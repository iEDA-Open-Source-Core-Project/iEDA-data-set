
module ysyx_040978_muler(
    input                   clock       ,
    input                   reset       ,// high active
    input                   in_valid    ,// 为高表示输入的数据有效，如果没有新的乘法输入，在乘法被接受的下一个周期要置低
    // input                   mulw        ,// 为高表示是 32 位乘法
    input     [1 : 0]       mul_signed  ,// 2'b11（signed x signed）；2'b10（signed x unsigned）；2'b00（unsigned x unsigned）；
    input     [63 : 0]      multiplicand,// 被乘数，xlen 表示乘法器位数
    input     [63 : 0]      multiplier  ,// 乘数

    output                  out_valid   ,// 高表示乘法器输出的结果有效
    output    [63 : 0]      result_hi   ,// 高 xlen bits 结果
    output    [63 : 0]      result_lo    // 低 xlen bits 结果    
  );
    //
    wire [64 : 0] multiplier_0;//符号位扩展
    wire [64 : 0] multiplicand_0;
    assign multiplier_0 = mul_signed[0] == 1'b1 ? {multiplier[63], multiplier} : {1'b0, multiplier};//1 is signed, 0 is unsigned
    assign multiplicand_0 = mul_signed[1] == 1'b1 ? {multiplicand[63], multiplicand} : {1'b0, multiplicand};//1 is signed, 0 is unsigned
    

    reg [5:0] cnt;
    reg mul_valid;
    wire mul_finish;
    reg  mul_ready, mul_busy;
    wire [128 : 0] p;//部分积

    always @(posedge clock) begin
        if(reset) cnt <= 6'd0;
        else if(cnt == 6'd32) cnt <= 6'd0;
        else if(mul_valid) cnt <= 6'd0;
        else if(in_valid | mul_busy) cnt <= cnt + 'h1;
        else cnt <= 6'd0;
    end

    reg  [65 : 0] multiplier_1;//乘数右移,取低三位
    wire [65 : 0] multiplier_2;

    always @(posedge clock) begin
        if(reset) multiplier_1 <= 'h0;
        else if(in_valid & mul_ready) multiplier_1 <= $signed({multiplier_0, 1'b0}) >>> 2;
        else if(mul_finish) multiplier_1 <= 'h0;
        else if(mul_busy) multiplier_1 <= $signed(multiplier_1) >>> 66'd2;
        else multiplier_1 <= 'h0;
    end


    reg [64 : 0] multiplicand_1;
    // wire [64 : 0] multiplicand_2;
    always @(posedge clock) begin
        if(reset) multiplicand_1 <= 'h0;
        else if(in_valid & mul_ready) multiplicand_1 <= multiplicand_0;
        else if(mul_finish) multiplicand_1 <= 'h0;
        else if(mul_busy) multiplicand_1 <= multiplicand_1;
        else multiplicand_1 <= 'h0;
    end

    assign multiplier_2 = (in_valid & mul_ready) ? {multiplier_0, 1'b0} : multiplier_1;
    // assign multiplicand_2 = (in_valid & mul_ready) ? multiplicand_0 : multiplicand_1;
    reg [128 : 0] result_buf;
    always @(posedge clock) begin
        if(reset) result_buf <= 'd0;
        else if(mul_busy) result_buf <= result_buf + p;
        else if(in_valid & mul_ready) result_buf <= p;
        else if(mul_valid) result_buf <= 'd0;
        else result_buf <= result_buf;
    end

    /* partial product */
    wire [128 : 0] pm_p;
    ysyx_040978_booth_pmgen u(.y_in(multiplier_2[2 : 0]), .x_in(multiplicand_0), .p(pm_p));
    assign p = pm_p << 2*cnt;
 

    /* control signal */

    always @(posedge clock) begin
        if(reset)begin
            mul_ready <= 1'b1;
        end else if(mul_finish)begin
            mul_ready <= 1'b1;
        end else if (in_valid)begin
            mul_ready <= 1'b0;
        end else begin
            mul_ready <= mul_ready;
        end
    end


    always @(posedge clock) begin
        if(reset)begin
            mul_busy <= 1'b0;
        end else if(mul_finish)begin
            mul_busy <= 1'b0;
        end else if(in_valid)begin
            mul_busy <= 1'b1;
        end else begin
            mul_busy <= mul_busy;
        end
    end

    assign mul_finish = cnt == 6'd32;
    
    /* output */

    always @(posedge clock) begin
        if(reset)   mul_valid <= 1'b0;
        else if(cnt == 6'd32) mul_valid <= 1'b1;
        else mul_valid <= 1'b0;
    end

    assign out_valid = mul_valid;

    assign result_hi = mul_valid ? result_buf[127 : 64] : 'd0;
    assign result_lo = mul_valid ? result_buf[63 : 0]   : 'd0;

endmodule

module ysyx_040978_mdu (
  input             clock   ,
  input             reset   ,
  input             mul     ,
  input             mulh    ,
  input             mulhu   ,
  input             mulhsu  ,
  input             div     ,
  input             divu    ,
  input             rem     ,
  input             remu    ,
  input   [63: 0]   src1    ,
  input   [63: 0]   src2    ,
  output  [63: 0]   result  ,
  output            ready 
);

  ///////////例化////////////
  wire    d_i_valid, d_i_signed;
  assign  d_i_valid = div | divu | rem | remu;
  assign  d_i_signed = div | rem;
  wire    d_o_valid;
  wire [63:0] d_o_q, d_o_r, d_res;
  ///////////除法器//////////
  ysyx_040978_diver du(
    .clock     (clock),
    .reset     (reset),
    .in_valid  (d_i_valid & ~d_o_valid),
    .div_signed(d_i_signed),
    .dividend  (src1),
    .divisor   (src2),
    
    .out_valid (d_o_valid),
    .quotient  (d_o_q),
    .remainder (d_o_r)
    );
  assign d_res = (div | divu) ? d_o_q : d_o_r;
  ///////////非法除法检查//////
  ///////////乘法器//////////
  wire m_i_valid;
  assign m_i_valid = mul | mulh | mulhu |mulhsu;
  wire [1:0] m_i_signed;
  assign m_i_signed[0] = mul | mulh;
  assign m_i_signed[1] = mul | mulh | mulhsu;
  wire [63:0] m_o_hi, m_o_lo, m_res;
  wire m_o_valid;

  ysyx_040978_muler mu(
    .clock       (clock),
    .reset       (reset),// high active
    .in_valid    (m_i_valid & ~m_o_valid),// 为高表示输入的数据有效，如果没有新的乘法输入，在乘法被接受的下一个周期要置低
    .mul_signed  (m_i_signed),// 2'b11（signed x signed）；2'b10（signed x unsigned）；2'b00（unsigned x unsigned）；
    .multiplicand(src1),// 被乘数，xlen 表示乘法器位数
    .multiplier  (src2),// 乘数

    .out_valid   (m_o_valid),// 高表示乘法器输出的结果有效
    .result_hi   (m_o_hi),// 高 xlen bits 结果
    .result_lo   (m_o_lo)// 低 xlen bits 结果    
  );
  assign m_res =  mul   ? m_o_lo : m_o_hi;

  ///////////输出////////////
  assign result = d_i_valid ? d_res : m_res;
  assign ready = d_o_valid | m_o_valid | ~(d_i_valid | m_i_valid) ;//d_o_ready & m_o_ready;

endmodule

module ysyx_040978_diver(
    input                   clock       ,
    input                   reset       ,// high active
    input                   in_valid   ,// 为高表示输入的数据有效，如果没有新的乘法输入，在乘法被接受的下一个周期要置低
    // input                   divw        ,// 为高表示是 32 位乘法
    input                   div_signed  ,// 表示是不是有符号除法，为高表示是有符号除法
    input     [63 : 0]      dividend    ,// 被除数，xlen 表示除法器位数
    input     [63 : 0]      divisor     ,// 除数

    output                  out_valid   ,// 高表示乘法器输出的结果有效
    output    [63 : 0]      quotient    ,// 商
    output    [63 : 0]      remainder    // 余数
  );
    //
    reg [6:0] cnt;
    reg valid;
    reg  ready, busy;
    wire finish;
    reg [191 : 0] dividend_1;

    always @(posedge clock) begin
        if(reset) cnt <= 'd63;
        else if(cnt == 'd0) cnt <= 'd63;
        else if(in_valid | busy) cnt <= cnt - 'd1;
        else cnt <= 'd63;
    end

    // 符号位缓存
    reg dsor_neg, dend_neg, div_signed_1;
    always @(posedge clock) begin
        if(reset)begin
            dsor_neg <= 1'b1;
            dend_neg <= 1'b1;
            div_signed_1 <= 1'b0;
        end else if(in_valid & ready)begin
            if(div_signed)begin
                dsor_neg <= divisor[63];
                dend_neg <= dividend[63];
                div_signed_1 <= 1'b1;
            end else begin
                dsor_neg <= 1'b0;
                dend_neg <= 1'b0;
                div_signed_1 <= 1'b0;
            end
        end else begin
            dsor_neg <= dsor_neg;
            dend_neg <= dend_neg;
            div_signed_1 <= div_signed_1;
        end
    end
    // 输入除数被除数绝对值计算
    wire [63:0] dividend_0;
    wire [63:0] divisor_0;
    ysyx_040978_MuxKey #(2, 1, 64) i2 (dividend_0, dividend[63] & div_signed, {1'b0, dividend, 1'b1, (~dividend + 64'b1)});
    ysyx_040978_MuxKey #(2, 1, 64) i3 (divisor_0,  divisor [63] & div_signed, {1'b0, divisor , 1'b1, (~divisor + 64'b1)});
    // assign dividend_0 = dividend[63] & div_signed ? (~dividend + 64'b1) : dividend;
    // assign divisor_0  = divisor [63] & div_signed ? (~divisor + 64'b1) : divisor;
    //除数缓存
    reg  [64 : 0] divisor_1;
    wire [64 : 0] divisor_2;
    always @(posedge clock) begin
        if(reset) divisor_1 <= 'h0;
        else if(in_valid & ready) divisor_1 <= {1'b0, divisor_0};
        else if(finish) divisor_1 <= 'h0;
        else divisor_1 <= divisor_1;
    end
    ysyx_040978_MuxKey #(2, 1, 65) i4 (divisor_2,  (in_valid==1'b1 && ready==1'b1), {1'b0, divisor_1 , 1'b1, {1'b0, divisor_0}});
    // assign divisor_2 = (in_valid==1'b1 && ready==1'b1) ? {1'b0, divisor_0} : divisor_1;
    //试商法,减数
    wire [64:0] subor;
    assign subor = divisor_2[64:0];
    wire [64:0] subend;
    ysyx_040978_MuxKey #(2, 1, 65) i5 (subend,  (in_valid & ready), {1'b0, dividend_1[127:63] , 1'b1, {64'h0, dividend_0[63]}});
    // assign subend = (in_valid & ready) ? {64'h0, dividend_0[63]} : dividend_1[127:63];
    wire [64:0] subres;
    assign subres = subend - subor;
    wire subneg;
    assign subneg = subres[64];

    //被除数,商,余数逻辑
    always @(posedge clock) begin
        if(reset) dividend_1 <= 'h0;
        else if(in_valid & ready)begin
            if(subneg) dividend_1 <= ({128'h0, dividend_0})<<1;//64 + 64 + 64
            else        dividend_1 <= ({64'h0, subres, dividend_0[62:0]})<<1;
        end else if(valid)begin
            dividend_1 <= 'h0;
        end else if(busy)begin
            if(subneg) dividend_1 <= dividend_1 << 1;
            else        dividend_1 <= ({dividend_1[191:128], subres, dividend_1[62:0]})<<1;
        end else begin
            dividend_1 <= dividend_1;
        end
    end

    reg [63:0] q;
    always @(posedge clock) begin
        if(reset)begin
            q <= 64'h0;
        end else if(in_valid & ready)begin
            if(subneg) q[cnt[5:0]] <= 1'b0;
            else q[cnt[5:0]] <= 1'b1;
        end else if(busy)begin
            if(subneg) q[cnt[5:0]] <= 1'b0;
            else q[cnt[5:0]] <= 1'b1;
        end else if(valid)begin
            q <= 64'h0;
        end else begin
            q <= q;
        end
    end

    /* control signal */
    always @(posedge clock) begin
        if(reset)begin
            ready <= 1'b1;
        end else if(finish)begin
            ready <= 1'b1;
        end else if (in_valid)begin
            ready <= 1'b0;
        end else begin
            ready <= ready;
        end
    end
    always @(posedge clock) begin
        if(reset)begin
            busy <= 1'b0;
        end else if(finish)begin
            busy <= 1'b0;
        end else if(in_valid)begin
            busy <= 1'b1;
        end else begin
            busy <= busy;
        end
    end

    assign finish = cnt == 'd0;
    
    /* output */
    always @(posedge clock) begin
        if(reset)   valid <= 1'b0;
        else if(cnt == 'd0) valid <= 1'b1;
        else valid <= 1'b0;
    end

    assign out_valid = valid;

    wire [63:0] q_neg;
    wire [63:0] r_neg;
    wire [63:0] q_pos;
    wire [63:0] r_pos;
    assign q_pos = q;
    assign r_pos = dividend_1[127:64];
    assign q_neg = (~q_pos) + 1'b1;
    assign r_neg = (~r_pos) + 1'b1;

    // assign remainder = dend_neg == 1'b1    ? r_neg : r_pos;
    // assign quotient  = dend_neg ^ dsor_neg ? q_neg : q_pos;
    ysyx_040978_MuxKey #(2, 1, 64) i0 (remainder, dend_neg, { 1'b0, r_pos, 1'b1, r_neg});

    wire den_neg_xor = dend_neg ^ dsor_neg;
    ysyx_040978_MuxKey #(2, 1, 64) i1 (quotient, den_neg_xor, { 1'b0, q_pos, 1'b1, q_neg});
endmodule

module ysyx_040978_booth_pmgen
(
  input     [2   : 0]     y_in,
  input     [64  : 0]     x_in,
  output    [128 : 0]     p
  // output                c//负数补码(-[X]补, -2[X]补), 末位+1信号
);

//booth选择信号的生成
    wire y_add,y,y_sub;
    assign {y_add,y,y_sub} = y_in;
    
    
    wire sel_neg, sel_dneg, sel_pos, sel_dpos;
    
    assign sel_neg =  y_add & (y & ~y_sub | ~y & y_sub);
    assign sel_pos = ~y_add & (y & ~y_sub | ~y & y_sub);
    assign sel_dneg =  y_add & ~y & ~y_sub;
    assign sel_dpos = ~y_add &  y &  y_sub;
    
    //结果选择逻辑
    wire [128 : 0] x_in_129;
    wire [128 : 0] p_pos, p_neg, p_dpos, p_dneg;

    assign x_in_129 = {{64{x_in[64]}}, x_in};
    assign p_pos = x_in_129;
    assign p_neg = ~x_in_129 + 128'b1;
    assign p_dpos = x_in_129 << 1;
    assign p_dneg = p_neg << 1; 
    
    assign p =  sel_pos ? p_pos :
                sel_dpos? p_dpos:
                sel_neg ? p_neg :
                sel_dneg? p_dneg: {129{1'b0}};

endmodule

module ysyx_040978_Interconnect3x1(
  input         clock,
  input         reset,
  input         io_maxi_ar_ready,
  output        io_maxi_ar_valid,
  output [31:0] io_maxi_ar_bits_addr,
  output [3:0]  io_maxi_ar_bits_id,
  output [7:0]  io_maxi_ar_bits_len,
  output [2:0]  io_maxi_ar_bits_size,
  input         io_maxi_r_valid,
  input  [63:0] io_maxi_r_bits_data,
  input  [3:0]  io_maxi_r_bits_id,
  input         io_maxi_r_bits_last,
  input         io_maxi_aw_ready,
  output        io_maxi_aw_valid,
  output [31:0] io_maxi_aw_bits_addr,
  output [3:0]  io_maxi_aw_bits_id,
  output [7:0]  io_maxi_aw_bits_len,
  output [2:0]  io_maxi_aw_bits_size,
  input         io_maxi_w_ready,
  output        io_maxi_w_valid,
  output [63:0] io_maxi_w_bits_data,
  output [7:0]  io_maxi_w_bits_strb,
  output        io_maxi_w_bits_last,
  input         io_maxi_b_valid,
  input  [3:0]  io_maxi_b_bits_id,
  output        io_ifu_ar_ready,
  input         io_ifu_ar_valid,
  input  [31:0] io_ifu_ar_bits_addr,
  input  [7:0]  io_ifu_ar_bits_len,
  input  [2:0]  io_ifu_ar_bits_size,
  output        io_ifu_r_valid,
  output [63:0] io_ifu_r_bits_data,
  output        io_ifu_r_bits_last,
  output        io_memu_ar_ready,
  input         io_memu_ar_valid,
  input  [31:0] io_memu_ar_bits_addr,
  input  [7:0]  io_memu_ar_bits_len,
  input  [2:0]  io_memu_ar_bits_size,
  output        io_memu_r_valid,
  output [63:0] io_memu_r_bits_data,
  output        io_memu_r_bits_last,
  output        io_memu_aw_ready,
  input         io_memu_aw_valid,
  input  [31:0] io_memu_aw_bits_addr,
  input  [7:0]  io_memu_aw_bits_len,
  input  [2:0]  io_memu_aw_bits_size,
  output        io_memu_w_ready,
  input         io_memu_w_valid,
  input  [63:0] io_memu_w_bits_data,
  input  [7:0]  io_memu_w_bits_strb,
  input         io_memu_w_bits_last,
  output        io_memu_b_valid,
  output        io_devu_ar_ready,
  input         io_devu_ar_valid,
  input  [31:0] io_devu_ar_bits_addr,
  input  [2:0]  io_devu_ar_bits_size,
  output        io_devu_r_valid,
  output [63:0] io_devu_r_bits_data,
  output        io_devu_r_bits_last,
  output        io_devu_aw_ready,
  input         io_devu_aw_valid,
  input  [31:0] io_devu_aw_bits_addr,
  input  [2:0]  io_devu_aw_bits_size,
  output        io_devu_w_ready,
  input         io_devu_w_valid,
  input  [63:0] io_devu_w_bits_data,
  input  [7:0]  io_devu_w_bits_strb,
  input         io_devu_w_bits_last,
  output        io_devu_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] axi_reading; // @[AXI.scala 131:36]
  wire  _T = axi_reading == 4'h0; // @[AXI.scala 133:35]
  wire  _io_memu_ar_ready_T = ~io_devu_ar_valid; // @[AXI.scala 140:37]
  wire [2:0] _GEN_2 = io_ifu_ar_valid ? io_ifu_ar_bits_size : 3'h0; // @[AXI.scala 152:27 AXI.scala 153:18 AXI.scala 310:19]
  wire [7:0] _GEN_3 = io_ifu_ar_valid ? io_ifu_ar_bits_len : 8'h0; // @[AXI.scala 152:27 AXI.scala 153:18 AXI.scala 311:19]
  wire [3:0] _GEN_4 = io_ifu_ar_valid ? 4'h1 : 4'h0; // @[AXI.scala 152:27 AXI.scala 155:21 AXI.scala 308:17]
  wire [31:0] _GEN_6 = io_ifu_ar_valid ? io_ifu_ar_bits_addr : 32'h0; // @[AXI.scala 152:27 AXI.scala 153:18 AXI.scala 309:19]
  wire [2:0] _GEN_8 = io_memu_ar_valid ? io_memu_ar_bits_size : _GEN_2; // @[AXI.scala 148:28 AXI.scala 149:18]
  wire [7:0] _GEN_9 = io_memu_ar_valid ? io_memu_ar_bits_len : _GEN_3; // @[AXI.scala 148:28 AXI.scala 149:18]
  wire [3:0] _GEN_10 = io_memu_ar_valid ? 4'h2 : _GEN_4; // @[AXI.scala 148:28 AXI.scala 151:21]
  wire [31:0] _GEN_12 = io_memu_ar_valid ? io_memu_ar_bits_addr : _GEN_6; // @[AXI.scala 148:28 AXI.scala 149:18]
  wire  _GEN_13 = io_memu_ar_valid | io_ifu_ar_valid; // @[AXI.scala 148:28 AXI.scala 150:19]
  wire [2:0] _GEN_14 = io_devu_ar_valid ? io_devu_ar_bits_size : _GEN_8; // @[AXI.scala 144:28 AXI.scala 145:18]
  wire [7:0] _GEN_15 = io_devu_ar_valid ? 8'h0 : _GEN_9; // @[AXI.scala 144:28 AXI.scala 145:18]
  wire [3:0] _GEN_16 = io_devu_ar_valid ? 4'h3 : _GEN_10; // @[AXI.scala 144:28 AXI.scala 147:21]
  wire [31:0] _GEN_18 = io_devu_ar_valid ? io_devu_ar_bits_addr : _GEN_12; // @[AXI.scala 144:28 AXI.scala 145:18]
  wire  _GEN_19 = io_devu_ar_valid | _GEN_13; // @[AXI.scala 144:28 AXI.scala 146:19]
  wire  _GEN_26 = io_maxi_r_bits_id == 4'h1 & io_maxi_r_valid; // @[AXI.scala 165:40 AXI.scala 166:18 AXI.scala 333:15]
  wire  _GEN_32 = io_maxi_r_bits_id == 4'h1 ? 1'h0 : io_maxi_r_bits_last; // @[AXI.scala 165:40 AXI.scala 337:19 AXI.scala 169:19]
  wire [63:0] _GEN_34 = io_maxi_r_bits_id == 4'h1 ? 64'h0 : io_maxi_r_bits_data; // @[AXI.scala 165:40 AXI.scala 336:19 AXI.scala 169:19]
  wire  _GEN_35 = io_maxi_r_bits_id == 4'h2 & io_maxi_r_valid; // @[AXI.scala 162:41 AXI.scala 163:19 AXI.scala 333:15]
  wire  _GEN_37 = io_maxi_r_bits_id == 4'h2 ? io_maxi_r_bits_last : _GEN_32; // @[AXI.scala 162:41 AXI.scala 164:19]
  wire [63:0] _GEN_39 = io_maxi_r_bits_id == 4'h2 ? io_maxi_r_bits_data : _GEN_34; // @[AXI.scala 162:41 AXI.scala 164:19]
  wire  _GEN_40 = io_maxi_r_bits_id == 4'h2 ? 1'h0 : _GEN_26; // @[AXI.scala 162:41 AXI.scala 333:15]
  wire  _GEN_42 = io_maxi_r_bits_id == 4'h2 ? 1'h0 : io_maxi_r_bits_last; // @[AXI.scala 162:41 AXI.scala 337:19]
  wire [63:0] _GEN_44 = io_maxi_r_bits_id == 4'h2 ? 64'h0 : io_maxi_r_bits_data; // @[AXI.scala 162:41 AXI.scala 336:19]
  wire  _GEN_46 = io_maxi_r_bits_id == 4'h2 ? 1'h0 : _GEN_32; // @[AXI.scala 162:41 AXI.scala 337:19]
  wire [63:0] _GEN_48 = io_maxi_r_bits_id == 4'h2 ? 64'h0 : _GEN_34; // @[AXI.scala 162:41 AXI.scala 336:19]
  reg  dev_writing; // @[AXI.scala 179:36]
  reg  mem_writing; // @[AXI.scala 180:36]
  wire  _T_10 = io_maxi_b_bits_id == 4'h3; // @[AXI.scala 183:46]
  wire  _GEN_64 = io_maxi_b_valid & io_maxi_b_bits_id == 4'h3 ? 1'h0 : dev_writing; // @[AXI.scala 183:59 AXI.scala 183:73 AXI.scala 179:36]
  wire  _GEN_65 = io_maxi_aw_valid & io_maxi_aw_bits_id == 4'h3 | _GEN_64; // @[AXI.scala 182:59 AXI.scala 182:73]
  wire  _GEN_66 = io_maxi_b_valid & io_maxi_b_bits_id == 4'h2 ? 1'h0 : mem_writing; // @[AXI.scala 185:59 AXI.scala 185:73 AXI.scala 180:36]
  wire  _GEN_67 = io_maxi_aw_valid & io_maxi_aw_bits_id == 4'h2 | _GEN_66; // @[AXI.scala 184:59 AXI.scala 184:73]
  wire  _io_devu_aw_ready_T = ~mem_writing; // @[AXI.scala 187:37]
  wire  _io_memu_aw_ready_T_2 = ~dev_writing; // @[AXI.scala 188:56]
  wire [2:0] _GEN_68 = io_memu_aw_valid ? io_memu_aw_bits_size : io_devu_aw_bits_size; // @[AXI.scala 193:28 AXI.scala 194:18 AXI.scala 174:11]
  wire [7:0] _GEN_69 = io_memu_aw_valid ? io_memu_aw_bits_len : 8'h0; // @[AXI.scala 193:28 AXI.scala 194:18 AXI.scala 174:11]
  wire [3:0] _GEN_70 = io_memu_aw_valid ? 4'h2 : 4'h0; // @[AXI.scala 193:28 AXI.scala 196:21 AXI.scala 174:11]
  wire [31:0] _GEN_72 = io_memu_aw_valid ? io_memu_aw_bits_addr : io_devu_aw_bits_addr; // @[AXI.scala 193:28 AXI.scala 194:18 AXI.scala 174:11]
  wire  _GEN_73 = io_memu_aw_valid | io_devu_aw_valid; // @[AXI.scala 193:28 AXI.scala 195:19 AXI.scala 174:11]
  wire  _GEN_80 = mem_writing ? io_memu_w_bits_last : io_devu_w_bits_last; // @[AXI.scala 204:26 AXI.scala 205:17 AXI.scala 175:10]
  wire [7:0] _GEN_81 = mem_writing ? io_memu_w_bits_strb : io_devu_w_bits_strb; // @[AXI.scala 204:26 AXI.scala 205:17 AXI.scala 175:10]
  wire [63:0] _GEN_82 = mem_writing ? io_memu_w_bits_data : io_devu_w_bits_data; // @[AXI.scala 204:26 AXI.scala 205:17 AXI.scala 175:10]
  wire  _GEN_83 = mem_writing ? io_memu_w_valid : io_devu_w_valid; // @[AXI.scala 204:26 AXI.scala 206:18 AXI.scala 175:10]
  assign io_maxi_ar_valid = axi_reading != 4'h0 ? 1'h0 : _GEN_19; // @[AXI.scala 142:32 AXI.scala 307:15]
  assign io_maxi_ar_bits_addr = axi_reading != 4'h0 ? 32'h0 : _GEN_18; // @[AXI.scala 142:32 AXI.scala 309:19]
  assign io_maxi_ar_bits_id = axi_reading != 4'h0 ? 4'h0 : _GEN_16; // @[AXI.scala 142:32 AXI.scala 308:17]
  assign io_maxi_ar_bits_len = axi_reading != 4'h0 ? 8'h0 : _GEN_15; // @[AXI.scala 142:32 AXI.scala 311:19]
  assign io_maxi_ar_bits_size = axi_reading != 4'h0 ? 3'h0 : _GEN_14; // @[AXI.scala 142:32 AXI.scala 310:19]
  assign io_maxi_aw_valid = io_devu_aw_valid | _GEN_73; // @[AXI.scala 189:22 AXI.scala 191:19]
  assign io_maxi_aw_bits_addr = io_devu_aw_valid ? io_devu_aw_bits_addr : _GEN_72; // @[AXI.scala 189:22 AXI.scala 190:18]
  assign io_maxi_aw_bits_id = io_devu_aw_valid ? 4'h3 : _GEN_70; // @[AXI.scala 189:22 AXI.scala 192:21]
  assign io_maxi_aw_bits_len = io_devu_aw_valid ? 8'h0 : _GEN_69; // @[AXI.scala 189:22 AXI.scala 190:18]
  assign io_maxi_aw_bits_size = io_devu_aw_valid ? io_devu_aw_bits_size : _GEN_68; // @[AXI.scala 189:22 AXI.scala 190:18]
  assign io_maxi_w_valid = dev_writing ? io_devu_w_valid : _GEN_83; // @[AXI.scala 201:20 AXI.scala 203:18]
  assign io_maxi_w_bits_data = dev_writing ? io_devu_w_bits_data : _GEN_82; // @[AXI.scala 201:20 AXI.scala 202:17]
  assign io_maxi_w_bits_strb = dev_writing ? io_devu_w_bits_strb : _GEN_81; // @[AXI.scala 201:20 AXI.scala 202:17]
  assign io_maxi_w_bits_last = dev_writing ? io_devu_w_bits_last : _GEN_80; // @[AXI.scala 201:20 AXI.scala 202:17]
  assign io_ifu_ar_ready = io_maxi_ar_ready & ~io_memu_ar_valid & _io_memu_ar_ready_T & _T; // @[AXI.scala 141:72]
  assign io_ifu_r_valid = io_maxi_r_bits_id == 4'h3 ? 1'h0 : _GEN_40; // @[AXI.scala 159:35 AXI.scala 333:15]
  assign io_ifu_r_bits_data = io_maxi_r_bits_id == 4'h3 ? 64'h0 : _GEN_44; // @[AXI.scala 159:35 AXI.scala 336:19]
  assign io_ifu_r_bits_last = io_maxi_r_bits_id == 4'h3 ? 1'h0 : _GEN_42; // @[AXI.scala 159:35 AXI.scala 337:19]
  assign io_memu_ar_ready = io_maxi_ar_ready & ~io_devu_ar_valid & _T; // @[AXI.scala 140:54]
  assign io_memu_r_valid = io_maxi_r_bits_id == 4'h3 ? 1'h0 : _GEN_35; // @[AXI.scala 159:35 AXI.scala 333:15]
  assign io_memu_r_bits_data = io_maxi_r_bits_id == 4'h3 ? 64'h0 : _GEN_39; // @[AXI.scala 159:35 AXI.scala 336:19]
  assign io_memu_r_bits_last = io_maxi_r_bits_id == 4'h3 ? 1'h0 : _GEN_37; // @[AXI.scala 159:35 AXI.scala 337:19]
  assign io_memu_aw_ready = io_maxi_aw_ready & ~io_devu_aw_valid & ~dev_writing; // @[AXI.scala 188:53]
  assign io_memu_w_ready = io_maxi_w_ready & _io_memu_aw_ready_T_2; // @[AXI.scala 200:32]
  assign io_memu_b_valid = _T_10 ? 1'h0 : io_maxi_b_valid; // @[AXI.scala 211:35 AXI.scala 379:15]
  assign io_devu_ar_ready = io_maxi_ar_ready & _T; // @[AXI.scala 139:34]
  assign io_devu_r_valid = io_maxi_r_bits_id == 4'h3 & io_maxi_r_valid; // @[AXI.scala 159:35 AXI.scala 160:19 AXI.scala 333:15]
  assign io_devu_r_bits_data = io_maxi_r_bits_id == 4'h3 ? io_maxi_r_bits_data : _GEN_48; // @[AXI.scala 159:35 AXI.scala 161:19]
  assign io_devu_r_bits_last = io_maxi_r_bits_id == 4'h3 ? io_maxi_r_bits_last : _GEN_46; // @[AXI.scala 159:35 AXI.scala 161:19]
  assign io_devu_aw_ready = io_maxi_aw_ready & ~mem_writing; // @[AXI.scala 187:34]
  assign io_devu_w_ready = io_maxi_w_ready & _io_devu_aw_ready_T; // @[AXI.scala 199:32]
  assign io_devu_b_valid = io_maxi_b_valid; // @[AXI.scala 211:35 AXI.scala 212:19 AXI.scala 176:10]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 131:36]
      axi_reading <= 4'h0; // @[AXI.scala 131:36]
    end else if (io_maxi_ar_valid & axi_reading == 4'h0 & io_maxi_ar_ready) begin // @[AXI.scala 133:62]
      axi_reading <= io_maxi_ar_bits_id; // @[AXI.scala 134:17]
    end else if (io_maxi_r_valid & io_maxi_r_bits_last) begin // @[AXI.scala 135:46]
      axi_reading <= 4'h0; // @[AXI.scala 136:17]
    end
    if (reset) begin // @[AXI.scala 179:36]
      dev_writing <= 1'h0; // @[AXI.scala 179:36]
    end else begin
      dev_writing <= _GEN_65;
    end
    if (reset) begin // @[AXI.scala 180:36]
      mem_writing <= 1'h0; // @[AXI.scala 180:36]
    end else begin
      mem_writing <= _GEN_67;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  axi_reading = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  dev_writing = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_writing = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_PC(
  input         clock,
  input         reset,
  input         io_jump0,
  input         io_jump,
  input  [63:0] io_npc,
  input         io_sys_ready,
  input         io_next_ready,
  output        io_next_valid,
  output [63:0] io_next_bits_pc2if_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pc_reg_x3 = (io_next_ready | io_jump) & io_sys_ready; // @[IFU.scala 27:109]
  reg [63:0] pc_reg; // @[Reg.scala 27:20]
  wire  _pc_reg_in_T = ~io_next_ready; // @[IFU.scala 33:6]
  wire [63:0] inc_pc_out = pc_reg + 64'h4; // @[IFU.scala 28:27]
  reg  start; // @[Reg.scala 27:20]
  wire  _GEN_1 = io_sys_ready | start; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _io_next_valid_T_1 = io_jump0 ? 1'h0 : start; // @[Mux.scala 98:16]
  assign io_next_valid = reset ? 1'h0 : _io_next_valid_T_1; // @[Mux.scala 98:16]
  assign io_next_bits_pc2if_pc = pc_reg; // @[IFU.scala 40:15]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      pc_reg <= 64'h30000000; // @[Reg.scala 27:20]
    end else if (pc_reg_x3) begin // @[Reg.scala 28:19]
      if (io_jump) begin // @[Mux.scala 98:16]
        pc_reg <= io_npc;
      end else if (!(_pc_reg_in_T)) begin // @[Mux.scala 98:16]
        pc_reg <= inc_pc_out;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      start <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      start <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_reg = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  start = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_IAXIManager(
  input          clock,
  input          reset,
  input          io_in_rd_en,
  input          io_in_dev,
  input  [31:0]  io_in_addr,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  output         io_out_finish,
  output         io_out_ready,
  output [127:0] io_out_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [127:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] curr_state; // @[AXI4Manager.scala 85:35]
  reg  stage_out2_rd_en; // @[Reg.scala 27:20]
  reg  stage_out2_dev; // @[Reg.scala 27:20]
  reg [31:0] stage_out2_addr; // @[Reg.scala 27:20]
  wire  stage_en = curr_state == 2'h0; // @[AXI4Manager.scala 110:26]
  wire [31:0] _GEN_0 = stage_en ? io_in_addr : stage_out2_addr; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_1 = stage_en ? io_in_dev : stage_out2_dev; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_2 = stage_en ? io_in_rd_en : stage_out2_rd_en; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  r_last = io_maxi_r_bits_last & io_maxi_r_valid; // @[AXI4Manager.scala 105:42]
  wire [7:0] a_len = _GEN_1 ? 8'h0 : 8'h1; // @[AXI4Manager.scala 115:31]
  wire [29:0] a_addr_hi = _GEN_0[31:2]; // @[AXI4Manager.scala 116:52]
  wire [31:0] _a_addr_T = {a_addr_hi,2'h0}; // @[Cat.scala 30:58]
  wire [27:0] a_addr_hi_1 = _GEN_0[31:4]; // @[AXI4Manager.scala 116:84]
  wire [31:0] _a_addr_T_1 = {a_addr_hi_1,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] a_addr = _GEN_1 ? _a_addr_T : _a_addr_T_1; // @[AXI4Manager.scala 116:31]
  wire [1:0] a_size = _GEN_1 ? 2'h2 : 2'h3; // @[AXI4Manager.scala 117:31]
  wire [5:0] _start_bit_T_1 = {_GEN_0[2:0], 3'h0}; // @[AXI4Manager.scala 118:55]
  wire [5:0] start_bit = _GEN_1 ? _start_bit_T_1 : _start_bit_T_1; // @[AXI4Manager.scala 118:31]
  wire  rdata64_x8 = io_maxi_r_valid & ~io_maxi_r_bits_last; // @[AXI4Manager.scala 120:101]
  reg [63:0] memory_data_lo; // @[Reg.scala 27:20]
  wire [63:0] _memory_data_T = io_maxi_r_bits_data >> start_bit; // @[AXI4Manager.scala 121:58]
  wire [127:0] _memory_data_T_1 = {io_maxi_r_bits_data,memory_data_lo}; // @[Cat.scala 30:58]
  wire [127:0] memory_data = _GEN_1 ? {{64'd0}, _memory_data_T} : _memory_data_T_1; // @[AXI4Manager.scala 121:32]
  wire  _T = 2'h0 == curr_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_4 = io_maxi_ar_ready ? 2'h2 : 2'h1; // @[AXI4Manager.scala 129:29 AXI4Manager.scala 129:42 AXI4Manager.scala 129:79]
  wire [1:0] _GEN_5 = _GEN_2 ? _GEN_4 : 2'h0; // @[AXI4Manager.scala 128:20 AXI4Manager.scala 130:42]
  wire  _T_1 = 2'h1 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == curr_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_6 = ~_GEN_1 ? 2'h3 : 2'h2; // @[AXI4Manager.scala 135:32 AXI4Manager.scala 135:45 AXI4Manager.scala 136:60]
  wire [1:0] _GEN_7 = r_last ? 2'h0 : _GEN_6; // @[AXI4Manager.scala 134:45 AXI4Manager.scala 134:58]
  wire  _T_4 = 2'h3 == curr_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_8 = r_last ? 2'h0 : 2'h3; // @[AXI4Manager.scala 139:47 AXI4Manager.scala 139:60 AXI4Manager.scala 140:60]
  wire [1:0] _GEN_9 = _T_4 ? _GEN_8 : 2'h0; // @[Conditional.scala 39:67 AXI4Manager.scala 125:14]
  wire [1:0] _GEN_10 = _T_2 ? _GEN_7 : _GEN_9; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_11 = _T_1 ? _GEN_4 : _GEN_10; // @[Conditional.scala 39:67]
  wire [1:0] next_state = _T ? _GEN_5 : _GEN_11; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_16 = next_state == 2'h2 | next_state == 2'h1 ? a_size : 2'h0; // @[AXI4Manager.scala 146:55 AXI.scala 318:19 AXI.scala 310:19]
  reg [127:0] memory_data_buffer; // @[AXI4Manager.scala 154:43]
  assign io_maxi_ar_valid = next_state == 2'h2 | next_state == 2'h1; // @[AXI4Manager.scala 146:30]
  assign io_maxi_ar_bits_addr = next_state == 2'h2 | next_state == 2'h1 ? a_addr : 32'h0; // @[AXI4Manager.scala 146:55 AXI.scala 317:19 AXI.scala 309:19]
  assign io_maxi_ar_bits_len = next_state == 2'h2 | next_state == 2'h1 ? a_len : 8'h0; // @[AXI4Manager.scala 146:55 AXI.scala 319:19 AXI.scala 311:19]
  assign io_maxi_ar_bits_size = {{1'd0}, _GEN_16}; // @[AXI4Manager.scala 146:55 AXI.scala 318:19 AXI.scala 310:19]
  assign io_out_finish = io_maxi_r_bits_last; // @[AXI4Manager.scala 153:34]
  assign io_out_ready = next_state == 2'h0 | stage_en; // @[AXI4Manager.scala 152:38]
  assign io_out_data = curr_state == 2'h2 | curr_state == 2'h3 ? memory_data : memory_data_buffer; // @[AXI4Manager.scala 156:18]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4Manager.scala 85:35]
      curr_state <= 2'h0; // @[AXI4Manager.scala 85:35]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_GEN_2) begin // @[AXI4Manager.scala 128:20]
        curr_state <= _GEN_4;
      end else begin
        curr_state <= 2'h0; // @[AXI4Manager.scala 130:42]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_4;
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_7;
    end else begin
      curr_state <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_dev <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_dev <= io_in_dev; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_addr <= io_in_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      memory_data_lo <= 64'h0; // @[Reg.scala 27:20]
    end else if (rdata64_x8) begin // @[Reg.scala 28:19]
      memory_data_lo <= io_maxi_r_bits_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[AXI4Manager.scala 154:43]
      memory_data_buffer <= 128'h0; // @[AXI4Manager.scala 154:43]
    end else if (io_out_finish) begin // @[AXI4Manager.scala 155:28]
      if (_GEN_1) begin // @[AXI4Manager.scala 121:32]
        memory_data_buffer <= {{64'd0}, _memory_data_T};
      end else begin
        memory_data_buffer <= _memory_data_T_1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  stage_out2_rd_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stage_out2_dev = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  stage_out2_addr = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  memory_data_lo = _RAND_4[63:0];
  _RAND_5 = {4{`RANDOM}};
  memory_data_buffer = _RAND_5[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_ICacheUnit(
  input          clock,
  input          reset,
  input          io_next_ready,
  output         io_next_valid,
  output [31:0]  io_next_bits_data_if2id_inst,
  output [63:0]  io_next_bits_data_if2id_pc,
  input          io_cache_reset,
  output         io_prev_ready,
  input          io_prev_valid,
  input  [38:0]  io_prev_bits_addr,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  output [5:0]   io_sram0_addr,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  input          fencei
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
`endif // RANDOMIZE_REG_INIT
  wire  maxi4_manager_clock; // @[ICache.scala 73:29]
  wire  maxi4_manager_reset; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_in_rd_en; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_in_dev; // @[ICache.scala 73:29]
  wire [31:0] maxi4_manager_io_in_addr; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_maxi_ar_ready; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_maxi_ar_valid; // @[ICache.scala 73:29]
  wire [31:0] maxi4_manager_io_maxi_ar_bits_addr; // @[ICache.scala 73:29]
  wire [7:0] maxi4_manager_io_maxi_ar_bits_len; // @[ICache.scala 73:29]
  wire [2:0] maxi4_manager_io_maxi_ar_bits_size; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_maxi_r_valid; // @[ICache.scala 73:29]
  wire [63:0] maxi4_manager_io_maxi_r_bits_data; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_maxi_r_bits_last; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_out_finish; // @[ICache.scala 73:29]
  wire  maxi4_manager_io_out_ready; // @[ICache.scala 73:29]
  wire [127:0] maxi4_manager_io_out_data; // @[ICache.scala 73:29]
  reg [2:0] curr_state; // @[ICache.scala 68:37]
  wire  _array_write_T = curr_state == 3'h4; // @[ICache.scala 278:29]
  wire  array_write = curr_state == 3'h4 & maxi4_manager_io_out_finish; // @[ICache.scala 278:39]
  reg [38:0] stage1_out_bits_addr; // @[Reg.scala 27:20]
  wire [5:0] stage1_index = stage1_out_bits_addr[9:4]; // @[ICache.scala 117:54]
  reg  lru_list_63; // @[ICache.scala 103:35]
  reg  lru_list_62; // @[ICache.scala 103:35]
  reg  lru_list_61; // @[ICache.scala 103:35]
  reg  lru_list_60; // @[ICache.scala 103:35]
  reg  lru_list_59; // @[ICache.scala 103:35]
  reg  lru_list_58; // @[ICache.scala 103:35]
  reg  lru_list_57; // @[ICache.scala 103:35]
  reg  lru_list_56; // @[ICache.scala 103:35]
  reg  lru_list_55; // @[ICache.scala 103:35]
  reg  lru_list_54; // @[ICache.scala 103:35]
  reg  lru_list_53; // @[ICache.scala 103:35]
  reg  lru_list_52; // @[ICache.scala 103:35]
  reg  lru_list_51; // @[ICache.scala 103:35]
  reg  lru_list_50; // @[ICache.scala 103:35]
  reg  lru_list_49; // @[ICache.scala 103:35]
  reg  lru_list_48; // @[ICache.scala 103:35]
  reg  lru_list_47; // @[ICache.scala 103:35]
  reg  lru_list_46; // @[ICache.scala 103:35]
  reg  lru_list_45; // @[ICache.scala 103:35]
  reg  lru_list_44; // @[ICache.scala 103:35]
  reg  lru_list_43; // @[ICache.scala 103:35]
  reg  lru_list_42; // @[ICache.scala 103:35]
  reg  lru_list_41; // @[ICache.scala 103:35]
  reg  lru_list_40; // @[ICache.scala 103:35]
  reg  lru_list_39; // @[ICache.scala 103:35]
  reg  lru_list_38; // @[ICache.scala 103:35]
  reg  lru_list_37; // @[ICache.scala 103:35]
  reg  lru_list_36; // @[ICache.scala 103:35]
  reg  lru_list_35; // @[ICache.scala 103:35]
  reg  lru_list_34; // @[ICache.scala 103:35]
  reg  lru_list_33; // @[ICache.scala 103:35]
  reg  lru_list_32; // @[ICache.scala 103:35]
  reg  lru_list_31; // @[ICache.scala 103:35]
  reg  lru_list_30; // @[ICache.scala 103:35]
  reg  lru_list_29; // @[ICache.scala 103:35]
  reg  lru_list_28; // @[ICache.scala 103:35]
  reg  lru_list_27; // @[ICache.scala 103:35]
  reg  lru_list_26; // @[ICache.scala 103:35]
  reg  lru_list_25; // @[ICache.scala 103:35]
  reg  lru_list_24; // @[ICache.scala 103:35]
  reg  lru_list_23; // @[ICache.scala 103:35]
  reg  lru_list_22; // @[ICache.scala 103:35]
  reg  lru_list_21; // @[ICache.scala 103:35]
  reg  lru_list_20; // @[ICache.scala 103:35]
  reg  lru_list_19; // @[ICache.scala 103:35]
  reg  lru_list_18; // @[ICache.scala 103:35]
  reg  lru_list_17; // @[ICache.scala 103:35]
  reg  lru_list_16; // @[ICache.scala 103:35]
  reg  lru_list_15; // @[ICache.scala 103:35]
  reg  lru_list_14; // @[ICache.scala 103:35]
  reg  lru_list_13; // @[ICache.scala 103:35]
  reg  lru_list_12; // @[ICache.scala 103:35]
  reg  lru_list_11; // @[ICache.scala 103:35]
  reg  lru_list_10; // @[ICache.scala 103:35]
  reg  lru_list_9; // @[ICache.scala 103:35]
  reg  lru_list_8; // @[ICache.scala 103:35]
  reg  lru_list_7; // @[ICache.scala 103:35]
  reg  lru_list_6; // @[ICache.scala 103:35]
  reg  lru_list_5; // @[ICache.scala 103:35]
  reg  lru_list_4; // @[ICache.scala 103:35]
  reg  lru_list_3; // @[ICache.scala 103:35]
  reg  lru_list_2; // @[ICache.scala 103:35]
  reg  lru_list_1; // @[ICache.scala 103:35]
  reg  lru_list_0; // @[ICache.scala 103:35]
  wire  _GEN_4 = 6'h1 == stage1_index ? lru_list_1 : lru_list_0; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_5 = 6'h2 == stage1_index ? lru_list_2 : _GEN_4; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_6 = 6'h3 == stage1_index ? lru_list_3 : _GEN_5; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_7 = 6'h4 == stage1_index ? lru_list_4 : _GEN_6; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_8 = 6'h5 == stage1_index ? lru_list_5 : _GEN_7; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_9 = 6'h6 == stage1_index ? lru_list_6 : _GEN_8; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_10 = 6'h7 == stage1_index ? lru_list_7 : _GEN_9; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_11 = 6'h8 == stage1_index ? lru_list_8 : _GEN_10; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_12 = 6'h9 == stage1_index ? lru_list_9 : _GEN_11; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_13 = 6'ha == stage1_index ? lru_list_10 : _GEN_12; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_14 = 6'hb == stage1_index ? lru_list_11 : _GEN_13; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_15 = 6'hc == stage1_index ? lru_list_12 : _GEN_14; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_16 = 6'hd == stage1_index ? lru_list_13 : _GEN_15; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_17 = 6'he == stage1_index ? lru_list_14 : _GEN_16; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_18 = 6'hf == stage1_index ? lru_list_15 : _GEN_17; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_19 = 6'h10 == stage1_index ? lru_list_16 : _GEN_18; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_20 = 6'h11 == stage1_index ? lru_list_17 : _GEN_19; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_21 = 6'h12 == stage1_index ? lru_list_18 : _GEN_20; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_22 = 6'h13 == stage1_index ? lru_list_19 : _GEN_21; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_23 = 6'h14 == stage1_index ? lru_list_20 : _GEN_22; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_24 = 6'h15 == stage1_index ? lru_list_21 : _GEN_23; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_25 = 6'h16 == stage1_index ? lru_list_22 : _GEN_24; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_26 = 6'h17 == stage1_index ? lru_list_23 : _GEN_25; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_27 = 6'h18 == stage1_index ? lru_list_24 : _GEN_26; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_28 = 6'h19 == stage1_index ? lru_list_25 : _GEN_27; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_29 = 6'h1a == stage1_index ? lru_list_26 : _GEN_28; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_30 = 6'h1b == stage1_index ? lru_list_27 : _GEN_29; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_31 = 6'h1c == stage1_index ? lru_list_28 : _GEN_30; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_32 = 6'h1d == stage1_index ? lru_list_29 : _GEN_31; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_33 = 6'h1e == stage1_index ? lru_list_30 : _GEN_32; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_34 = 6'h1f == stage1_index ? lru_list_31 : _GEN_33; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_35 = 6'h20 == stage1_index ? lru_list_32 : _GEN_34; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_36 = 6'h21 == stage1_index ? lru_list_33 : _GEN_35; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_37 = 6'h22 == stage1_index ? lru_list_34 : _GEN_36; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_38 = 6'h23 == stage1_index ? lru_list_35 : _GEN_37; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_39 = 6'h24 == stage1_index ? lru_list_36 : _GEN_38; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_40 = 6'h25 == stage1_index ? lru_list_37 : _GEN_39; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_41 = 6'h26 == stage1_index ? lru_list_38 : _GEN_40; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_42 = 6'h27 == stage1_index ? lru_list_39 : _GEN_41; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_43 = 6'h28 == stage1_index ? lru_list_40 : _GEN_42; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_44 = 6'h29 == stage1_index ? lru_list_41 : _GEN_43; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_45 = 6'h2a == stage1_index ? lru_list_42 : _GEN_44; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_46 = 6'h2b == stage1_index ? lru_list_43 : _GEN_45; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_47 = 6'h2c == stage1_index ? lru_list_44 : _GEN_46; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_48 = 6'h2d == stage1_index ? lru_list_45 : _GEN_47; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_49 = 6'h2e == stage1_index ? lru_list_46 : _GEN_48; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_50 = 6'h2f == stage1_index ? lru_list_47 : _GEN_49; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_51 = 6'h30 == stage1_index ? lru_list_48 : _GEN_50; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_52 = 6'h31 == stage1_index ? lru_list_49 : _GEN_51; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_53 = 6'h32 == stage1_index ? lru_list_50 : _GEN_52; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_54 = 6'h33 == stage1_index ? lru_list_51 : _GEN_53; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_55 = 6'h34 == stage1_index ? lru_list_52 : _GEN_54; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_56 = 6'h35 == stage1_index ? lru_list_53 : _GEN_55; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_57 = 6'h36 == stage1_index ? lru_list_54 : _GEN_56; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_58 = 6'h37 == stage1_index ? lru_list_55 : _GEN_57; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_59 = 6'h38 == stage1_index ? lru_list_56 : _GEN_58; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_60 = 6'h39 == stage1_index ? lru_list_57 : _GEN_59; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_61 = 6'h3a == stage1_index ? lru_list_58 : _GEN_60; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_62 = 6'h3b == stage1_index ? lru_list_59 : _GEN_61; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_63 = 6'h3c == stage1_index ? lru_list_60 : _GEN_62; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_64 = 6'h3d == stage1_index ? lru_list_61 : _GEN_63; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_65 = 6'h3e == stage1_index ? lru_list_62 : _GEN_64; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  _GEN_66 = 6'h3f == stage1_index ? lru_list_63 : _GEN_65; // @[ICache.scala 124:35 ICache.scala 124:35]
  wire  next_way = ~_GEN_66; // @[ICache.scala 124:35]
  wire [29:0] tag_array_out_0 = io_sram2_rdata[29:0]; // @[ICache.scala 97:50]
  wire [29:0] tag_array_out_1 = io_sram3_rdata[29:0]; // @[ICache.scala 98:50]
  reg  valid_array_0_0; // @[ICache.scala 99:44]
  reg  valid_array_0_1; // @[ICache.scala 99:44]
  reg  valid_array_0_2; // @[ICache.scala 99:44]
  reg  valid_array_0_3; // @[ICache.scala 99:44]
  reg  valid_array_0_4; // @[ICache.scala 99:44]
  reg  valid_array_0_5; // @[ICache.scala 99:44]
  reg  valid_array_0_6; // @[ICache.scala 99:44]
  reg  valid_array_0_7; // @[ICache.scala 99:44]
  reg  valid_array_0_8; // @[ICache.scala 99:44]
  reg  valid_array_0_9; // @[ICache.scala 99:44]
  reg  valid_array_0_10; // @[ICache.scala 99:44]
  reg  valid_array_0_11; // @[ICache.scala 99:44]
  reg  valid_array_0_12; // @[ICache.scala 99:44]
  reg  valid_array_0_13; // @[ICache.scala 99:44]
  reg  valid_array_0_14; // @[ICache.scala 99:44]
  reg  valid_array_0_15; // @[ICache.scala 99:44]
  reg  valid_array_0_16; // @[ICache.scala 99:44]
  reg  valid_array_0_17; // @[ICache.scala 99:44]
  reg  valid_array_0_18; // @[ICache.scala 99:44]
  reg  valid_array_0_19; // @[ICache.scala 99:44]
  reg  valid_array_0_20; // @[ICache.scala 99:44]
  reg  valid_array_0_21; // @[ICache.scala 99:44]
  reg  valid_array_0_22; // @[ICache.scala 99:44]
  reg  valid_array_0_23; // @[ICache.scala 99:44]
  reg  valid_array_0_24; // @[ICache.scala 99:44]
  reg  valid_array_0_25; // @[ICache.scala 99:44]
  reg  valid_array_0_26; // @[ICache.scala 99:44]
  reg  valid_array_0_27; // @[ICache.scala 99:44]
  reg  valid_array_0_28; // @[ICache.scala 99:44]
  reg  valid_array_0_29; // @[ICache.scala 99:44]
  reg  valid_array_0_30; // @[ICache.scala 99:44]
  reg  valid_array_0_31; // @[ICache.scala 99:44]
  reg  valid_array_0_32; // @[ICache.scala 99:44]
  reg  valid_array_0_33; // @[ICache.scala 99:44]
  reg  valid_array_0_34; // @[ICache.scala 99:44]
  reg  valid_array_0_35; // @[ICache.scala 99:44]
  reg  valid_array_0_36; // @[ICache.scala 99:44]
  reg  valid_array_0_37; // @[ICache.scala 99:44]
  reg  valid_array_0_38; // @[ICache.scala 99:44]
  reg  valid_array_0_39; // @[ICache.scala 99:44]
  reg  valid_array_0_40; // @[ICache.scala 99:44]
  reg  valid_array_0_41; // @[ICache.scala 99:44]
  reg  valid_array_0_42; // @[ICache.scala 99:44]
  reg  valid_array_0_43; // @[ICache.scala 99:44]
  reg  valid_array_0_44; // @[ICache.scala 99:44]
  reg  valid_array_0_45; // @[ICache.scala 99:44]
  reg  valid_array_0_46; // @[ICache.scala 99:44]
  reg  valid_array_0_47; // @[ICache.scala 99:44]
  reg  valid_array_0_48; // @[ICache.scala 99:44]
  reg  valid_array_0_49; // @[ICache.scala 99:44]
  reg  valid_array_0_50; // @[ICache.scala 99:44]
  reg  valid_array_0_51; // @[ICache.scala 99:44]
  reg  valid_array_0_52; // @[ICache.scala 99:44]
  reg  valid_array_0_53; // @[ICache.scala 99:44]
  reg  valid_array_0_54; // @[ICache.scala 99:44]
  reg  valid_array_0_55; // @[ICache.scala 99:44]
  reg  valid_array_0_56; // @[ICache.scala 99:44]
  reg  valid_array_0_57; // @[ICache.scala 99:44]
  reg  valid_array_0_58; // @[ICache.scala 99:44]
  reg  valid_array_0_59; // @[ICache.scala 99:44]
  reg  valid_array_0_60; // @[ICache.scala 99:44]
  reg  valid_array_0_61; // @[ICache.scala 99:44]
  reg  valid_array_0_62; // @[ICache.scala 99:44]
  reg  valid_array_0_63; // @[ICache.scala 99:44]
  reg  valid_array_1_0; // @[ICache.scala 100:44]
  reg  valid_array_1_1; // @[ICache.scala 100:44]
  reg  valid_array_1_2; // @[ICache.scala 100:44]
  reg  valid_array_1_3; // @[ICache.scala 100:44]
  reg  valid_array_1_4; // @[ICache.scala 100:44]
  reg  valid_array_1_5; // @[ICache.scala 100:44]
  reg  valid_array_1_6; // @[ICache.scala 100:44]
  reg  valid_array_1_7; // @[ICache.scala 100:44]
  reg  valid_array_1_8; // @[ICache.scala 100:44]
  reg  valid_array_1_9; // @[ICache.scala 100:44]
  reg  valid_array_1_10; // @[ICache.scala 100:44]
  reg  valid_array_1_11; // @[ICache.scala 100:44]
  reg  valid_array_1_12; // @[ICache.scala 100:44]
  reg  valid_array_1_13; // @[ICache.scala 100:44]
  reg  valid_array_1_14; // @[ICache.scala 100:44]
  reg  valid_array_1_15; // @[ICache.scala 100:44]
  reg  valid_array_1_16; // @[ICache.scala 100:44]
  reg  valid_array_1_17; // @[ICache.scala 100:44]
  reg  valid_array_1_18; // @[ICache.scala 100:44]
  reg  valid_array_1_19; // @[ICache.scala 100:44]
  reg  valid_array_1_20; // @[ICache.scala 100:44]
  reg  valid_array_1_21; // @[ICache.scala 100:44]
  reg  valid_array_1_22; // @[ICache.scala 100:44]
  reg  valid_array_1_23; // @[ICache.scala 100:44]
  reg  valid_array_1_24; // @[ICache.scala 100:44]
  reg  valid_array_1_25; // @[ICache.scala 100:44]
  reg  valid_array_1_26; // @[ICache.scala 100:44]
  reg  valid_array_1_27; // @[ICache.scala 100:44]
  reg  valid_array_1_28; // @[ICache.scala 100:44]
  reg  valid_array_1_29; // @[ICache.scala 100:44]
  reg  valid_array_1_30; // @[ICache.scala 100:44]
  reg  valid_array_1_31; // @[ICache.scala 100:44]
  reg  valid_array_1_32; // @[ICache.scala 100:44]
  reg  valid_array_1_33; // @[ICache.scala 100:44]
  reg  valid_array_1_34; // @[ICache.scala 100:44]
  reg  valid_array_1_35; // @[ICache.scala 100:44]
  reg  valid_array_1_36; // @[ICache.scala 100:44]
  reg  valid_array_1_37; // @[ICache.scala 100:44]
  reg  valid_array_1_38; // @[ICache.scala 100:44]
  reg  valid_array_1_39; // @[ICache.scala 100:44]
  reg  valid_array_1_40; // @[ICache.scala 100:44]
  reg  valid_array_1_41; // @[ICache.scala 100:44]
  reg  valid_array_1_42; // @[ICache.scala 100:44]
  reg  valid_array_1_43; // @[ICache.scala 100:44]
  reg  valid_array_1_44; // @[ICache.scala 100:44]
  reg  valid_array_1_45; // @[ICache.scala 100:44]
  reg  valid_array_1_46; // @[ICache.scala 100:44]
  reg  valid_array_1_47; // @[ICache.scala 100:44]
  reg  valid_array_1_48; // @[ICache.scala 100:44]
  reg  valid_array_1_49; // @[ICache.scala 100:44]
  reg  valid_array_1_50; // @[ICache.scala 100:44]
  reg  valid_array_1_51; // @[ICache.scala 100:44]
  reg  valid_array_1_52; // @[ICache.scala 100:44]
  reg  valid_array_1_53; // @[ICache.scala 100:44]
  reg  valid_array_1_54; // @[ICache.scala 100:44]
  reg  valid_array_1_55; // @[ICache.scala 100:44]
  reg  valid_array_1_56; // @[ICache.scala 100:44]
  reg  valid_array_1_57; // @[ICache.scala 100:44]
  reg  valid_array_1_58; // @[ICache.scala 100:44]
  reg  valid_array_1_59; // @[ICache.scala 100:44]
  reg  valid_array_1_60; // @[ICache.scala 100:44]
  reg  valid_array_1_61; // @[ICache.scala 100:44]
  reg  valid_array_1_62; // @[ICache.scala 100:44]
  reg  valid_array_1_63; // @[ICache.scala 100:44]
  reg  stage1_out_valid; // @[Reg.scala 27:20]
  wire  _T_4 = 3'h0 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1208 = io_next_ready & io_prev_valid ? 3'h2 : curr_state; // @[ICache.scala 206:36 ICache.scala 206:49 ICache.scala 203:14]
  wire  _T_6 = 3'h1 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1209 = maxi4_manager_io_out_finish ? 3'h0 : curr_state; // @[ICache.scala 210:31 ICache.scala 210:44 ICache.scala 203:14]
  wire [2:0] _GEN_1210 = maxi4_manager_io_out_finish & io_next_ready ? 3'h2 : _GEN_1209; // @[ICache.scala 209:37 ICache.scala 209:50]
  wire  _T_8 = 3'h2 == curr_state; // @[Conditional.scala 37:30]
  wire  addr_underflow = ~stage1_out_bits_addr[31]; // @[ICache.scala 128:60]
  wire [2:0] _GEN_1211 = maxi4_manager_io_out_ready ? 3'h7 : 3'h6; // @[ICache.scala 218:25 ICache.scala 218:38 ICache.scala 219:38]
  wire [28:0] stage1_tag = stage1_out_bits_addr[38:10]; // @[ICache.scala 118:54]
  wire [29:0] _GEN_1235 = {{1'd0}, stage1_tag}; // @[ICache.scala 125:52]
  wire  _GEN_74 = 6'h1 == stage1_index ? valid_array_0_1 : valid_array_0_0; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_75 = 6'h2 == stage1_index ? valid_array_0_2 : _GEN_74; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_76 = 6'h3 == stage1_index ? valid_array_0_3 : _GEN_75; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_77 = 6'h4 == stage1_index ? valid_array_0_4 : _GEN_76; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_78 = 6'h5 == stage1_index ? valid_array_0_5 : _GEN_77; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_79 = 6'h6 == stage1_index ? valid_array_0_6 : _GEN_78; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_80 = 6'h7 == stage1_index ? valid_array_0_7 : _GEN_79; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_81 = 6'h8 == stage1_index ? valid_array_0_8 : _GEN_80; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_82 = 6'h9 == stage1_index ? valid_array_0_9 : _GEN_81; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_83 = 6'ha == stage1_index ? valid_array_0_10 : _GEN_82; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_84 = 6'hb == stage1_index ? valid_array_0_11 : _GEN_83; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_85 = 6'hc == stage1_index ? valid_array_0_12 : _GEN_84; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_86 = 6'hd == stage1_index ? valid_array_0_13 : _GEN_85; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_87 = 6'he == stage1_index ? valid_array_0_14 : _GEN_86; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_88 = 6'hf == stage1_index ? valid_array_0_15 : _GEN_87; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_89 = 6'h10 == stage1_index ? valid_array_0_16 : _GEN_88; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_90 = 6'h11 == stage1_index ? valid_array_0_17 : _GEN_89; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_91 = 6'h12 == stage1_index ? valid_array_0_18 : _GEN_90; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_92 = 6'h13 == stage1_index ? valid_array_0_19 : _GEN_91; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_93 = 6'h14 == stage1_index ? valid_array_0_20 : _GEN_92; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_94 = 6'h15 == stage1_index ? valid_array_0_21 : _GEN_93; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_95 = 6'h16 == stage1_index ? valid_array_0_22 : _GEN_94; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_96 = 6'h17 == stage1_index ? valid_array_0_23 : _GEN_95; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_97 = 6'h18 == stage1_index ? valid_array_0_24 : _GEN_96; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_98 = 6'h19 == stage1_index ? valid_array_0_25 : _GEN_97; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_99 = 6'h1a == stage1_index ? valid_array_0_26 : _GEN_98; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_100 = 6'h1b == stage1_index ? valid_array_0_27 : _GEN_99; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_101 = 6'h1c == stage1_index ? valid_array_0_28 : _GEN_100; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_102 = 6'h1d == stage1_index ? valid_array_0_29 : _GEN_101; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_103 = 6'h1e == stage1_index ? valid_array_0_30 : _GEN_102; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_104 = 6'h1f == stage1_index ? valid_array_0_31 : _GEN_103; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_105 = 6'h20 == stage1_index ? valid_array_0_32 : _GEN_104; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_106 = 6'h21 == stage1_index ? valid_array_0_33 : _GEN_105; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_107 = 6'h22 == stage1_index ? valid_array_0_34 : _GEN_106; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_108 = 6'h23 == stage1_index ? valid_array_0_35 : _GEN_107; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_109 = 6'h24 == stage1_index ? valid_array_0_36 : _GEN_108; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_110 = 6'h25 == stage1_index ? valid_array_0_37 : _GEN_109; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_111 = 6'h26 == stage1_index ? valid_array_0_38 : _GEN_110; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_112 = 6'h27 == stage1_index ? valid_array_0_39 : _GEN_111; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_113 = 6'h28 == stage1_index ? valid_array_0_40 : _GEN_112; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_114 = 6'h29 == stage1_index ? valid_array_0_41 : _GEN_113; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_115 = 6'h2a == stage1_index ? valid_array_0_42 : _GEN_114; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_116 = 6'h2b == stage1_index ? valid_array_0_43 : _GEN_115; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_117 = 6'h2c == stage1_index ? valid_array_0_44 : _GEN_116; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_118 = 6'h2d == stage1_index ? valid_array_0_45 : _GEN_117; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_119 = 6'h2e == stage1_index ? valid_array_0_46 : _GEN_118; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_120 = 6'h2f == stage1_index ? valid_array_0_47 : _GEN_119; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_121 = 6'h30 == stage1_index ? valid_array_0_48 : _GEN_120; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_122 = 6'h31 == stage1_index ? valid_array_0_49 : _GEN_121; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_123 = 6'h32 == stage1_index ? valid_array_0_50 : _GEN_122; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_124 = 6'h33 == stage1_index ? valid_array_0_51 : _GEN_123; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_125 = 6'h34 == stage1_index ? valid_array_0_52 : _GEN_124; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_126 = 6'h35 == stage1_index ? valid_array_0_53 : _GEN_125; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_127 = 6'h36 == stage1_index ? valid_array_0_54 : _GEN_126; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_128 = 6'h37 == stage1_index ? valid_array_0_55 : _GEN_127; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_129 = 6'h38 == stage1_index ? valid_array_0_56 : _GEN_128; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_130 = 6'h39 == stage1_index ? valid_array_0_57 : _GEN_129; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_131 = 6'h3a == stage1_index ? valid_array_0_58 : _GEN_130; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_132 = 6'h3b == stage1_index ? valid_array_0_59 : _GEN_131; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_133 = 6'h3c == stage1_index ? valid_array_0_60 : _GEN_132; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_134 = 6'h3d == stage1_index ? valid_array_0_61 : _GEN_133; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_135 = 6'h3e == stage1_index ? valid_array_0_62 : _GEN_134; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  _GEN_136 = 6'h3f == stage1_index ? valid_array_0_63 : _GEN_135; // @[ICache.scala 171:21 ICache.scala 171:21]
  wire  valid_array_0_out = fencei ? 1'h0 : _GEN_136; // @[ICache.scala 189:26 ICache.scala 192:23 ICache.scala 171:21]
  wire  tag0_hit = tag_array_out_0 == _GEN_1235 & valid_array_0_out; // @[ICache.scala 125:68]
  wire  _GEN_138 = 6'h1 == stage1_index ? valid_array_1_1 : valid_array_1_0; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_139 = 6'h2 == stage1_index ? valid_array_1_2 : _GEN_138; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_140 = 6'h3 == stage1_index ? valid_array_1_3 : _GEN_139; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_141 = 6'h4 == stage1_index ? valid_array_1_4 : _GEN_140; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_142 = 6'h5 == stage1_index ? valid_array_1_5 : _GEN_141; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_143 = 6'h6 == stage1_index ? valid_array_1_6 : _GEN_142; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_144 = 6'h7 == stage1_index ? valid_array_1_7 : _GEN_143; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_145 = 6'h8 == stage1_index ? valid_array_1_8 : _GEN_144; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_146 = 6'h9 == stage1_index ? valid_array_1_9 : _GEN_145; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_147 = 6'ha == stage1_index ? valid_array_1_10 : _GEN_146; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_148 = 6'hb == stage1_index ? valid_array_1_11 : _GEN_147; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_149 = 6'hc == stage1_index ? valid_array_1_12 : _GEN_148; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_150 = 6'hd == stage1_index ? valid_array_1_13 : _GEN_149; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_151 = 6'he == stage1_index ? valid_array_1_14 : _GEN_150; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_152 = 6'hf == stage1_index ? valid_array_1_15 : _GEN_151; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_153 = 6'h10 == stage1_index ? valid_array_1_16 : _GEN_152; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_154 = 6'h11 == stage1_index ? valid_array_1_17 : _GEN_153; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_155 = 6'h12 == stage1_index ? valid_array_1_18 : _GEN_154; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_156 = 6'h13 == stage1_index ? valid_array_1_19 : _GEN_155; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_157 = 6'h14 == stage1_index ? valid_array_1_20 : _GEN_156; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_158 = 6'h15 == stage1_index ? valid_array_1_21 : _GEN_157; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_159 = 6'h16 == stage1_index ? valid_array_1_22 : _GEN_158; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_160 = 6'h17 == stage1_index ? valid_array_1_23 : _GEN_159; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_161 = 6'h18 == stage1_index ? valid_array_1_24 : _GEN_160; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_162 = 6'h19 == stage1_index ? valid_array_1_25 : _GEN_161; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_163 = 6'h1a == stage1_index ? valid_array_1_26 : _GEN_162; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_164 = 6'h1b == stage1_index ? valid_array_1_27 : _GEN_163; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_165 = 6'h1c == stage1_index ? valid_array_1_28 : _GEN_164; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_166 = 6'h1d == stage1_index ? valid_array_1_29 : _GEN_165; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_167 = 6'h1e == stage1_index ? valid_array_1_30 : _GEN_166; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_168 = 6'h1f == stage1_index ? valid_array_1_31 : _GEN_167; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_169 = 6'h20 == stage1_index ? valid_array_1_32 : _GEN_168; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_170 = 6'h21 == stage1_index ? valid_array_1_33 : _GEN_169; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_171 = 6'h22 == stage1_index ? valid_array_1_34 : _GEN_170; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_172 = 6'h23 == stage1_index ? valid_array_1_35 : _GEN_171; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_173 = 6'h24 == stage1_index ? valid_array_1_36 : _GEN_172; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_174 = 6'h25 == stage1_index ? valid_array_1_37 : _GEN_173; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_175 = 6'h26 == stage1_index ? valid_array_1_38 : _GEN_174; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_176 = 6'h27 == stage1_index ? valid_array_1_39 : _GEN_175; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_177 = 6'h28 == stage1_index ? valid_array_1_40 : _GEN_176; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_178 = 6'h29 == stage1_index ? valid_array_1_41 : _GEN_177; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_179 = 6'h2a == stage1_index ? valid_array_1_42 : _GEN_178; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_180 = 6'h2b == stage1_index ? valid_array_1_43 : _GEN_179; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_181 = 6'h2c == stage1_index ? valid_array_1_44 : _GEN_180; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_182 = 6'h2d == stage1_index ? valid_array_1_45 : _GEN_181; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_183 = 6'h2e == stage1_index ? valid_array_1_46 : _GEN_182; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_184 = 6'h2f == stage1_index ? valid_array_1_47 : _GEN_183; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_185 = 6'h30 == stage1_index ? valid_array_1_48 : _GEN_184; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_186 = 6'h31 == stage1_index ? valid_array_1_49 : _GEN_185; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_187 = 6'h32 == stage1_index ? valid_array_1_50 : _GEN_186; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_188 = 6'h33 == stage1_index ? valid_array_1_51 : _GEN_187; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_189 = 6'h34 == stage1_index ? valid_array_1_52 : _GEN_188; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_190 = 6'h35 == stage1_index ? valid_array_1_53 : _GEN_189; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_191 = 6'h36 == stage1_index ? valid_array_1_54 : _GEN_190; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_192 = 6'h37 == stage1_index ? valid_array_1_55 : _GEN_191; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_193 = 6'h38 == stage1_index ? valid_array_1_56 : _GEN_192; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_194 = 6'h39 == stage1_index ? valid_array_1_57 : _GEN_193; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_195 = 6'h3a == stage1_index ? valid_array_1_58 : _GEN_194; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_196 = 6'h3b == stage1_index ? valid_array_1_59 : _GEN_195; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_197 = 6'h3c == stage1_index ? valid_array_1_60 : _GEN_196; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_198 = 6'h3d == stage1_index ? valid_array_1_61 : _GEN_197; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_199 = 6'h3e == stage1_index ? valid_array_1_62 : _GEN_198; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  _GEN_200 = 6'h3f == stage1_index ? valid_array_1_63 : _GEN_199; // @[ICache.scala 172:21 ICache.scala 172:21]
  wire  valid_array_1_out = fencei ? 1'h0 : _GEN_200; // @[ICache.scala 189:26 ICache.scala 193:23 ICache.scala 172:21]
  wire  tag1_hit = tag_array_out_1 == _GEN_1235 & valid_array_1_out; // @[ICache.scala 126:68]
  wire  miss = ~(tag0_hit | tag1_hit); // @[ICache.scala 127:35]
  wire [2:0] _GEN_1212 = maxi4_manager_io_out_ready ? 3'h4 : 3'h3; // @[ICache.scala 221:25 ICache.scala 221:38 ICache.scala 222:38]
  wire [2:0] _GEN_1213 = miss ? _GEN_1212 : curr_state; // @[ICache.scala 220:24 ICache.scala 203:14]
  wire [2:0] _GEN_1214 = addr_underflow ? _GEN_1211 : _GEN_1213; // @[ICache.scala 217:33]
  wire [2:0] _GEN_1215 = ~io_prev_valid ? 3'h2 : _GEN_1214; // @[ICache.scala 215:30 ICache.scala 216:20]
  wire [2:0] _GEN_1216 = io_cache_reset ? 3'h2 : _GEN_1215; // @[ICache.scala 213:24 ICache.scala 214:20]
  wire  _T_10 = 3'h3 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1217 = maxi4_manager_io_out_ready ? 3'h4 : curr_state; // @[ICache.scala 228:30 ICache.scala 229:20 ICache.scala 203:14]
  wire [2:0] _GEN_1218 = io_cache_reset ? 3'h2 : _GEN_1217; // @[ICache.scala 226:24 ICache.scala 227:20]
  wire  _T_11 = 3'h4 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1219 = maxi4_manager_io_out_finish ? 3'h5 : curr_state; // @[ICache.scala 237:30 ICache.scala 238:20 ICache.scala 203:14]
  wire [2:0] _GEN_1220 = io_cache_reset ? 3'h1 : _GEN_1219; // @[ICache.scala 235:30 ICache.scala 236:20]
  wire [2:0] _GEN_1221 = io_cache_reset & maxi4_manager_io_out_finish ? 3'h2 : _GEN_1220; // @[ICache.scala 233:38 ICache.scala 234:20]
  wire  _T_13 = 3'h6 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1222 = maxi4_manager_io_out_ready ? 3'h7 : curr_state; // @[ICache.scala 244:30 ICache.scala 245:20 ICache.scala 203:14]
  wire [2:0] _GEN_1223 = io_cache_reset ? 3'h2 : _GEN_1222; // @[ICache.scala 242:24 ICache.scala 243:20]
  wire  _T_14 = 3'h7 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h5 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_1225 = io_next_ready ? 3'h2 : curr_state; // @[ICache.scala 260:29 ICache.scala 261:20 ICache.scala 263:20]
  wire [2:0] _GEN_1226 = io_cache_reset ? 3'h2 : _GEN_1225; // @[ICache.scala 258:24 ICache.scala 259:20]
  wire [2:0] _GEN_1227 = _T_16 ? _GEN_1226 : curr_state; // @[Conditional.scala 39:67 ICache.scala 203:14]
  wire [2:0] _GEN_1228 = _T_14 ? _GEN_1221 : _GEN_1227; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1229 = _T_13 ? _GEN_1223 : _GEN_1228; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1230 = _T_11 ? _GEN_1221 : _GEN_1229; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1231 = _T_10 ? _GEN_1218 : _GEN_1230; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1232 = _T_8 ? _GEN_1216 : _GEN_1231; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_1233 = _T_6 ? _GEN_1210 : _GEN_1232; // @[Conditional.scala 39:67]
  wire [2:0] next_state = _T_4 ? _GEN_1208 : _GEN_1233; // @[Conditional.scala 40:58]
  wire  go_on = next_state == 3'h2 & io_next_ready | io_cache_reset; // @[ICache.scala 129:73]
  wire [5:0] prev_index = io_prev_bits_addr[9:4]; // @[ICache.scala 115:48]
  wire [127:0] _cache_line_data_out_T = tag1_hit ? io_sram1_rdata : 128'h0; // @[Mux.scala 98:16]
  wire [127:0] cache_line_data_out = tag0_hit ? io_sram0_rdata : _cache_line_data_out_T; // @[Mux.scala 98:16]
  wire  _T = curr_state == 3'h2; // @[ICache.scala 151:25]
  wire  _GEN_68 = addr_underflow | miss; // @[ICache.scala 152:26 ICache.scala 153:18]
  wire  _T_2 = curr_state == 3'h6; // @[ICache.scala 159:25]
  wire  _GEN_70 = curr_state == 3'h3 | _T_2; // @[ICache.scala 157:36 ICache.scala 158:16]
  wire  _GEN_71 = curr_state == 3'h2 ? _GEN_68 : _GEN_70; // @[ICache.scala 151:37]
  wire [34:0] maxi4_manager_io_in_addr_hi = stage1_out_bits_addr[38:4]; // @[ICache.scala 162:93]
  wire [38:0] _maxi4_manager_io_in_addr_T_1 = {maxi4_manager_io_in_addr_hi,4'h0}; // @[Cat.scala 30:58]
  wire [38:0] _maxi4_manager_io_in_addr_T_2 = addr_underflow ? stage1_out_bits_addr : _maxi4_manager_io_in_addr_T_1; // @[ICache.scala 162:18]
  wire  _GEN_1237 = 6'h0 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_201 = 6'h0 == stage1_index | lru_list_0; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1238 = 6'h1 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_202 = 6'h1 == stage1_index | lru_list_1; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1239 = 6'h2 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_203 = 6'h2 == stage1_index | lru_list_2; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1240 = 6'h3 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_204 = 6'h3 == stage1_index | lru_list_3; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1241 = 6'h4 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_205 = 6'h4 == stage1_index | lru_list_4; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1242 = 6'h5 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_206 = 6'h5 == stage1_index | lru_list_5; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1243 = 6'h6 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_207 = 6'h6 == stage1_index | lru_list_6; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1244 = 6'h7 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_208 = 6'h7 == stage1_index | lru_list_7; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1245 = 6'h8 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_209 = 6'h8 == stage1_index | lru_list_8; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1246 = 6'h9 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_210 = 6'h9 == stage1_index | lru_list_9; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1247 = 6'ha == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_211 = 6'ha == stage1_index | lru_list_10; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1248 = 6'hb == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_212 = 6'hb == stage1_index | lru_list_11; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1249 = 6'hc == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_213 = 6'hc == stage1_index | lru_list_12; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1250 = 6'hd == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_214 = 6'hd == stage1_index | lru_list_13; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1251 = 6'he == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_215 = 6'he == stage1_index | lru_list_14; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1252 = 6'hf == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_216 = 6'hf == stage1_index | lru_list_15; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1253 = 6'h10 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_217 = 6'h10 == stage1_index | lru_list_16; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1254 = 6'h11 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_218 = 6'h11 == stage1_index | lru_list_17; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1255 = 6'h12 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_219 = 6'h12 == stage1_index | lru_list_18; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1256 = 6'h13 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_220 = 6'h13 == stage1_index | lru_list_19; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1257 = 6'h14 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_221 = 6'h14 == stage1_index | lru_list_20; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1258 = 6'h15 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_222 = 6'h15 == stage1_index | lru_list_21; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1259 = 6'h16 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_223 = 6'h16 == stage1_index | lru_list_22; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1260 = 6'h17 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_224 = 6'h17 == stage1_index | lru_list_23; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1261 = 6'h18 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_225 = 6'h18 == stage1_index | lru_list_24; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1262 = 6'h19 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_226 = 6'h19 == stage1_index | lru_list_25; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1263 = 6'h1a == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_227 = 6'h1a == stage1_index | lru_list_26; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1264 = 6'h1b == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_228 = 6'h1b == stage1_index | lru_list_27; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1265 = 6'h1c == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_229 = 6'h1c == stage1_index | lru_list_28; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1266 = 6'h1d == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_230 = 6'h1d == stage1_index | lru_list_29; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1267 = 6'h1e == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_231 = 6'h1e == stage1_index | lru_list_30; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1268 = 6'h1f == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_232 = 6'h1f == stage1_index | lru_list_31; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1269 = 6'h20 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_233 = 6'h20 == stage1_index | lru_list_32; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1270 = 6'h21 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_234 = 6'h21 == stage1_index | lru_list_33; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1271 = 6'h22 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_235 = 6'h22 == stage1_index | lru_list_34; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1272 = 6'h23 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_236 = 6'h23 == stage1_index | lru_list_35; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1273 = 6'h24 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_237 = 6'h24 == stage1_index | lru_list_36; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1274 = 6'h25 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_238 = 6'h25 == stage1_index | lru_list_37; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1275 = 6'h26 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_239 = 6'h26 == stage1_index | lru_list_38; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1276 = 6'h27 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_240 = 6'h27 == stage1_index | lru_list_39; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1277 = 6'h28 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_241 = 6'h28 == stage1_index | lru_list_40; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1278 = 6'h29 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_242 = 6'h29 == stage1_index | lru_list_41; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1279 = 6'h2a == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_243 = 6'h2a == stage1_index | lru_list_42; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1280 = 6'h2b == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_244 = 6'h2b == stage1_index | lru_list_43; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1281 = 6'h2c == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_245 = 6'h2c == stage1_index | lru_list_44; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1282 = 6'h2d == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_246 = 6'h2d == stage1_index | lru_list_45; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1283 = 6'h2e == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_247 = 6'h2e == stage1_index | lru_list_46; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1284 = 6'h2f == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_248 = 6'h2f == stage1_index | lru_list_47; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1285 = 6'h30 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_249 = 6'h30 == stage1_index | lru_list_48; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1286 = 6'h31 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_250 = 6'h31 == stage1_index | lru_list_49; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1287 = 6'h32 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_251 = 6'h32 == stage1_index | lru_list_50; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1288 = 6'h33 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_252 = 6'h33 == stage1_index | lru_list_51; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1289 = 6'h34 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_253 = 6'h34 == stage1_index | lru_list_52; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1290 = 6'h35 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_254 = 6'h35 == stage1_index | lru_list_53; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1291 = 6'h36 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_255 = 6'h36 == stage1_index | lru_list_54; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1292 = 6'h37 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_256 = 6'h37 == stage1_index | lru_list_55; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1293 = 6'h38 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_257 = 6'h38 == stage1_index | lru_list_56; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1294 = 6'h39 == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_258 = 6'h39 == stage1_index | lru_list_57; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1295 = 6'h3a == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_259 = 6'h3a == stage1_index | lru_list_58; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1296 = 6'h3b == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_260 = 6'h3b == stage1_index | lru_list_59; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1297 = 6'h3c == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_261 = 6'h3c == stage1_index | lru_list_60; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1298 = 6'h3d == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_262 = 6'h3d == stage1_index | lru_list_61; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1299 = 6'h3e == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_263 = 6'h3e == stage1_index | lru_list_62; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_1300 = 6'h3f == stage1_index; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_264 = 6'h3f == stage1_index | lru_list_63; // @[ICache.scala 176:34 ICache.scala 176:34 ICache.scala 103:35]
  wire  _GEN_265 = _GEN_1237 | valid_array_1_0; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_266 = _GEN_1238 | valid_array_1_1; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_267 = _GEN_1239 | valid_array_1_2; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_268 = _GEN_1240 | valid_array_1_3; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_269 = _GEN_1241 | valid_array_1_4; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_270 = _GEN_1242 | valid_array_1_5; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_271 = _GEN_1243 | valid_array_1_6; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_272 = _GEN_1244 | valid_array_1_7; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_273 = _GEN_1245 | valid_array_1_8; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_274 = _GEN_1246 | valid_array_1_9; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_275 = _GEN_1247 | valid_array_1_10; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_276 = _GEN_1248 | valid_array_1_11; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_277 = _GEN_1249 | valid_array_1_12; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_278 = _GEN_1250 | valid_array_1_13; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_279 = _GEN_1251 | valid_array_1_14; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_280 = _GEN_1252 | valid_array_1_15; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_281 = _GEN_1253 | valid_array_1_16; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_282 = _GEN_1254 | valid_array_1_17; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_283 = _GEN_1255 | valid_array_1_18; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_284 = _GEN_1256 | valid_array_1_19; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_285 = _GEN_1257 | valid_array_1_20; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_286 = _GEN_1258 | valid_array_1_21; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_287 = _GEN_1259 | valid_array_1_22; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_288 = _GEN_1260 | valid_array_1_23; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_289 = _GEN_1261 | valid_array_1_24; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_290 = _GEN_1262 | valid_array_1_25; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_291 = _GEN_1263 | valid_array_1_26; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_292 = _GEN_1264 | valid_array_1_27; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_293 = _GEN_1265 | valid_array_1_28; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_294 = _GEN_1266 | valid_array_1_29; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_295 = _GEN_1267 | valid_array_1_30; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_296 = _GEN_1268 | valid_array_1_31; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_297 = _GEN_1269 | valid_array_1_32; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_298 = _GEN_1270 | valid_array_1_33; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_299 = _GEN_1271 | valid_array_1_34; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_300 = _GEN_1272 | valid_array_1_35; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_301 = _GEN_1273 | valid_array_1_36; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_302 = _GEN_1274 | valid_array_1_37; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_303 = _GEN_1275 | valid_array_1_38; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_304 = _GEN_1276 | valid_array_1_39; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_305 = _GEN_1277 | valid_array_1_40; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_306 = _GEN_1278 | valid_array_1_41; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_307 = _GEN_1279 | valid_array_1_42; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_308 = _GEN_1280 | valid_array_1_43; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_309 = _GEN_1281 | valid_array_1_44; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_310 = _GEN_1282 | valid_array_1_45; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_311 = _GEN_1283 | valid_array_1_46; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_312 = _GEN_1284 | valid_array_1_47; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_313 = _GEN_1285 | valid_array_1_48; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_314 = _GEN_1286 | valid_array_1_49; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_315 = _GEN_1287 | valid_array_1_50; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_316 = _GEN_1288 | valid_array_1_51; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_317 = _GEN_1289 | valid_array_1_52; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_318 = _GEN_1290 | valid_array_1_53; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_319 = _GEN_1291 | valid_array_1_54; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_320 = _GEN_1292 | valid_array_1_55; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_321 = _GEN_1293 | valid_array_1_56; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_322 = _GEN_1294 | valid_array_1_57; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_323 = _GEN_1295 | valid_array_1_58; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_324 = _GEN_1296 | valid_array_1_59; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_325 = _GEN_1297 | valid_array_1_60; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_326 = _GEN_1298 | valid_array_1_61; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_327 = _GEN_1299 | valid_array_1_62; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_328 = _GEN_1300 | valid_array_1_63; // @[ICache.scala 179:39 ICache.scala 179:39 ICache.scala 100:44]
  wire  _GEN_329 = 6'h0 == stage1_index ? 1'h0 : lru_list_0; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_330 = 6'h1 == stage1_index ? 1'h0 : lru_list_1; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_331 = 6'h2 == stage1_index ? 1'h0 : lru_list_2; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_332 = 6'h3 == stage1_index ? 1'h0 : lru_list_3; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_333 = 6'h4 == stage1_index ? 1'h0 : lru_list_4; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_334 = 6'h5 == stage1_index ? 1'h0 : lru_list_5; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_335 = 6'h6 == stage1_index ? 1'h0 : lru_list_6; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_336 = 6'h7 == stage1_index ? 1'h0 : lru_list_7; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_337 = 6'h8 == stage1_index ? 1'h0 : lru_list_8; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_338 = 6'h9 == stage1_index ? 1'h0 : lru_list_9; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_339 = 6'ha == stage1_index ? 1'h0 : lru_list_10; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_340 = 6'hb == stage1_index ? 1'h0 : lru_list_11; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_341 = 6'hc == stage1_index ? 1'h0 : lru_list_12; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_342 = 6'hd == stage1_index ? 1'h0 : lru_list_13; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_343 = 6'he == stage1_index ? 1'h0 : lru_list_14; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_344 = 6'hf == stage1_index ? 1'h0 : lru_list_15; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_345 = 6'h10 == stage1_index ? 1'h0 : lru_list_16; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_346 = 6'h11 == stage1_index ? 1'h0 : lru_list_17; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_347 = 6'h12 == stage1_index ? 1'h0 : lru_list_18; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_348 = 6'h13 == stage1_index ? 1'h0 : lru_list_19; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_349 = 6'h14 == stage1_index ? 1'h0 : lru_list_20; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_350 = 6'h15 == stage1_index ? 1'h0 : lru_list_21; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_351 = 6'h16 == stage1_index ? 1'h0 : lru_list_22; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_352 = 6'h17 == stage1_index ? 1'h0 : lru_list_23; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_353 = 6'h18 == stage1_index ? 1'h0 : lru_list_24; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_354 = 6'h19 == stage1_index ? 1'h0 : lru_list_25; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_355 = 6'h1a == stage1_index ? 1'h0 : lru_list_26; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_356 = 6'h1b == stage1_index ? 1'h0 : lru_list_27; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_357 = 6'h1c == stage1_index ? 1'h0 : lru_list_28; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_358 = 6'h1d == stage1_index ? 1'h0 : lru_list_29; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_359 = 6'h1e == stage1_index ? 1'h0 : lru_list_30; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_360 = 6'h1f == stage1_index ? 1'h0 : lru_list_31; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_361 = 6'h20 == stage1_index ? 1'h0 : lru_list_32; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_362 = 6'h21 == stage1_index ? 1'h0 : lru_list_33; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_363 = 6'h22 == stage1_index ? 1'h0 : lru_list_34; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_364 = 6'h23 == stage1_index ? 1'h0 : lru_list_35; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_365 = 6'h24 == stage1_index ? 1'h0 : lru_list_36; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_366 = 6'h25 == stage1_index ? 1'h0 : lru_list_37; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_367 = 6'h26 == stage1_index ? 1'h0 : lru_list_38; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_368 = 6'h27 == stage1_index ? 1'h0 : lru_list_39; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_369 = 6'h28 == stage1_index ? 1'h0 : lru_list_40; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_370 = 6'h29 == stage1_index ? 1'h0 : lru_list_41; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_371 = 6'h2a == stage1_index ? 1'h0 : lru_list_42; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_372 = 6'h2b == stage1_index ? 1'h0 : lru_list_43; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_373 = 6'h2c == stage1_index ? 1'h0 : lru_list_44; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_374 = 6'h2d == stage1_index ? 1'h0 : lru_list_45; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_375 = 6'h2e == stage1_index ? 1'h0 : lru_list_46; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_376 = 6'h2f == stage1_index ? 1'h0 : lru_list_47; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_377 = 6'h30 == stage1_index ? 1'h0 : lru_list_48; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_378 = 6'h31 == stage1_index ? 1'h0 : lru_list_49; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_379 = 6'h32 == stage1_index ? 1'h0 : lru_list_50; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_380 = 6'h33 == stage1_index ? 1'h0 : lru_list_51; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_381 = 6'h34 == stage1_index ? 1'h0 : lru_list_52; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_382 = 6'h35 == stage1_index ? 1'h0 : lru_list_53; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_383 = 6'h36 == stage1_index ? 1'h0 : lru_list_54; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_384 = 6'h37 == stage1_index ? 1'h0 : lru_list_55; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_385 = 6'h38 == stage1_index ? 1'h0 : lru_list_56; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_386 = 6'h39 == stage1_index ? 1'h0 : lru_list_57; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_387 = 6'h3a == stage1_index ? 1'h0 : lru_list_58; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_388 = 6'h3b == stage1_index ? 1'h0 : lru_list_59; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_389 = 6'h3c == stage1_index ? 1'h0 : lru_list_60; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_390 = 6'h3d == stage1_index ? 1'h0 : lru_list_61; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_391 = 6'h3e == stage1_index ? 1'h0 : lru_list_62; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_392 = 6'h3f == stage1_index ? 1'h0 : lru_list_63; // @[ICache.scala 181:34 ICache.scala 181:34 ICache.scala 103:35]
  wire  _GEN_393 = _GEN_1237 | valid_array_0_0; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_394 = _GEN_1238 | valid_array_0_1; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_395 = _GEN_1239 | valid_array_0_2; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_396 = _GEN_1240 | valid_array_0_3; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_397 = _GEN_1241 | valid_array_0_4; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_398 = _GEN_1242 | valid_array_0_5; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_399 = _GEN_1243 | valid_array_0_6; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_400 = _GEN_1244 | valid_array_0_7; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_401 = _GEN_1245 | valid_array_0_8; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_402 = _GEN_1246 | valid_array_0_9; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_403 = _GEN_1247 | valid_array_0_10; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_404 = _GEN_1248 | valid_array_0_11; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_405 = _GEN_1249 | valid_array_0_12; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_406 = _GEN_1250 | valid_array_0_13; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_407 = _GEN_1251 | valid_array_0_14; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_408 = _GEN_1252 | valid_array_0_15; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_409 = _GEN_1253 | valid_array_0_16; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_410 = _GEN_1254 | valid_array_0_17; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_411 = _GEN_1255 | valid_array_0_18; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_412 = _GEN_1256 | valid_array_0_19; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_413 = _GEN_1257 | valid_array_0_20; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_414 = _GEN_1258 | valid_array_0_21; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_415 = _GEN_1259 | valid_array_0_22; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_416 = _GEN_1260 | valid_array_0_23; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_417 = _GEN_1261 | valid_array_0_24; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_418 = _GEN_1262 | valid_array_0_25; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_419 = _GEN_1263 | valid_array_0_26; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_420 = _GEN_1264 | valid_array_0_27; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_421 = _GEN_1265 | valid_array_0_28; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_422 = _GEN_1266 | valid_array_0_29; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_423 = _GEN_1267 | valid_array_0_30; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_424 = _GEN_1268 | valid_array_0_31; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_425 = _GEN_1269 | valid_array_0_32; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_426 = _GEN_1270 | valid_array_0_33; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_427 = _GEN_1271 | valid_array_0_34; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_428 = _GEN_1272 | valid_array_0_35; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_429 = _GEN_1273 | valid_array_0_36; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_430 = _GEN_1274 | valid_array_0_37; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_431 = _GEN_1275 | valid_array_0_38; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_432 = _GEN_1276 | valid_array_0_39; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_433 = _GEN_1277 | valid_array_0_40; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_434 = _GEN_1278 | valid_array_0_41; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_435 = _GEN_1279 | valid_array_0_42; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_436 = _GEN_1280 | valid_array_0_43; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_437 = _GEN_1281 | valid_array_0_44; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_438 = _GEN_1282 | valid_array_0_45; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_439 = _GEN_1283 | valid_array_0_46; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_440 = _GEN_1284 | valid_array_0_47; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_441 = _GEN_1285 | valid_array_0_48; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_442 = _GEN_1286 | valid_array_0_49; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_443 = _GEN_1287 | valid_array_0_50; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_444 = _GEN_1288 | valid_array_0_51; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_445 = _GEN_1289 | valid_array_0_52; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_446 = _GEN_1290 | valid_array_0_53; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_447 = _GEN_1291 | valid_array_0_54; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_448 = _GEN_1292 | valid_array_0_55; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_449 = _GEN_1293 | valid_array_0_56; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_450 = _GEN_1294 | valid_array_0_57; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_451 = _GEN_1295 | valid_array_0_58; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_452 = _GEN_1296 | valid_array_0_59; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_453 = _GEN_1297 | valid_array_0_60; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_454 = _GEN_1298 | valid_array_0_61; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_455 = _GEN_1299 | valid_array_0_62; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_456 = _GEN_1300 | valid_array_0_63; // @[ICache.scala 184:39 ICache.scala 184:39 ICache.scala 99:44]
  wire  _GEN_522 = next_way ? 1'h0 : 1'h1; // @[ICache.scala 175:21 CacheBase.scala 72:13 CacheBase.scala 81:13]
  wire  _array_rd_index_T = next_state == 3'h5; // @[ICache.scala 281:17]
  wire [5:0] _array_rd_index_T_1 = _array_rd_index_T ? prev_index : stage1_index; // @[Mux.scala 98:16]
  wire [5:0] array_rd_index = go_on ? prev_index : _array_rd_index_T_1; // @[Mux.scala 98:16]
  wire [5:0] _GEN_523 = next_way ? stage1_index : array_rd_index; // @[ICache.scala 175:21 CacheBase.scala 73:14 CacheBase.scala 82:14]
  wire [127:0] data_array_in = maxi4_manager_io_out_data; // @[ICache.scala 143:39 ICache.scala 284:18]
  wire [127:0] _GEN_524 = next_way ? data_array_in : 128'h0; // @[ICache.scala 175:21 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire [127:0] _GEN_525 = next_way ? 128'h0 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 175:21 CacheBase.scala 75:15 CacheBase.scala 84:15]
  wire [127:0] tag_array_in = {{99'd0}, stage1_tag}; // @[ICache.scala 144:39 ICache.scala 285:18]
  wire [127:0] _GEN_527 = next_way ? tag_array_in : 128'h0; // @[ICache.scala 175:21 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire  _GEN_529 = next_way ? _GEN_265 : valid_array_1_0; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_530 = next_way ? _GEN_266 : valid_array_1_1; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_531 = next_way ? _GEN_267 : valid_array_1_2; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_532 = next_way ? _GEN_268 : valid_array_1_3; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_533 = next_way ? _GEN_269 : valid_array_1_4; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_534 = next_way ? _GEN_270 : valid_array_1_5; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_535 = next_way ? _GEN_271 : valid_array_1_6; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_536 = next_way ? _GEN_272 : valid_array_1_7; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_537 = next_way ? _GEN_273 : valid_array_1_8; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_538 = next_way ? _GEN_274 : valid_array_1_9; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_539 = next_way ? _GEN_275 : valid_array_1_10; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_540 = next_way ? _GEN_276 : valid_array_1_11; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_541 = next_way ? _GEN_277 : valid_array_1_12; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_542 = next_way ? _GEN_278 : valid_array_1_13; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_543 = next_way ? _GEN_279 : valid_array_1_14; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_544 = next_way ? _GEN_280 : valid_array_1_15; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_545 = next_way ? _GEN_281 : valid_array_1_16; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_546 = next_way ? _GEN_282 : valid_array_1_17; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_547 = next_way ? _GEN_283 : valid_array_1_18; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_548 = next_way ? _GEN_284 : valid_array_1_19; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_549 = next_way ? _GEN_285 : valid_array_1_20; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_550 = next_way ? _GEN_286 : valid_array_1_21; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_551 = next_way ? _GEN_287 : valid_array_1_22; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_552 = next_way ? _GEN_288 : valid_array_1_23; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_553 = next_way ? _GEN_289 : valid_array_1_24; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_554 = next_way ? _GEN_290 : valid_array_1_25; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_555 = next_way ? _GEN_291 : valid_array_1_26; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_556 = next_way ? _GEN_292 : valid_array_1_27; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_557 = next_way ? _GEN_293 : valid_array_1_28; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_558 = next_way ? _GEN_294 : valid_array_1_29; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_559 = next_way ? _GEN_295 : valid_array_1_30; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_560 = next_way ? _GEN_296 : valid_array_1_31; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_561 = next_way ? _GEN_297 : valid_array_1_32; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_562 = next_way ? _GEN_298 : valid_array_1_33; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_563 = next_way ? _GEN_299 : valid_array_1_34; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_564 = next_way ? _GEN_300 : valid_array_1_35; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_565 = next_way ? _GEN_301 : valid_array_1_36; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_566 = next_way ? _GEN_302 : valid_array_1_37; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_567 = next_way ? _GEN_303 : valid_array_1_38; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_568 = next_way ? _GEN_304 : valid_array_1_39; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_569 = next_way ? _GEN_305 : valid_array_1_40; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_570 = next_way ? _GEN_306 : valid_array_1_41; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_571 = next_way ? _GEN_307 : valid_array_1_42; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_572 = next_way ? _GEN_308 : valid_array_1_43; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_573 = next_way ? _GEN_309 : valid_array_1_44; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_574 = next_way ? _GEN_310 : valid_array_1_45; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_575 = next_way ? _GEN_311 : valid_array_1_46; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_576 = next_way ? _GEN_312 : valid_array_1_47; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_577 = next_way ? _GEN_313 : valid_array_1_48; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_578 = next_way ? _GEN_314 : valid_array_1_49; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_579 = next_way ? _GEN_315 : valid_array_1_50; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_580 = next_way ? _GEN_316 : valid_array_1_51; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_581 = next_way ? _GEN_317 : valid_array_1_52; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_582 = next_way ? _GEN_318 : valid_array_1_53; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_583 = next_way ? _GEN_319 : valid_array_1_54; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_584 = next_way ? _GEN_320 : valid_array_1_55; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_585 = next_way ? _GEN_321 : valid_array_1_56; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_586 = next_way ? _GEN_322 : valid_array_1_57; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_587 = next_way ? _GEN_323 : valid_array_1_58; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_588 = next_way ? _GEN_324 : valid_array_1_59; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_589 = next_way ? _GEN_325 : valid_array_1_60; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_590 = next_way ? _GEN_326 : valid_array_1_61; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_591 = next_way ? _GEN_327 : valid_array_1_62; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire  _GEN_592 = next_way ? _GEN_328 : valid_array_1_63; // @[ICache.scala 175:21 ICache.scala 100:44]
  wire [5:0] _GEN_594 = next_way ? array_rd_index : stage1_index; // @[ICache.scala 175:21 CacheBase.scala 82:14 CacheBase.scala 73:14]
  wire [127:0] _GEN_595 = next_way ? 128'h0 : data_array_in; // @[ICache.scala 175:21 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire [127:0] _GEN_596 = next_way ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[ICache.scala 175:21 CacheBase.scala 84:15 CacheBase.scala 75:15]
  wire [127:0] _GEN_598 = next_way ? 128'h0 : tag_array_in; // @[ICache.scala 175:21 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire  _GEN_600 = next_way ? valid_array_0_0 : _GEN_393; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_601 = next_way ? valid_array_0_1 : _GEN_394; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_602 = next_way ? valid_array_0_2 : _GEN_395; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_603 = next_way ? valid_array_0_3 : _GEN_396; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_604 = next_way ? valid_array_0_4 : _GEN_397; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_605 = next_way ? valid_array_0_5 : _GEN_398; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_606 = next_way ? valid_array_0_6 : _GEN_399; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_607 = next_way ? valid_array_0_7 : _GEN_400; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_608 = next_way ? valid_array_0_8 : _GEN_401; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_609 = next_way ? valid_array_0_9 : _GEN_402; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_610 = next_way ? valid_array_0_10 : _GEN_403; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_611 = next_way ? valid_array_0_11 : _GEN_404; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_612 = next_way ? valid_array_0_12 : _GEN_405; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_613 = next_way ? valid_array_0_13 : _GEN_406; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_614 = next_way ? valid_array_0_14 : _GEN_407; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_615 = next_way ? valid_array_0_15 : _GEN_408; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_616 = next_way ? valid_array_0_16 : _GEN_409; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_617 = next_way ? valid_array_0_17 : _GEN_410; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_618 = next_way ? valid_array_0_18 : _GEN_411; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_619 = next_way ? valid_array_0_19 : _GEN_412; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_620 = next_way ? valid_array_0_20 : _GEN_413; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_621 = next_way ? valid_array_0_21 : _GEN_414; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_622 = next_way ? valid_array_0_22 : _GEN_415; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_623 = next_way ? valid_array_0_23 : _GEN_416; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_624 = next_way ? valid_array_0_24 : _GEN_417; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_625 = next_way ? valid_array_0_25 : _GEN_418; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_626 = next_way ? valid_array_0_26 : _GEN_419; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_627 = next_way ? valid_array_0_27 : _GEN_420; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_628 = next_way ? valid_array_0_28 : _GEN_421; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_629 = next_way ? valid_array_0_29 : _GEN_422; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_630 = next_way ? valid_array_0_30 : _GEN_423; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_631 = next_way ? valid_array_0_31 : _GEN_424; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_632 = next_way ? valid_array_0_32 : _GEN_425; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_633 = next_way ? valid_array_0_33 : _GEN_426; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_634 = next_way ? valid_array_0_34 : _GEN_427; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_635 = next_way ? valid_array_0_35 : _GEN_428; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_636 = next_way ? valid_array_0_36 : _GEN_429; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_637 = next_way ? valid_array_0_37 : _GEN_430; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_638 = next_way ? valid_array_0_38 : _GEN_431; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_639 = next_way ? valid_array_0_39 : _GEN_432; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_640 = next_way ? valid_array_0_40 : _GEN_433; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_641 = next_way ? valid_array_0_41 : _GEN_434; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_642 = next_way ? valid_array_0_42 : _GEN_435; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_643 = next_way ? valid_array_0_43 : _GEN_436; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_644 = next_way ? valid_array_0_44 : _GEN_437; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_645 = next_way ? valid_array_0_45 : _GEN_438; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_646 = next_way ? valid_array_0_46 : _GEN_439; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_647 = next_way ? valid_array_0_47 : _GEN_440; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_648 = next_way ? valid_array_0_48 : _GEN_441; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_649 = next_way ? valid_array_0_49 : _GEN_442; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_650 = next_way ? valid_array_0_50 : _GEN_443; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_651 = next_way ? valid_array_0_51 : _GEN_444; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_652 = next_way ? valid_array_0_52 : _GEN_445; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_653 = next_way ? valid_array_0_53 : _GEN_446; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_654 = next_way ? valid_array_0_54 : _GEN_447; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_655 = next_way ? valid_array_0_55 : _GEN_448; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_656 = next_way ? valid_array_0_56 : _GEN_449; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_657 = next_way ? valid_array_0_57 : _GEN_450; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_658 = next_way ? valid_array_0_58 : _GEN_451; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_659 = next_way ? valid_array_0_59 : _GEN_452; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_660 = next_way ? valid_array_0_60 : _GEN_453; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_661 = next_way ? valid_array_0_61 : _GEN_454; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_662 = next_way ? valid_array_0_62 : _GEN_455; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_663 = next_way ? valid_array_0_63 : _GEN_456; // @[ICache.scala 175:21 ICache.scala 99:44]
  wire  _GEN_729 = _array_write_T ? _GEN_522 : 1'h1; // @[ICache.scala 174:31 CacheBase.scala 81:13]
  wire [5:0] _GEN_730 = _array_write_T ? _GEN_523 : array_rd_index; // @[ICache.scala 174:31 CacheBase.scala 82:14]
  wire [127:0] _GEN_731 = _array_write_T ? _GEN_524 : 128'h0; // @[ICache.scala 174:31 CacheBase.scala 83:15]
  wire [127:0] _GEN_732 = _array_write_T ? _GEN_525 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 174:31 CacheBase.scala 84:15]
  wire [127:0] _GEN_734 = _array_write_T ? _GEN_527 : 128'h0; // @[ICache.scala 174:31 CacheBase.scala 83:15]
  wire  _GEN_800 = _array_write_T ? next_way : 1'h1; // @[ICache.scala 174:31 CacheBase.scala 81:13]
  wire [5:0] _GEN_801 = _array_write_T ? _GEN_594 : array_rd_index; // @[ICache.scala 174:31 CacheBase.scala 82:14]
  wire [127:0] _GEN_802 = _array_write_T ? _GEN_595 : 128'h0; // @[ICache.scala 174:31 CacheBase.scala 83:15]
  wire [127:0] _GEN_803 = _array_write_T ? _GEN_596 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 174:31 CacheBase.scala 84:15]
  wire [127:0] _GEN_805 = _array_write_T ? _GEN_598 : 128'h0; // @[ICache.scala 174:31 CacheBase.scala 83:15]
  wire [3:0] start_byte = stage1_out_bits_addr[3:0]; // @[ICache.scala 269:51]
  wire [6:0] start_bit = {start_byte, 3'h0}; // @[ICache.scala 270:44]
  wire [127:0] read_data_128 = _T ? cache_line_data_out : maxi4_manager_io_out_data; // @[Mux.scala 98:16]
  wire [127:0] _read_data_T_1 = read_data_128 >> start_bit; // @[ICache.scala 274:84]
  wire  _io_next_bits_data_if2id_pc_T_3 = curr_state != 3'h1 & ~io_cache_reset & go_on; // @[ICache.scala 290:73]
  wire [38:0] _io_next_bits_data_if2id_pc_T_4 = curr_state != 3'h1 & ~io_cache_reset & go_on ? stage1_out_bits_addr : 39'h0
    ; // @[ICache.scala 290:35]
  ysyx_040978_IAXIManager maxi4_manager ( // @[ICache.scala 73:29]
    .clock(maxi4_manager_clock),
    .reset(maxi4_manager_reset),
    .io_in_rd_en(maxi4_manager_io_in_rd_en),
    .io_in_dev(maxi4_manager_io_in_dev),
    .io_in_addr(maxi4_manager_io_in_addr),
    .io_maxi_ar_ready(maxi4_manager_io_maxi_ar_ready),
    .io_maxi_ar_valid(maxi4_manager_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(maxi4_manager_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(maxi4_manager_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(maxi4_manager_io_maxi_ar_bits_size),
    .io_maxi_r_valid(maxi4_manager_io_maxi_r_valid),
    .io_maxi_r_bits_data(maxi4_manager_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(maxi4_manager_io_maxi_r_bits_last),
    .io_out_finish(maxi4_manager_io_out_finish),
    .io_out_ready(maxi4_manager_io_out_ready),
    .io_out_data(maxi4_manager_io_out_data)
  );
  assign io_next_valid = _io_next_bits_data_if2id_pc_T_3 & stage1_out_valid; // @[ICache.scala 291:35]
  assign io_next_bits_data_if2id_inst = addr_underflow ? read_data_128[31:0] : _read_data_T_1[31:0]; // @[ICache.scala 274:30]
  assign io_next_bits_data_if2id_pc = {{25'd0}, _io_next_bits_data_if2id_pc_T_4}; // @[ICache.scala 290:35]
  assign io_prev_ready = next_state == 3'h2 & io_next_ready | io_cache_reset; // @[ICache.scala 129:73]
  assign io_maxi_ar_valid = maxi4_manager_io_maxi_ar_valid; // @[ICache.scala 74:25]
  assign io_maxi_ar_bits_addr = maxi4_manager_io_maxi_ar_bits_addr; // @[ICache.scala 74:25]
  assign io_maxi_ar_bits_len = maxi4_manager_io_maxi_ar_bits_len; // @[ICache.scala 74:25]
  assign io_maxi_ar_bits_size = maxi4_manager_io_maxi_ar_bits_size; // @[ICache.scala 74:25]
  assign io_sram0_addr = array_write ? _GEN_801 : array_rd_index; // @[ICache.scala 173:20 CacheBase.scala 82:14]
  assign io_sram0_wen = array_write ? _GEN_800 : 1'h1; // @[ICache.scala 173:20 CacheBase.scala 81:13]
  assign io_sram0_wmask = array_write ? _GEN_803 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 173:20 CacheBase.scala 84:15]
  assign io_sram0_wdata = array_write ? _GEN_802 : 128'h0; // @[ICache.scala 173:20 CacheBase.scala 83:15]
  assign io_sram1_addr = array_write ? _GEN_730 : array_rd_index; // @[ICache.scala 173:20 CacheBase.scala 82:14]
  assign io_sram1_wen = array_write ? _GEN_729 : 1'h1; // @[ICache.scala 173:20 CacheBase.scala 81:13]
  assign io_sram1_wmask = array_write ? _GEN_732 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 173:20 CacheBase.scala 84:15]
  assign io_sram1_wdata = array_write ? _GEN_731 : 128'h0; // @[ICache.scala 173:20 CacheBase.scala 83:15]
  assign io_sram2_addr = array_write ? _GEN_801 : array_rd_index; // @[ICache.scala 173:20 CacheBase.scala 82:14]
  assign io_sram2_wen = array_write ? _GEN_800 : 1'h1; // @[ICache.scala 173:20 CacheBase.scala 81:13]
  assign io_sram2_wmask = array_write ? _GEN_803 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 173:20 CacheBase.scala 84:15]
  assign io_sram2_wdata = array_write ? _GEN_805 : 128'h0; // @[ICache.scala 173:20 CacheBase.scala 83:15]
  assign io_sram3_addr = array_write ? _GEN_730 : array_rd_index; // @[ICache.scala 173:20 CacheBase.scala 82:14]
  assign io_sram3_wen = array_write ? _GEN_729 : 1'h1; // @[ICache.scala 173:20 CacheBase.scala 81:13]
  assign io_sram3_wmask = array_write ? _GEN_732 : 128'hffffffffffffffffffffffffffffffff; // @[ICache.scala 173:20 CacheBase.scala 84:15]
  assign io_sram3_wdata = array_write ? _GEN_734 : 128'h0; // @[ICache.scala 173:20 CacheBase.scala 83:15]
  assign maxi4_manager_clock = clock;
  assign maxi4_manager_reset = reset;
  assign maxi4_manager_io_in_rd_en = io_cache_reset ? 1'h0 : _GEN_71; // @[ICache.scala 149:20 ICache.scala 150:16]
  assign maxi4_manager_io_in_dev = ~stage1_out_bits_addr[31]; // @[ICache.scala 128:60]
  assign maxi4_manager_io_in_addr = _maxi4_manager_io_in_addr_T_2[31:0]; // @[ICache.scala 162:12]
  assign maxi4_manager_io_maxi_ar_ready = io_maxi_ar_ready; // @[ICache.scala 74:25]
  assign maxi4_manager_io_maxi_r_valid = io_maxi_r_valid; // @[ICache.scala 74:25]
  assign maxi4_manager_io_maxi_r_bits_data = io_maxi_r_bits_data; // @[ICache.scala 74:25]
  assign maxi4_manager_io_maxi_r_bits_last = io_maxi_r_bits_last; // @[ICache.scala 74:25]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 68:37]
      curr_state <= 3'h0; // @[ICache.scala 68:37]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (io_next_ready & io_prev_valid) begin // @[ICache.scala 206:36]
        curr_state <= 3'h2; // @[ICache.scala 206:49]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (maxi4_manager_io_out_finish & io_next_ready) begin // @[ICache.scala 209:37]
        curr_state <= 3'h2; // @[ICache.scala 209:50]
      end else begin
        curr_state <= _GEN_1209;
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_1216;
    end else begin
      curr_state <= _GEN_1231;
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_addr <= 39'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_addr <= io_prev_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_63 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_63 <= _GEN_264;
        end else begin
          lru_list_63 <= _GEN_392;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_62 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_62 <= _GEN_263;
        end else begin
          lru_list_62 <= _GEN_391;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_61 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_61 <= _GEN_262;
        end else begin
          lru_list_61 <= _GEN_390;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_60 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_60 <= _GEN_261;
        end else begin
          lru_list_60 <= _GEN_389;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_59 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_59 <= _GEN_260;
        end else begin
          lru_list_59 <= _GEN_388;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_58 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_58 <= _GEN_259;
        end else begin
          lru_list_58 <= _GEN_387;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_57 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_57 <= _GEN_258;
        end else begin
          lru_list_57 <= _GEN_386;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_56 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_56 <= _GEN_257;
        end else begin
          lru_list_56 <= _GEN_385;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_55 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_55 <= _GEN_256;
        end else begin
          lru_list_55 <= _GEN_384;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_54 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_54 <= _GEN_255;
        end else begin
          lru_list_54 <= _GEN_383;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_53 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_53 <= _GEN_254;
        end else begin
          lru_list_53 <= _GEN_382;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_52 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_52 <= _GEN_253;
        end else begin
          lru_list_52 <= _GEN_381;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_51 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_51 <= _GEN_252;
        end else begin
          lru_list_51 <= _GEN_380;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_50 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_50 <= _GEN_251;
        end else begin
          lru_list_50 <= _GEN_379;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_49 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_49 <= _GEN_250;
        end else begin
          lru_list_49 <= _GEN_378;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_48 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_48 <= _GEN_249;
        end else begin
          lru_list_48 <= _GEN_377;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_47 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_47 <= _GEN_248;
        end else begin
          lru_list_47 <= _GEN_376;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_46 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_46 <= _GEN_247;
        end else begin
          lru_list_46 <= _GEN_375;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_45 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_45 <= _GEN_246;
        end else begin
          lru_list_45 <= _GEN_374;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_44 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_44 <= _GEN_245;
        end else begin
          lru_list_44 <= _GEN_373;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_43 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_43 <= _GEN_244;
        end else begin
          lru_list_43 <= _GEN_372;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_42 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_42 <= _GEN_243;
        end else begin
          lru_list_42 <= _GEN_371;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_41 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_41 <= _GEN_242;
        end else begin
          lru_list_41 <= _GEN_370;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_40 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_40 <= _GEN_241;
        end else begin
          lru_list_40 <= _GEN_369;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_39 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_39 <= _GEN_240;
        end else begin
          lru_list_39 <= _GEN_368;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_38 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_38 <= _GEN_239;
        end else begin
          lru_list_38 <= _GEN_367;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_37 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_37 <= _GEN_238;
        end else begin
          lru_list_37 <= _GEN_366;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_36 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_36 <= _GEN_237;
        end else begin
          lru_list_36 <= _GEN_365;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_35 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_35 <= _GEN_236;
        end else begin
          lru_list_35 <= _GEN_364;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_34 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_34 <= _GEN_235;
        end else begin
          lru_list_34 <= _GEN_363;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_33 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_33 <= _GEN_234;
        end else begin
          lru_list_33 <= _GEN_362;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_32 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_32 <= _GEN_233;
        end else begin
          lru_list_32 <= _GEN_361;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_31 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_31 <= _GEN_232;
        end else begin
          lru_list_31 <= _GEN_360;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_30 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_30 <= _GEN_231;
        end else begin
          lru_list_30 <= _GEN_359;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_29 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_29 <= _GEN_230;
        end else begin
          lru_list_29 <= _GEN_358;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_28 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_28 <= _GEN_229;
        end else begin
          lru_list_28 <= _GEN_357;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_27 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_27 <= _GEN_228;
        end else begin
          lru_list_27 <= _GEN_356;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_26 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_26 <= _GEN_227;
        end else begin
          lru_list_26 <= _GEN_355;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_25 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_25 <= _GEN_226;
        end else begin
          lru_list_25 <= _GEN_354;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_24 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_24 <= _GEN_225;
        end else begin
          lru_list_24 <= _GEN_353;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_23 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_23 <= _GEN_224;
        end else begin
          lru_list_23 <= _GEN_352;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_22 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_22 <= _GEN_223;
        end else begin
          lru_list_22 <= _GEN_351;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_21 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_21 <= _GEN_222;
        end else begin
          lru_list_21 <= _GEN_350;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_20 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_20 <= _GEN_221;
        end else begin
          lru_list_20 <= _GEN_349;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_19 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_19 <= _GEN_220;
        end else begin
          lru_list_19 <= _GEN_348;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_18 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_18 <= _GEN_219;
        end else begin
          lru_list_18 <= _GEN_347;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_17 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_17 <= _GEN_218;
        end else begin
          lru_list_17 <= _GEN_346;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_16 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_16 <= _GEN_217;
        end else begin
          lru_list_16 <= _GEN_345;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_15 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_15 <= _GEN_216;
        end else begin
          lru_list_15 <= _GEN_344;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_14 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_14 <= _GEN_215;
        end else begin
          lru_list_14 <= _GEN_343;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_13 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_13 <= _GEN_214;
        end else begin
          lru_list_13 <= _GEN_342;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_12 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_12 <= _GEN_213;
        end else begin
          lru_list_12 <= _GEN_341;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_11 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_11 <= _GEN_212;
        end else begin
          lru_list_11 <= _GEN_340;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_10 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_10 <= _GEN_211;
        end else begin
          lru_list_10 <= _GEN_339;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_9 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_9 <= _GEN_210;
        end else begin
          lru_list_9 <= _GEN_338;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_8 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_8 <= _GEN_209;
        end else begin
          lru_list_8 <= _GEN_337;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_7 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_7 <= _GEN_208;
        end else begin
          lru_list_7 <= _GEN_336;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_6 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_6 <= _GEN_207;
        end else begin
          lru_list_6 <= _GEN_335;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_5 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_5 <= _GEN_206;
        end else begin
          lru_list_5 <= _GEN_334;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_4 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_4 <= _GEN_205;
        end else begin
          lru_list_4 <= _GEN_333;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_3 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_3 <= _GEN_204;
        end else begin
          lru_list_3 <= _GEN_332;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_2 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_2 <= _GEN_203;
        end else begin
          lru_list_2 <= _GEN_331;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_1 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_1 <= _GEN_202;
        end else begin
          lru_list_1 <= _GEN_330;
        end
      end
    end
    if (reset) begin // @[ICache.scala 103:35]
      lru_list_0 <= 1'h0; // @[ICache.scala 103:35]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        if (next_way) begin // @[ICache.scala 175:21]
          lru_list_0 <= _GEN_201;
        end else begin
          lru_list_0 <= _GEN_329;
        end
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_0 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_0 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_0 <= _GEN_600;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_1 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_1 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_1 <= _GEN_601;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_2 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_2 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_2 <= _GEN_602;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_3 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_3 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_3 <= _GEN_603;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_4 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_4 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_4 <= _GEN_604;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_5 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_5 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_5 <= _GEN_605;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_6 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_6 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_6 <= _GEN_606;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_7 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_7 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_7 <= _GEN_607;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_8 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_8 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_8 <= _GEN_608;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_9 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_9 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_9 <= _GEN_609;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_10 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_10 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_10 <= _GEN_610;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_11 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_11 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_11 <= _GEN_611;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_12 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_12 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_12 <= _GEN_612;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_13 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_13 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_13 <= _GEN_613;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_14 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_14 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_14 <= _GEN_614;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_15 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_15 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_15 <= _GEN_615;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_16 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_16 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_16 <= _GEN_616;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_17 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_17 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_17 <= _GEN_617;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_18 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_18 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_18 <= _GEN_618;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_19 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_19 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_19 <= _GEN_619;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_20 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_20 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_20 <= _GEN_620;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_21 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_21 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_21 <= _GEN_621;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_22 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_22 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_22 <= _GEN_622;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_23 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_23 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_23 <= _GEN_623;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_24 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_24 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_24 <= _GEN_624;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_25 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_25 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_25 <= _GEN_625;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_26 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_26 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_26 <= _GEN_626;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_27 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_27 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_27 <= _GEN_627;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_28 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_28 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_28 <= _GEN_628;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_29 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_29 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_29 <= _GEN_629;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_30 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_30 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_30 <= _GEN_630;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_31 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_31 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_31 <= _GEN_631;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_32 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_32 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_32 <= _GEN_632;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_33 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_33 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_33 <= _GEN_633;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_34 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_34 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_34 <= _GEN_634;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_35 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_35 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_35 <= _GEN_635;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_36 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_36 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_36 <= _GEN_636;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_37 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_37 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_37 <= _GEN_637;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_38 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_38 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_38 <= _GEN_638;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_39 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_39 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_39 <= _GEN_639;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_40 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_40 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_40 <= _GEN_640;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_41 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_41 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_41 <= _GEN_641;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_42 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_42 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_42 <= _GEN_642;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_43 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_43 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_43 <= _GEN_643;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_44 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_44 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_44 <= _GEN_644;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_45 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_45 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_45 <= _GEN_645;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_46 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_46 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_46 <= _GEN_646;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_47 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_47 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_47 <= _GEN_647;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_48 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_48 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_48 <= _GEN_648;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_49 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_49 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_49 <= _GEN_649;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_50 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_50 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_50 <= _GEN_650;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_51 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_51 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_51 <= _GEN_651;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_52 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_52 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_52 <= _GEN_652;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_53 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_53 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_53 <= _GEN_653;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_54 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_54 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_54 <= _GEN_654;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_55 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_55 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_55 <= _GEN_655;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_56 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_56 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_56 <= _GEN_656;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_57 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_57 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_57 <= _GEN_657;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_58 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_58 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_58 <= _GEN_658;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_59 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_59 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_59 <= _GEN_659;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_60 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_60 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_60 <= _GEN_660;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_61 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_61 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_61 <= _GEN_661;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_62 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_62 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_62 <= _GEN_662;
      end
    end
    if (reset) begin // @[ICache.scala 99:44]
      valid_array_0_63 <= 1'h0; // @[ICache.scala 99:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_0_63 <= 1'h0; // @[ICache.scala 190:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_0_63 <= _GEN_663;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_0 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_0 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_0 <= _GEN_529;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_1 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_1 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_1 <= _GEN_530;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_2 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_2 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_2 <= _GEN_531;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_3 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_3 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_3 <= _GEN_532;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_4 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_4 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_4 <= _GEN_533;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_5 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_5 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_5 <= _GEN_534;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_6 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_6 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_6 <= _GEN_535;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_7 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_7 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_7 <= _GEN_536;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_8 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_8 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_8 <= _GEN_537;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_9 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_9 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_9 <= _GEN_538;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_10 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_10 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_10 <= _GEN_539;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_11 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_11 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_11 <= _GEN_540;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_12 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_12 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_12 <= _GEN_541;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_13 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_13 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_13 <= _GEN_542;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_14 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_14 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_14 <= _GEN_543;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_15 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_15 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_15 <= _GEN_544;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_16 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_16 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_16 <= _GEN_545;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_17 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_17 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_17 <= _GEN_546;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_18 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_18 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_18 <= _GEN_547;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_19 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_19 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_19 <= _GEN_548;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_20 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_20 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_20 <= _GEN_549;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_21 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_21 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_21 <= _GEN_550;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_22 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_22 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_22 <= _GEN_551;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_23 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_23 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_23 <= _GEN_552;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_24 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_24 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_24 <= _GEN_553;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_25 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_25 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_25 <= _GEN_554;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_26 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_26 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_26 <= _GEN_555;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_27 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_27 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_27 <= _GEN_556;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_28 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_28 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_28 <= _GEN_557;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_29 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_29 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_29 <= _GEN_558;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_30 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_30 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_30 <= _GEN_559;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_31 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_31 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_31 <= _GEN_560;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_32 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_32 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_32 <= _GEN_561;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_33 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_33 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_33 <= _GEN_562;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_34 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_34 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_34 <= _GEN_563;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_35 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_35 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_35 <= _GEN_564;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_36 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_36 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_36 <= _GEN_565;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_37 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_37 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_37 <= _GEN_566;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_38 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_38 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_38 <= _GEN_567;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_39 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_39 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_39 <= _GEN_568;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_40 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_40 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_40 <= _GEN_569;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_41 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_41 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_41 <= _GEN_570;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_42 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_42 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_42 <= _GEN_571;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_43 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_43 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_43 <= _GEN_572;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_44 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_44 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_44 <= _GEN_573;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_45 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_45 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_45 <= _GEN_574;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_46 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_46 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_46 <= _GEN_575;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_47 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_47 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_47 <= _GEN_576;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_48 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_48 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_48 <= _GEN_577;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_49 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_49 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_49 <= _GEN_578;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_50 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_50 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_50 <= _GEN_579;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_51 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_51 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_51 <= _GEN_580;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_52 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_52 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_52 <= _GEN_581;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_53 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_53 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_53 <= _GEN_582;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_54 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_54 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_54 <= _GEN_583;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_55 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_55 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_55 <= _GEN_584;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_56 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_56 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_56 <= _GEN_585;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_57 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_57 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_57 <= _GEN_586;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_58 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_58 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_58 <= _GEN_587;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_59 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_59 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_59 <= _GEN_588;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_60 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_60 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_60 <= _GEN_589;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_61 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_61 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_61 <= _GEN_590;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_62 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_62 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_62 <= _GEN_591;
      end
    end
    if (reset) begin // @[ICache.scala 100:44]
      valid_array_1_63 <= 1'h0; // @[ICache.scala 100:44]
    end else if (fencei) begin // @[ICache.scala 189:26]
      valid_array_1_63 <= 1'h0; // @[ICache.scala 191:19]
    end else if (array_write) begin // @[ICache.scala 173:20]
      if (_array_write_T) begin // @[ICache.scala 174:31]
        valid_array_1_63 <= _GEN_592;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      if (io_cache_reset) begin // @[ICache.scala 111:25]
        stage1_out_valid <= 1'h0;
      end else begin
        stage1_out_valid <= io_prev_valid;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  stage1_out_bits_addr = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  lru_list_63 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_list_62 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_list_61 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_list_60 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_list_59 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_list_58 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_list_57 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_list_56 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_list_55 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_list_54 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_list_53 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_list_52 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_list_51 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_list_50 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_list_49 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_list_48 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_list_47 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_list_46 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_list_45 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_list_44 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_list_43 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_list_42 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_list_41 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_list_40 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_list_39 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_list_38 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_list_37 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_list_36 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_list_35 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_list_34 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_list_33 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_list_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_list_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_list_30 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_list_29 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_list_28 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_list_27 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_list_26 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_list_25 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_list_24 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_list_23 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_list_22 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_list_21 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_list_20 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_list_19 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_list_18 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_list_17 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_list_16 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_list_15 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_list_14 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_list_13 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_list_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_list_11 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_list_10 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_list_9 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_list_8 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_list_7 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_list_6 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_list_5 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_list_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_list_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_list_2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_list_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_list_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_array_0_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_array_0_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_array_0_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_array_0_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_array_0_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_array_0_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_array_0_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_array_0_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_array_0_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_array_0_9 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_array_0_10 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_array_0_11 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_array_0_12 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_array_0_13 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_array_0_14 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_array_0_15 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_array_0_16 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_array_0_17 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_array_0_18 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_array_0_19 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_array_0_20 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_array_0_21 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_array_0_22 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_array_0_23 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_array_0_24 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_array_0_25 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_array_0_26 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_array_0_27 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_array_0_28 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_array_0_29 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_array_0_30 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_array_0_31 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_array_0_32 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_array_0_33 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_array_0_34 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_array_0_35 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_array_0_36 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_array_0_37 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_array_0_38 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_array_0_39 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_array_0_40 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_array_0_41 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_array_0_42 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_array_0_43 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_array_0_44 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_array_0_45 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_array_0_46 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_array_0_47 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_array_0_48 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_array_0_49 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_array_0_50 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_array_0_51 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_array_0_52 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_array_0_53 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_array_0_54 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_array_0_55 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_array_0_56 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_array_0_57 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_array_0_58 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_array_0_59 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_array_0_60 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_array_0_61 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_array_0_62 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_array_0_63 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_array_1_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_array_1_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_array_1_2 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_array_1_3 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_array_1_4 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_array_1_5 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_array_1_6 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_array_1_7 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_array_1_8 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_array_1_9 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_array_1_10 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_array_1_11 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_array_1_12 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_array_1_13 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_array_1_14 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_array_1_15 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_array_1_16 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_array_1_17 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_array_1_18 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_array_1_19 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_array_1_20 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_array_1_21 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_array_1_22 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_array_1_23 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_array_1_24 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_array_1_25 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_array_1_26 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_array_1_27 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_array_1_28 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_array_1_29 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_array_1_30 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_array_1_31 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_array_1_32 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_array_1_33 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_array_1_34 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_array_1_35 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_array_1_36 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_array_1_37 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_array_1_38 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_array_1_39 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_array_1_40 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_array_1_41 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_array_1_42 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_array_1_43 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_array_1_44 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_array_1_45 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_array_1_46 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_array_1_47 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_array_1_48 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_array_1_49 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_array_1_50 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_array_1_51 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_array_1_52 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_array_1_53 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_array_1_54 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_array_1_55 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_array_1_56 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_array_1_57 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_array_1_58 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_array_1_59 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_array_1_60 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_array_1_61 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_array_1_62 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_array_1_63 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  stage1_out_valid = _RAND_194[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_IFU(
  input          clock,
  input          reset,
  input          io_cache_reset,
  output         io_prev_ready,
  input          io_prev_valid,
  input  [63:0]  io_prev_bits_pc2if_pc,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  input          io_next_ready,
  output         io_next_valid,
  output [31:0]  io_next_bits_if2id_inst,
  output [63:0]  io_next_bits_if2id_pc,
  output [5:0]   io_sram0_addr,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  input          fenceiing
);
  wire  icache_clock; // @[IFU.scala 65:30]
  wire  icache_reset; // @[IFU.scala 65:30]
  wire  icache_io_next_ready; // @[IFU.scala 65:30]
  wire  icache_io_next_valid; // @[IFU.scala 65:30]
  wire [31:0] icache_io_next_bits_data_if2id_inst; // @[IFU.scala 65:30]
  wire [63:0] icache_io_next_bits_data_if2id_pc; // @[IFU.scala 65:30]
  wire  icache_io_cache_reset; // @[IFU.scala 65:30]
  wire  icache_io_prev_ready; // @[IFU.scala 65:30]
  wire  icache_io_prev_valid; // @[IFU.scala 65:30]
  wire [38:0] icache_io_prev_bits_addr; // @[IFU.scala 65:30]
  wire  icache_io_maxi_ar_ready; // @[IFU.scala 65:30]
  wire  icache_io_maxi_ar_valid; // @[IFU.scala 65:30]
  wire [31:0] icache_io_maxi_ar_bits_addr; // @[IFU.scala 65:30]
  wire [7:0] icache_io_maxi_ar_bits_len; // @[IFU.scala 65:30]
  wire [2:0] icache_io_maxi_ar_bits_size; // @[IFU.scala 65:30]
  wire  icache_io_maxi_r_valid; // @[IFU.scala 65:30]
  wire [63:0] icache_io_maxi_r_bits_data; // @[IFU.scala 65:30]
  wire  icache_io_maxi_r_bits_last; // @[IFU.scala 65:30]
  wire [5:0] icache_io_sram0_addr; // @[IFU.scala 65:30]
  wire  icache_io_sram0_wen; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram0_wmask; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram0_wdata; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram0_rdata; // @[IFU.scala 65:30]
  wire [5:0] icache_io_sram1_addr; // @[IFU.scala 65:30]
  wire  icache_io_sram1_wen; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram1_wmask; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram1_wdata; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram1_rdata; // @[IFU.scala 65:30]
  wire [5:0] icache_io_sram2_addr; // @[IFU.scala 65:30]
  wire  icache_io_sram2_wen; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram2_wmask; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram2_wdata; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram2_rdata; // @[IFU.scala 65:30]
  wire [5:0] icache_io_sram3_addr; // @[IFU.scala 65:30]
  wire  icache_io_sram3_wen; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram3_wmask; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram3_wdata; // @[IFU.scala 65:30]
  wire [127:0] icache_io_sram3_rdata; // @[IFU.scala 65:30]
  wire  icache_fencei; // @[IFU.scala 65:30]
  wire  pc_hi = &io_prev_bits_pc2if_pc[63:38]; // @[IFU.scala 59:46]
  wire [37:0] pc2addr_lo = io_prev_bits_pc2if_pc[37:0]; // @[IFU.scala 61:43]
  ysyx_040978_ICacheUnit icache ( // @[IFU.scala 65:30]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_next_ready(icache_io_next_ready),
    .io_next_valid(icache_io_next_valid),
    .io_next_bits_data_if2id_inst(icache_io_next_bits_data_if2id_inst),
    .io_next_bits_data_if2id_pc(icache_io_next_bits_data_if2id_pc),
    .io_cache_reset(icache_io_cache_reset),
    .io_prev_ready(icache_io_prev_ready),
    .io_prev_valid(icache_io_prev_valid),
    .io_prev_bits_addr(icache_io_prev_bits_addr),
    .io_maxi_ar_ready(icache_io_maxi_ar_ready),
    .io_maxi_ar_valid(icache_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(icache_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(icache_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(icache_io_maxi_ar_bits_size),
    .io_maxi_r_valid(icache_io_maxi_r_valid),
    .io_maxi_r_bits_data(icache_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(icache_io_maxi_r_bits_last),
    .io_sram0_addr(icache_io_sram0_addr),
    .io_sram0_wen(icache_io_sram0_wen),
    .io_sram0_wmask(icache_io_sram0_wmask),
    .io_sram0_wdata(icache_io_sram0_wdata),
    .io_sram0_rdata(icache_io_sram0_rdata),
    .io_sram1_addr(icache_io_sram1_addr),
    .io_sram1_wen(icache_io_sram1_wen),
    .io_sram1_wmask(icache_io_sram1_wmask),
    .io_sram1_wdata(icache_io_sram1_wdata),
    .io_sram1_rdata(icache_io_sram1_rdata),
    .io_sram2_addr(icache_io_sram2_addr),
    .io_sram2_wen(icache_io_sram2_wen),
    .io_sram2_wmask(icache_io_sram2_wmask),
    .io_sram2_wdata(icache_io_sram2_wdata),
    .io_sram2_rdata(icache_io_sram2_rdata),
    .io_sram3_addr(icache_io_sram3_addr),
    .io_sram3_wen(icache_io_sram3_wen),
    .io_sram3_wmask(icache_io_sram3_wmask),
    .io_sram3_wdata(icache_io_sram3_wdata),
    .io_sram3_rdata(icache_io_sram3_rdata),
    .fencei(icache_fencei)
  );
  assign io_prev_ready = io_next_ready & icache_io_prev_ready; // @[IFU.scala 83:34]
  assign io_maxi_ar_valid = icache_io_maxi_ar_valid; // @[IFU.scala 74:18]
  assign io_maxi_ar_bits_addr = icache_io_maxi_ar_bits_addr; // @[IFU.scala 74:18]
  assign io_maxi_ar_bits_len = icache_io_maxi_ar_bits_len; // @[IFU.scala 74:18]
  assign io_maxi_ar_bits_size = icache_io_maxi_ar_bits_size; // @[IFU.scala 74:18]
  assign io_next_valid = io_prev_valid & icache_io_next_valid; // @[IFU.scala 84:34]
  assign io_next_bits_if2id_inst = icache_io_next_bits_data_if2id_inst; // @[IFU.scala 70:19]
  assign io_next_bits_if2id_pc = icache_io_next_bits_data_if2id_pc; // @[IFU.scala 70:19]
  assign io_sram0_addr = icache_io_sram0_addr; // @[IFU.scala 78:19]
  assign io_sram0_wen = icache_io_sram0_wen; // @[IFU.scala 78:19]
  assign io_sram0_wmask = icache_io_sram0_wmask; // @[IFU.scala 78:19]
  assign io_sram0_wdata = icache_io_sram0_wdata; // @[IFU.scala 78:19]
  assign io_sram1_addr = icache_io_sram1_addr; // @[IFU.scala 79:19]
  assign io_sram1_wen = icache_io_sram1_wen; // @[IFU.scala 79:19]
  assign io_sram1_wmask = icache_io_sram1_wmask; // @[IFU.scala 79:19]
  assign io_sram1_wdata = icache_io_sram1_wdata; // @[IFU.scala 79:19]
  assign io_sram2_addr = icache_io_sram2_addr; // @[IFU.scala 80:19]
  assign io_sram2_wen = icache_io_sram2_wen; // @[IFU.scala 80:19]
  assign io_sram2_wmask = icache_io_sram2_wmask; // @[IFU.scala 80:19]
  assign io_sram2_wdata = icache_io_sram2_wdata; // @[IFU.scala 80:19]
  assign io_sram3_addr = icache_io_sram3_addr; // @[IFU.scala 81:19]
  assign io_sram3_wen = icache_io_sram3_wen; // @[IFU.scala 81:19]
  assign io_sram3_wmask = icache_io_sram3_wmask; // @[IFU.scala 81:19]
  assign io_sram3_wdata = icache_io_sram3_wdata; // @[IFU.scala 81:19]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_next_ready = io_next_ready; // @[IFU.scala 71:24]
  assign icache_io_cache_reset = io_cache_reset; // @[IFU.scala 73:25]
  assign icache_io_prev_valid = io_prev_valid; // @[IFU.scala 68:24]
  assign icache_io_prev_bits_addr = {pc_hi,pc2addr_lo}; // @[Cat.scala 30:58]
  assign icache_io_maxi_ar_ready = io_maxi_ar_ready; // @[IFU.scala 75:27]
  assign icache_io_maxi_r_valid = io_maxi_r_valid; // @[IFU.scala 74:18]
  assign icache_io_maxi_r_bits_data = io_maxi_r_bits_data; // @[IFU.scala 74:18]
  assign icache_io_maxi_r_bits_last = io_maxi_r_bits_last; // @[IFU.scala 74:18]
  assign icache_io_sram0_rdata = io_sram0_rdata; // @[IFU.scala 78:19]
  assign icache_io_sram1_rdata = io_sram1_rdata; // @[IFU.scala 79:19]
  assign icache_io_sram2_rdata = io_sram2_rdata; // @[IFU.scala 80:19]
  assign icache_io_sram3_rdata = io_sram3_rdata; // @[IFU.scala 81:19]
  assign icache_fencei = fenceiing;
endmodule
module ysyx_040978_IDReg(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_if2id_inst,
  input  [63:0] io_prev_bits_if2id_pc,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_if2id_inst,
  output [63:0] io_next_bits_if2id_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  io_next_valid_r; // @[Reg.scala 27:20]
  reg [31:0] reg_inst; // @[Reg.scala 27:20]
  reg [63:0] reg_pc; // @[Reg.scala 27:20]
  assign io_prev_ready = io_next_ready; // @[IDU.scala 23:11]
  assign io_next_valid = io_next_valid_r; // @[IDU.scala 25:11]
  assign io_next_bits_if2id_inst = reg_inst; // @[IDU.scala 29:12]
  assign io_next_bits_if2id_pc = reg_pc; // @[IDU.scala 29:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      io_next_valid_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      io_next_valid_r <= io_prev_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[IDU.scala 27:17]
        reg_inst <= io_prev_bits_if2id_inst;
      end else begin
        reg_inst <= 32'h13;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[IDU.scala 27:17]
        reg_pc <= io_prev_bits_if2id_pc;
      end else begin
        reg_pc <= 64'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_next_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_inst = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  reg_pc = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_CsrHitCtrl(
  input  [11:0] io_csr_idx,
  output        io_csr_hit_is_mepc,
  output        io_csr_hit_is_mtvec,
  output        io_csr_hit_is_mstatus,
  output        io_csr_hit_is_mie,
  output        io_csr_hit_is_mcause,
  output        io_csr_hit_is_mip,
  output        io_csr_hit_is_mtime,
  output        io_csr_hit_is_mcycle,
  output        io_csr_hit_is_mhartid
);
  assign io_csr_hit_is_mepc = io_csr_idx == 12'h341; // @[Controller.scala 84:41]
  assign io_csr_hit_is_mtvec = io_csr_idx == 12'h305; // @[Controller.scala 85:41]
  assign io_csr_hit_is_mstatus = io_csr_idx == 12'h300; // @[Controller.scala 86:41]
  assign io_csr_hit_is_mie = io_csr_idx == 12'h304; // @[Controller.scala 87:41]
  assign io_csr_hit_is_mcause = io_csr_idx == 12'h342; // @[Controller.scala 88:41]
  assign io_csr_hit_is_mip = io_csr_idx == 12'h344; // @[Controller.scala 89:41]
  assign io_csr_hit_is_mtime = io_csr_idx == 12'h305; // @[Controller.scala 90:41]
  assign io_csr_hit_is_mcycle = io_csr_idx == 12'hb00; // @[Controller.scala 91:41]
  assign io_csr_hit_is_mhartid = io_csr_idx == 12'hf14; // @[Controller.scala 92:41]
endmodule
module ysyx_040978_Controller(
  input  [31:0] io_inst,
  output        io_operator_auipc,
  output        io_operator_lui,
  output        io_operator_jal,
  output        io_operator_jalr,
  output        io_operator_lb,
  output        io_operator_lh,
  output        io_operator_lw,
  output        io_operator_lbu,
  output        io_operator_lhu,
  output        io_operator_ld,
  output        io_operator_lwu,
  output        io_operator_sb,
  output        io_operator_sh,
  output        io_operator_sw,
  output        io_operator_sd,
  output        io_operator_beq,
  output        io_operator_bne,
  output        io_operator_blt,
  output        io_operator_bge,
  output        io_operator_bltu,
  output        io_operator_bgeu,
  output        io_operator_add,
  output        io_operator_sub,
  output        io_operator_sll,
  output        io_operator_slt,
  output        io_operator_sltu,
  output        io_operator_xor,
  output        io_operator_srl,
  output        io_operator_sra,
  output        io_operator_or,
  output        io_operator_and,
  output        io_operator_mul,
  output        io_operator_mulh,
  output        io_operator_mulhu,
  output        io_operator_mulhsu,
  output        io_operator_div,
  output        io_operator_divu,
  output        io_operator_rem,
  output        io_operator_remu,
  output        io_operator_ecall,
  output        io_operator_mret,
  output        io_operator_fencei,
  output        io_operator_csr_is_csr,
  output        io_operator_csr_csrrw,
  output        io_operator_csr_csrrs,
  output        io_operator_csr_csrrc,
  output        io_operator_csr_csrrwi,
  output        io_operator_csr_csrrsi,
  output        io_operator_csr_csrrci,
  output        io_optype_Btype,
  output        io_optype_Jtype,
  output        io_optype_Stype,
  output        io_optype_Rtype,
  output        io_optype_Utype,
  output        io_optype_Itype,
  output        io_srcsize_byte,
  output        io_srcsize_hword,
  output        io_srcsize_word,
  output        io_srcsize_dword,
  output        io_is_load,
  output        io_is_save,
  output        io_csr_hit_is_mepc,
  output        io_csr_hit_is_mtvec,
  output        io_csr_hit_is_mstatus,
  output        io_csr_hit_is_mie,
  output        io_csr_hit_is_mcause,
  output        io_csr_hit_is_mip,
  output        io_csr_hit_is_mtime,
  output        io_csr_hit_is_mcycle,
  output        io_csr_hit_is_mhartid
);
  wire [11:0] csr_hit_ctrl_io_csr_idx; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mepc; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mtvec; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mstatus; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mie; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mcause; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mip; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mtime; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mcycle; // @[Controller.scala 234:36]
  wire  csr_hit_ctrl_io_csr_hit_is_mhartid; // @[Controller.scala 234:36]
  wire [6:0] opcode = io_inst[6:0]; // @[Controller.scala 131:31]
  wire [2:0] fun3 = io_inst[14:12]; // @[Controller.scala 132:29]
  wire [6:0] fun7 = io_inst[31:25]; // @[Controller.scala 133:29]
  wire [5:0] fun6 = io_inst[31:26]; // @[Controller.scala 134:29]
  wire  fun3_000 = fun3 == 3'h0; // @[Controller.scala 141:31]
  wire  fun3_001 = fun3 == 3'h1; // @[Controller.scala 142:31]
  wire  fun3_010 = fun3 == 3'h2; // @[Controller.scala 143:31]
  wire  fun3_011 = fun3 == 3'h3; // @[Controller.scala 144:31]
  wire  fun3_100 = fun3 == 3'h4; // @[Controller.scala 145:31]
  wire  fun3_101 = fun3 == 3'h5; // @[Controller.scala 146:31]
  wire  fun3_110 = fun3 == 3'h6; // @[Controller.scala 147:31]
  wire  fun3_111 = fun3 == 3'h7; // @[Controller.scala 148:31]
  wire  fun7_0000000 = fun7 == 7'h0; // @[Controller.scala 149:35]
  wire  fun7_0000001 = fun7 == 7'h1; // @[Controller.scala 150:35]
  wire  fun7_0100000 = fun7 == 7'h20; // @[Controller.scala 151:35]
  wire  fun6_000000 = fun6 == 6'h0; // @[Controller.scala 152:34]
  wire  fun6_010000 = fun6 == 6'h10; // @[Controller.scala 153:34]
  wire  _io_optype_Rtype_T = opcode == 7'h33; // @[Controller.scala 159:27]
  wire  _io_optype_Rtype_T_1 = opcode == 7'h3b; // @[Controller.scala 159:55]
  wire  _io_optype_Rtype_T_2 = opcode == 7'h33 | opcode == 7'h3b; // @[Controller.scala 159:45]
  wire  _io_optype_Itype_T_1 = opcode == 7'h13; // @[Controller.scala 161:55]
  wire  _io_optype_Itype_T_3 = opcode == 7'h1b; // @[Controller.scala 161:83]
  wire  _io_optype_Itype_T_5 = opcode == 7'h67; // @[Controller.scala 161:111]
  wire  _io_operator_add_T = _io_optype_Rtype_T & fun7_0000000; // @[Controller.scala 193:51]
  wire  _io_operator_add_T_1 = _io_optype_Itype_T_1 | _io_optype_Rtype_T & fun7_0000000; // @[Controller.scala 193:41]
  wire  _io_operator_add_T_3 = _io_optype_Rtype_T_1 & fun7_0000000; // @[Controller.scala 193:87]
  wire  _io_operator_sub_T = _io_optype_Rtype_T & fun7_0100000; // @[Controller.scala 194:42]
  wire  _io_operator_sub_T_1 = _io_optype_Rtype_T_1 & fun7_0100000; // @[Controller.scala 194:68]
  wire  _io_operator_sll_T_6 = _io_optype_Itype_T_1 & fun6_000000 | _io_operator_add_T | _io_optype_Itype_T_3 &
    fun7_0000000 | _io_operator_add_T_3; // @[Controller.scala 195:110]
  wire  fun7_1110011 = opcode == 7'h73; // @[Controller.scala 212:37]
  wire  zero_19_7 = io_inst[19:7] == 13'h0; // @[Controller.scala 221:40]
  ysyx_040978_CsrHitCtrl csr_hit_ctrl ( // @[Controller.scala 234:36]
    .io_csr_idx(csr_hit_ctrl_io_csr_idx),
    .io_csr_hit_is_mepc(csr_hit_ctrl_io_csr_hit_is_mepc),
    .io_csr_hit_is_mtvec(csr_hit_ctrl_io_csr_hit_is_mtvec),
    .io_csr_hit_is_mstatus(csr_hit_ctrl_io_csr_hit_is_mstatus),
    .io_csr_hit_is_mie(csr_hit_ctrl_io_csr_hit_is_mie),
    .io_csr_hit_is_mcause(csr_hit_ctrl_io_csr_hit_is_mcause),
    .io_csr_hit_is_mip(csr_hit_ctrl_io_csr_hit_is_mip),
    .io_csr_hit_is_mtime(csr_hit_ctrl_io_csr_hit_is_mtime),
    .io_csr_hit_is_mcycle(csr_hit_ctrl_io_csr_hit_is_mcycle),
    .io_csr_hit_is_mhartid(csr_hit_ctrl_io_csr_hit_is_mhartid)
  );
  assign io_operator_auipc = opcode == 7'h17; // @[Controller.scala 164:29]
  assign io_operator_lui = opcode == 7'h37; // @[Controller.scala 165:29]
  assign io_operator_jal = opcode == 7'h6f; // @[Controller.scala 166:29]
  assign io_operator_jalr = _io_optype_Itype_T_5 & fun3_000; // @[Controller.scala 167:47]
  assign io_operator_lb = fun3_000 & io_is_load; // @[Controller.scala 170:28]
  assign io_operator_lh = fun3_001 & io_is_load; // @[Controller.scala 171:28]
  assign io_operator_lw = fun3_010 & io_is_load; // @[Controller.scala 172:28]
  assign io_operator_lbu = fun3_100 & io_is_load; // @[Controller.scala 173:28]
  assign io_operator_lhu = fun3_101 & io_is_load; // @[Controller.scala 174:28]
  assign io_operator_ld = fun3_011 & io_is_load; // @[Controller.scala 175:28]
  assign io_operator_lwu = fun3_110 & io_is_load; // @[Controller.scala 176:28]
  assign io_operator_sb = fun3_000 & io_is_save; // @[Controller.scala 178:28]
  assign io_operator_sh = fun3_001 & io_is_save; // @[Controller.scala 179:28]
  assign io_operator_sw = fun3_010 & io_is_save; // @[Controller.scala 180:28]
  assign io_operator_sd = fun3_011 & io_is_save; // @[Controller.scala 181:28]
  assign io_operator_beq = fun3_000 & io_optype_Btype; // @[Controller.scala 182:28]
  assign io_operator_bne = fun3_001 & io_optype_Btype; // @[Controller.scala 183:28]
  assign io_operator_blt = fun3_100 & io_optype_Btype; // @[Controller.scala 184:28]
  assign io_operator_bge = fun3_101 & io_optype_Btype; // @[Controller.scala 185:28]
  assign io_operator_bltu = fun3_110 & io_optype_Btype; // @[Controller.scala 186:28]
  assign io_operator_bgeu = fun3_111 & io_optype_Btype; // @[Controller.scala 187:28]
  assign io_operator_add = fun3_000 & (_io_optype_Itype_T_1 | _io_optype_Rtype_T & fun7_0000000 | _io_optype_Itype_T_3
     | _io_optype_Rtype_T_1 & fun7_0000000); // @[Controller.scala 193:31]
  assign io_operator_sub = fun3_000 & (_io_optype_Rtype_T & fun7_0100000 | _io_optype_Rtype_T_1 & fun7_0100000); // @[Controller.scala 194:31]
  assign io_operator_sll = fun3_001 & (_io_optype_Itype_T_1 & fun6_000000 | _io_operator_add_T | _io_optype_Itype_T_3 &
    fun7_0000000 | _io_operator_add_T_3); // @[Controller.scala 195:31]
  assign io_operator_slt = fun3_010 & _io_operator_add_T_1; // @[Controller.scala 196:31]
  assign io_operator_sltu = fun3_011 & _io_operator_add_T_1; // @[Controller.scala 197:31]
  assign io_operator_xor = fun3_100 & _io_operator_add_T_1; // @[Controller.scala 198:31]
  assign io_operator_srl = fun3_101 & _io_operator_sll_T_6; // @[Controller.scala 199:31]
  assign io_operator_sra = fun3_101 & (_io_optype_Itype_T_1 & fun6_010000 | _io_operator_sub_T | _io_optype_Itype_T_3 &
    fun7_0100000 | _io_operator_sub_T_1); // @[Controller.scala 200:31]
  assign io_operator_or = fun3_110 & _io_operator_add_T_1; // @[Controller.scala 201:31]
  assign io_operator_and = fun3_111 & _io_operator_add_T_1; // @[Controller.scala 202:31]
  assign io_operator_mul = fun3_000 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 203:46]
  assign io_operator_mulh = fun3_001 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 204:46]
  assign io_operator_mulhu = fun3_011 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 206:46]
  assign io_operator_mulhsu = fun3_010 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 205:46]
  assign io_operator_div = fun3_100 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 207:46]
  assign io_operator_divu = fun3_101 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 208:46]
  assign io_operator_rem = fun3_110 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 209:46]
  assign io_operator_remu = fun3_111 & fun7_0000001 & _io_optype_Rtype_T_2; // @[Controller.scala 210:46]
  assign io_operator_ecall = io_inst[31:20] == 12'h0 & zero_19_7 & fun7_1110011; // @[Controller.scala 222:63]
  assign io_operator_mret = io_inst[31:20] == 12'h302 & zero_19_7 & fun7_1110011; // @[Controller.scala 225:72]
  assign io_operator_fencei = io_inst == 32'h100f; // @[Controller.scala 227:27]
  assign io_operator_csr_is_csr = fun7_1110011 & (fun3_001 | fun3_010 | fun3_011 | fun3_101 | fun3_110 | fun3_111); // @[Controller.scala 219:39]
  assign io_operator_csr_csrrw = fun3_001 & fun7_1110011; // @[Controller.scala 213:35]
  assign io_operator_csr_csrrs = fun3_010 & fun7_1110011; // @[Controller.scala 214:35]
  assign io_operator_csr_csrrc = fun3_011 & fun7_1110011; // @[Controller.scala 215:35]
  assign io_operator_csr_csrrwi = fun3_101 & fun7_1110011; // @[Controller.scala 216:35]
  assign io_operator_csr_csrrsi = fun3_110 & fun7_1110011; // @[Controller.scala 217:35]
  assign io_operator_csr_csrrci = fun3_111 & fun7_1110011; // @[Controller.scala 218:35]
  assign io_optype_Btype = opcode == 7'h63; // @[Controller.scala 156:27]
  assign io_optype_Jtype = opcode == 7'h6f; // @[Controller.scala 157:27]
  assign io_optype_Stype = opcode == 7'h23; // @[Controller.scala 158:27]
  assign io_optype_Rtype = opcode == 7'h33 | opcode == 7'h3b; // @[Controller.scala 159:45]
  assign io_optype_Utype = opcode == 7'h17 | opcode == 7'h37; // @[Controller.scala 160:45]
  assign io_optype_Itype = opcode == 7'h3 | opcode == 7'h13 | opcode == 7'h1b | opcode == 7'h67; // @[Controller.scala 161:101]
  assign io_srcsize_byte = io_operator_lb | io_operator_lbu | io_operator_sb; // @[Controller.scala 229:47]
  assign io_srcsize_hword = io_operator_lh | io_operator_lhu | io_operator_sh; // @[Controller.scala 230:47]
  assign io_srcsize_word = io_operator_lw | io_operator_lwu | io_operator_sw | _io_optype_Itype_T_3 |
    _io_optype_Rtype_T_1; // @[Controller.scala 231:71]
  assign io_srcsize_dword = ~(io_srcsize_byte | io_srcsize_hword | io_srcsize_word); // @[Controller.scala 232:20]
  assign io_is_load = opcode == 7'h3; // @[Controller.scala 169:22]
  assign io_is_save = opcode == 7'h23; // @[Controller.scala 177:22]
  assign io_csr_hit_is_mepc = csr_hit_ctrl_io_csr_hit_is_mepc; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mtvec = csr_hit_ctrl_io_csr_hit_is_mtvec; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mstatus = csr_hit_ctrl_io_csr_hit_is_mstatus; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mie = csr_hit_ctrl_io_csr_hit_is_mie; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mcause = csr_hit_ctrl_io_csr_hit_is_mcause; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mip = csr_hit_ctrl_io_csr_hit_is_mip; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mtime = csr_hit_ctrl_io_csr_hit_is_mtime; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mcycle = csr_hit_ctrl_io_csr_hit_is_mcycle; // @[Controller.scala 236:14]
  assign io_csr_hit_is_mhartid = csr_hit_ctrl_io_csr_hit_is_mhartid; // @[Controller.scala 236:14]
  assign csr_hit_ctrl_io_csr_idx = io_inst[31:20]; // @[Controller.scala 235:34]
endmodule
module ysyx_040978_MduCtrl(
  input        io_operator_mul,
  input        io_operator_mulh,
  input        io_operator_mulhu,
  input        io_operator_mulhsu,
  input        io_operator_div,
  input        io_operator_divu,
  input        io_operator_rem,
  input        io_operator_remu,
  output       io_mdu_op_mul_signed,
  output       io_mdu_op_is_mu,
  output       io_mdu_op_mul_32,
  output [1:0] io_mdu_op_div_signed,
  output       io_mdu_op_is_div,
  output       io_mdu_op_is_du
);
  wire  _io_mdu_op_is_mu_T = io_operator_mul | io_operator_mulh; // @[Controller.scala 111:36]
  wire  io_mdu_op_mul_signed_hi = _io_mdu_op_is_mu_T | io_operator_mulhsu; // @[Controller.scala 112:60]
  wire [1:0] _io_mdu_op_mul_signed_T_1 = {io_mdu_op_mul_signed_hi,_io_mdu_op_is_mu_T}; // @[Cat.scala 30:58]
  wire  _io_mdu_op_div_signed_T = io_operator_div | io_operator_rem; // @[Controller.scala 116:40]
  assign io_mdu_op_mul_signed = _io_mdu_op_mul_signed_T_1[0]; // @[Controller.scala 112:24]
  assign io_mdu_op_is_mu = io_operator_mul | io_operator_mulh | io_operator_mulhu | io_operator_mulhsu; // @[Controller.scala 111:69]
  assign io_mdu_op_mul_32 = io_operator_mul; // @[Controller.scala 113:20]
  assign io_mdu_op_div_signed = {{1'd0}, _io_mdu_op_div_signed_T}; // @[Controller.scala 116:40]
  assign io_mdu_op_is_div = io_operator_div | io_operator_divu; // @[Controller.scala 115:36]
  assign io_mdu_op_is_du = io_operator_div | io_operator_divu | io_operator_rem | io_operator_remu; // @[Controller.scala 114:67]
endmodule
module ysyx_040978_IDU(
  input         clock,
  input         reset,
  output [4:0]  io_regfile_addr1,
  input  [63:0] io_regfile_data1,
  output [4:0]  io_regfile_addr2,
  input  [63:0] io_regfile_data2,
  input  [63:0] io_fwu_fw_src1_data,
  input  [63:0] io_fwu_fw_src2_data,
  output        io_fwu_optype_Itype,
  output [4:0]  io_fwu_src1_addr,
  output [4:0]  io_fwu_src2_addr,
  output [63:0] io_fwu_src1_data,
  output [63:0] io_fwu_src2_data,
  output        io_bru_brh,
  output        io_bru_jal,
  output        io_bru_jalr,
  output [63:0] io_bru_pc,
  output [63:0] io_bru_src1,
  output [63:0] io_bru_src2,
  output [63:0] io_bru_imm,
  input  [63:0] io_csr_out_mepc,
  input  [63:0] io_csr_out_mtvec,
  input         io_csr_out_mie,
  input         io_csr_out_mtie,
  input         io_csr_out_msie,
  input         io_csr_out_meie,
  input         io_csr_out_mtip,
  input         io_csr_out_msip,
  input         io_csr_out_meip,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_if2id_inst,
  input  [63:0] io_prev_bits_if2id_pc,
  input         io_next_ready,
  output        io_next_valid,
  output [63:0] io_next_bits_id2ex_alu_src1,
  output [63:0] io_next_bits_id2ex_alu_src2,
  output [63:0] io_next_bits_id2ex_salu_src1,
  output [63:0] io_next_bits_id2ex_salu_src2,
  output [63:0] io_next_bits_id2ex_src1,
  output [63:0] io_next_bits_id2ex_src2,
  output [63:0] io_next_bits_id2ex_src3,
  output        io_next_bits_id2ex_operator_auipc,
  output        io_next_bits_id2ex_operator_lui,
  output        io_next_bits_id2ex_operator_jal,
  output        io_next_bits_id2ex_operator_jalr,
  output        io_next_bits_id2ex_operator_sb,
  output        io_next_bits_id2ex_operator_sh,
  output        io_next_bits_id2ex_operator_sw,
  output        io_next_bits_id2ex_operator_sd,
  output        io_next_bits_id2ex_operator_add,
  output        io_next_bits_id2ex_operator_sub,
  output        io_next_bits_id2ex_operator_sll,
  output        io_next_bits_id2ex_operator_slt,
  output        io_next_bits_id2ex_operator_sltu,
  output        io_next_bits_id2ex_operator_xor,
  output        io_next_bits_id2ex_operator_srl,
  output        io_next_bits_id2ex_operator_sra,
  output        io_next_bits_id2ex_operator_or,
  output        io_next_bits_id2ex_operator_and,
  output        io_next_bits_id2ex_operator_csr_is_csr,
  output        io_next_bits_id2ex_operator_csr_csrrw,
  output        io_next_bits_id2ex_operator_csr_csrrs,
  output        io_next_bits_id2ex_operator_csr_csrrc,
  output        io_next_bits_id2ex_operator_csr_csrrwi,
  output        io_next_bits_id2ex_operator_csr_csrrsi,
  output        io_next_bits_id2ex_operator_csr_csrrci,
  output        io_next_bits_id2ex_srcsize_byte,
  output        io_next_bits_id2ex_srcsize_hword,
  output        io_next_bits_id2ex_srcsize_word,
  output        io_next_bits_id2ex_srcsize_dword,
  output        io_next_bits_id2ex_is_load,
  output        io_next_bits_id2ex_is_save,
  output        io_next_bits_id2ex_div_inf,
  output        io_next_bits_id2ex_csr_we,
  output        io_next_bits_id2ex_csr_hit_is_mepc,
  output        io_next_bits_id2ex_csr_hit_is_mtvec,
  output        io_next_bits_id2ex_csr_hit_is_mstatus,
  output        io_next_bits_id2ex_csr_hit_is_mie,
  output        io_next_bits_id2ex_csr_hit_is_mcause,
  output        io_next_bits_id2ex_csr_hit_is_mip,
  output        io_next_bits_id2ex_csr_hit_is_mtime,
  output        io_next_bits_id2ex_csr_hit_is_mcycle,
  output        io_next_bits_id2ex_csr_hit_is_mhartid,
  output        io_next_bits_id2ex_mdu_op_mul_signed,
  output        io_next_bits_id2ex_mdu_op_is_mu,
  output        io_next_bits_id2ex_mdu_op_mul_32,
  output [1:0]  io_next_bits_id2ex_mdu_op_div_signed,
  output        io_next_bits_id2ex_mdu_op_is_div,
  output        io_next_bits_id2ex_mdu_op_is_du,
  output [4:0]  io_next_bits_id2ex_zimm,
  output        io_next_bits_id2ex_intr,
  output        io_next_bits_id2ex_exec,
  output        io_next_bits_id2ex_mret,
  output [3:0]  io_next_bits_id2ex_exce_code,
  output [63:0] io_next_bits_id2ex_pc,
  output        io_next_bits_id2ex_is_iem,
  output        io_next_bits_id2mem_fencei,
  output        io_next_bits_id2mem_size_byte,
  output        io_next_bits_id2mem_size_hword,
  output        io_next_bits_id2mem_size_word,
  output        io_next_bits_id2mem_size_dword,
  output        io_next_bits_id2mem_sext_flag,
  output        io_next_bits_id2mem_memory_rd_en,
  output        io_next_bits_id2mem_memory_we_en,
  output        io_next_bits_id2wb_intr_exce_ret,
  output        io_next_bits_id2wb_fencei,
  output        io_next_bits_id2wb_wb_sel,
  output        io_next_bits_id2wb_regfile_we_en,
  output [4:0]  io_next_bits_id2wb_regfile_we_addr,
  input         wb_fencei_0,
  input         wb_intr_exce_ret_0,
  output        fenceiing_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] ctrl_io_inst; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_auipc; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lui; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_jal; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_jalr; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lb; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lh; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lw; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lbu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lhu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_ld; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_lwu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sb; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sh; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sw; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sd; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_beq; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_bne; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_blt; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_bge; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_bltu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_bgeu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_add; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sub; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sll; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_slt; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sltu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_xor; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_srl; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_sra; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_or; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_and; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_mul; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_mulh; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_mulhu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_mulhsu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_div; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_divu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_rem; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_remu; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_ecall; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_mret; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_fencei; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_is_csr; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrw; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrs; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrc; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrwi; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrsi; // @[IDU.scala 53:20]
  wire  ctrl_io_operator_csr_csrrci; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Btype; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Jtype; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Stype; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Rtype; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Utype; // @[IDU.scala 53:20]
  wire  ctrl_io_optype_Itype; // @[IDU.scala 53:20]
  wire  ctrl_io_srcsize_byte; // @[IDU.scala 53:20]
  wire  ctrl_io_srcsize_hword; // @[IDU.scala 53:20]
  wire  ctrl_io_srcsize_word; // @[IDU.scala 53:20]
  wire  ctrl_io_srcsize_dword; // @[IDU.scala 53:20]
  wire  ctrl_io_is_load; // @[IDU.scala 53:20]
  wire  ctrl_io_is_save; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mepc; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mtvec; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mstatus; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mie; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mcause; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mip; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mtime; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mcycle; // @[IDU.scala 53:20]
  wire  ctrl_io_csr_hit_is_mhartid; // @[IDU.scala 53:20]
  wire  mdu_ctrl_io_operator_mul; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_mulh; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_mulhu; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_mulhsu; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_div; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_divu; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_rem; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_operator_remu; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_mdu_op_mul_signed; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_mdu_op_is_mu; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_mdu_op_mul_32; // @[IDU.scala 143:32]
  wire [1:0] mdu_ctrl_io_mdu_op_div_signed; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_mdu_op_is_div; // @[IDU.scala 143:32]
  wire  mdu_ctrl_io_mdu_op_is_du; // @[IDU.scala 143:32]
  wire  _io_next_bits_id2ex_csr_we_T = ctrl_io_operator_csr_csrrw | ctrl_io_operator_csr_csrrwi; // @[IDU.scala 108:26]
  wire  _io_next_bits_id2ex_csr_we_T_1 = ctrl_io_operator_csr_csrrs | ctrl_io_operator_csr_csrrc; // @[IDU.scala 109:26]
  wire  _io_next_bits_id2ex_csr_we_T_2 = io_next_bits_id2ex_zimm != 5'h0; // @[IDU.scala 109:62]
  wire  _io_next_bits_id2ex_csr_we_T_3 = ctrl_io_operator_csr_csrrsi | ctrl_io_operator_csr_csrrci; // @[IDU.scala 110:26]
  wire  _io_next_bits_id2ex_csr_we_T_6 = _io_next_bits_id2ex_csr_we_T_1 ? _io_next_bits_id2ex_csr_we_T_2 :
    _io_next_bits_id2ex_csr_we_T_3 & _io_next_bits_id2ex_csr_we_T_2; // @[Mux.scala 98:16]
  wire [19:0] exb_src1_Utype_hi = io_prev_bits_if2id_inst[31:12]; // @[IDU.scala 116:29]
  wire [31:0] _exb_src1_Utype_T_1 = {exb_src1_Utype_hi,12'h0}; // @[IDU.scala 116:54]
  wire  _io_next_bits_id2ex_src1_T = ctrl_io_optype_Rtype | ctrl_io_optype_Itype; // @[IDU.scala 119:22]
  wire  _io_next_bits_id2ex_src1_T_1 = _io_next_bits_id2ex_src1_T | ctrl_io_optype_Btype; // @[IDU.scala 120:22]
  wire  _io_next_bits_id2ex_src1_T_2 = _io_next_bits_id2ex_src1_T_1 | ctrl_io_optype_Stype; // @[IDU.scala 121:22]
  wire  _io_next_bits_id2ex_src1_T_3 = _io_next_bits_id2ex_src1_T_2 | ctrl_io_operator_csr_is_csr; // @[IDU.scala 122:22]
  wire [63:0] _io_next_bits_id2ex_src1_T_4 = {{32{_exb_src1_Utype_T_1[31]}},_exb_src1_Utype_T_1}; // @[IDU.scala 125:38]
  wire [63:0] _io_next_bits_id2ex_src1_T_5 = ctrl_io_optype_Utype ? _io_next_bits_id2ex_src1_T_4 : 64'h0; // @[Mux.scala 98:16]
  wire [11:0] _exb_src2_Itype_T_1 = io_prev_bits_if2id_inst[31:20]; // @[IDU.scala 129:39]
  wire  _io_next_bits_id2ex_src2_T_1 = ctrl_io_optype_Rtype | ctrl_io_optype_Stype | ctrl_io_optype_Btype; // @[IDU.scala 132:36]
  wire [63:0] _io_next_bits_id2ex_src2_T_2 = {{52{_exb_src2_Itype_T_1[11]}},_exb_src2_Itype_T_1}; // @[IDU.scala 133:40]
  wire [63:0] _io_next_bits_id2ex_src2_T_3 = ctrl_io_optype_Itype ? _io_next_bits_id2ex_src2_T_2 : 64'h0; // @[Mux.scala 98:16]
  wire [31:0] _io_next_bits_id2ex_salu_src1_T_1 = io_fwu_fw_src1_data[31:0]; // @[IDU.scala 138:61]
  wire [31:0] _io_next_bits_id2ex_salu_src2_T_1 = io_next_bits_id2ex_src2[31:0]; // @[IDU.scala 139:60]
  wire  _io_next_bits_id2ex_div_inf_T = io_next_bits_id2ex_src2 == 64'h0; // @[IDU.scala 141:27]
  wire  _mdu_ctrl_io_operator_div_T = ~_io_next_bits_id2ex_div_inf_T; // @[IDU.scala 148:39]
  wire [6:0] exb_src3_false_hi = io_prev_bits_if2id_inst[31:25]; // @[IDU.scala 155:29]
  wire [11:0] _exb_src3_false_T_1 = {exb_src3_false_hi,io_prev_bits_if2id_inst[11:7]}; // @[IDU.scala 155:52]
  wire [63:0] _io_next_bits_id2ex_src3_T_2 = {{52{_exb_src3_false_T_1[11]}},_exb_src3_false_T_1}; // @[IDU.scala 156:83]
  wire  beq_jump = ctrl_io_operator_beq & io_fwu_fw_src1_data == io_fwu_fw_src2_data; // @[IDU.scala 158:31]
  wire  bne_jump = ctrl_io_operator_bne & io_fwu_fw_src1_data != io_fwu_fw_src2_data; // @[IDU.scala 159:31]
  wire  blt_jump = ctrl_io_operator_blt & $signed(io_fwu_fw_src1_data) < $signed(io_fwu_fw_src2_data); // @[IDU.scala 160:31]
  wire  bge_jump = ctrl_io_operator_bge & $signed(io_fwu_fw_src1_data) >= $signed(io_fwu_fw_src2_data); // @[IDU.scala 161:31]
  wire  bltu_jump = ctrl_io_operator_bltu & io_fwu_fw_src1_data < io_fwu_fw_src2_data; // @[IDU.scala 162:33]
  wire  bgeu_jump = ctrl_io_operator_bgeu & io_fwu_fw_src1_data >= io_fwu_fw_src2_data; // @[IDU.scala 163:33]
  wire  branch = beq_jump | bne_jump | blt_jump | bge_jump | bltu_jump | bgeu_jump; // @[IDU.scala 164:70]
  wire  brb_imm_jal_hi_hi_hi = io_prev_bits_if2id_inst[31]; // @[IDU.scala 172:26]
  wire [7:0] brb_imm_jal_hi_hi_lo = io_prev_bits_if2id_inst[19:12]; // @[IDU.scala 172:36]
  wire  brb_imm_jal_hi_lo = io_prev_bits_if2id_inst[20]; // @[IDU.scala 172:50]
  wire [5:0] brb_imm_jal_lo_hi_hi = io_prev_bits_if2id_inst[30:25]; // @[IDU.scala 172:60]
  wire [3:0] brb_imm_jal_lo_hi_lo = io_prev_bits_if2id_inst[24:21]; // @[IDU.scala 172:74]
  wire [20:0] _brb_imm_jal_T_1 = {brb_imm_jal_hi_hi_hi,brb_imm_jal_hi_hi_lo,brb_imm_jal_hi_lo,brb_imm_jal_lo_hi_hi,
    brb_imm_jal_lo_hi_lo,1'h0}; // @[IDU.scala 172:94]
  wire  brb_imm_branch_hi_hi_lo = io_prev_bits_if2id_inst[7]; // @[IDU.scala 174:39]
  wire [3:0] brb_imm_branch_lo_hi = io_prev_bits_if2id_inst[11:8]; // @[IDU.scala 174:62]
  wire [12:0] _brb_imm_branch_T_1 = {brb_imm_jal_hi_hi_hi,brb_imm_branch_hi_hi_lo,brb_imm_jal_lo_hi_hi,
    brb_imm_branch_lo_hi,1'h0}; // @[IDU.scala 174:76]
  wire [63:0] _io_bru_imm_T = {{43{_brb_imm_jal_T_1[20]}},_brb_imm_jal_T_1}; // @[IDU.scala 177:35]
  wire [63:0] _io_bru_imm_T_1 = {{51{_brb_imm_branch_T_1[12]}},_brb_imm_branch_T_1}; // @[IDU.scala 178:32]
  wire [63:0] _io_bru_imm_T_2 = branch ? _io_bru_imm_T_1 : 64'h0; // @[Mux.scala 98:16]
  reg  fenceiing; // @[IDU.scala 184:26]
  wire  _GEN_0 = ctrl_io_operator_fencei & io_next_ready | fenceiing; // @[IDU.scala 189:46 IDU.scala 190:15 IDU.scala 184:26]
  reg  exce_flushing; // @[IDU.scala 197:38]
  wire  _T_10 = io_csr_out_mie & io_csr_out_meie & io_csr_out_meip; // @[IDU.scala 222:45]
  wire [3:0] _GEN_3 = io_csr_out_mie & io_csr_out_meie & io_csr_out_meip ? 4'hb : 4'h0; // @[IDU.scala 222:61 IDU.scala 224:25 IDU.scala 203:21]
  wire  _GEN_4 = io_csr_out_mie & io_csr_out_mtie & io_csr_out_mtip | _T_10; // @[IDU.scala 219:61 IDU.scala 220:20]
  wire [3:0] _GEN_5 = io_csr_out_mie & io_csr_out_mtie & io_csr_out_mtip ? 4'h7 : _GEN_3; // @[IDU.scala 219:61 IDU.scala 221:25]
  wire  _GEN_6 = io_csr_out_mie & io_csr_out_msie & io_csr_out_msip | _GEN_4; // @[IDU.scala 216:61 IDU.scala 217:20]
  wire [3:0] _GEN_7 = io_csr_out_mie & io_csr_out_msie & io_csr_out_msip ? 4'h3 : _GEN_5; // @[IDU.scala 216:61 IDU.scala 218:25]
  wire  _GEN_8 = ctrl_io_operator_ecall; // @[IDU.scala 213:39 IDU.scala 214:20 IDU.scala 200:16]
  wire [3:0] _GEN_9 = ctrl_io_operator_ecall ? 4'hb : _GEN_7; // @[IDU.scala 213:39 IDU.scala 215:25]
  wire  _GEN_10 = ctrl_io_operator_ecall ? 1'h0 : _GEN_6; // @[IDU.scala 213:39 IDU.scala 199:16]
  wire  _GEN_11 = ctrl_io_operator_mret; // @[IDU.scala 211:38 IDU.scala 212:20 IDU.scala 202:16]
  wire  _GEN_12 = ctrl_io_operator_mret ? 1'h0 : _GEN_8; // @[IDU.scala 211:38 IDU.scala 200:16]
  wire [3:0] _GEN_13 = ctrl_io_operator_mret ? 4'h0 : _GEN_9; // @[IDU.scala 211:38 IDU.scala 203:21]
  wire  _GEN_14 = ctrl_io_operator_mret ? 1'h0 : _GEN_10; // @[IDU.scala 211:38 IDU.scala 199:16]
  wire  _GEN_15 = ctrl_io_operator_jal | ctrl_io_operator_jalr | branch ? 1'h0 : _GEN_14; // @[IDU.scala 207:70 IDU.scala 208:20]
  wire  _GEN_16 = ctrl_io_operator_jal | ctrl_io_operator_jalr | branch ? 1'h0 : _GEN_12; // @[IDU.scala 207:70 IDU.scala 209:20]
  wire  _GEN_17 = ctrl_io_operator_jal | ctrl_io_operator_jalr | branch ? 1'h0 : _GEN_11; // @[IDU.scala 207:70 IDU.scala 210:20]
  wire [3:0] _GEN_18 = ctrl_io_operator_jal | ctrl_io_operator_jalr | branch ? 4'h0 : _GEN_13; // @[IDU.scala 207:70 IDU.scala 203:21]
  wire [3:0] _GEN_19 = exce_flushing ? 4'h0 : _GEN_18; // @[IDU.scala 205:24 IDU.scala 206:25]
  wire  _GEN_20 = exce_flushing ? 1'h0 : _GEN_15; // @[IDU.scala 205:24 IDU.scala 199:16]
  wire  _GEN_21 = exce_flushing ? 1'h0 : _GEN_16; // @[IDU.scala 205:24 IDU.scala 200:16]
  wire  _GEN_22 = exce_flushing ? 1'h0 : _GEN_17; // @[IDU.scala 205:24 IDU.scala 202:16]
  wire  intr_exce_ret = ctrl_io_operator_mret | io_next_bits_id2ex_exec | io_next_bits_id2ex_intr; // @[IDU.scala 229:68]
  wire [63:0] _GEN_27 = ctrl_io_operator_mret ? io_csr_out_mepc : io_next_bits_id2ex_src1; // @[IDU.scala 237:36 IDU.scala 238:15 IDU.scala 169:12]
  wire [63:0] _GEN_28 = ctrl_io_operator_mret ? 64'h0 : io_next_bits_id2ex_src2; // @[IDU.scala 237:36 IDU.scala 239:15 IDU.scala 170:12]
  wire  _GEN_29 = ctrl_io_operator_mret | ctrl_io_operator_jalr & io_next_ready; // @[IDU.scala 237:36 IDU.scala 240:15 IDU.scala 167:12]
  wire  _GEN_30 = ctrl_io_operator_mret ? 1'h0 : ctrl_io_operator_jal & io_next_ready; // @[IDU.scala 237:36 IDU.scala 241:15 IDU.scala 166:12]
  wire  _GEN_31 = ctrl_io_operator_mret ? 1'h0 : branch & io_next_ready; // @[IDU.scala 237:36 IDU.scala 242:15 IDU.scala 165:12]
  wire  _GEN_37 = intr_exce_ret & io_next_ready | exce_flushing; // @[IDU.scala 252:43 IDU.scala 252:59 IDU.scala 197:38]
  wire  _GEN_39 = wb_intr_exce_ret_0 | io_next_ready; // @[IDU.scala 263:31 IDU.scala 264:19 IDU.scala 267:19]
  wire  _GEN_40 = wb_intr_exce_ret_0 ? 1'h0 : io_prev_valid; // @[IDU.scala 263:31 IDU.scala 265:19 IDU.scala 268:19]
  wire  _GEN_41 = intr_exce_ret ? io_next_ready : _GEN_39; // @[IDU.scala 260:28 IDU.scala 261:19]
  wire  _GEN_42 = intr_exce_ret | _GEN_40; // @[IDU.scala 260:28 IDU.scala 262:19]
  wire  _GEN_43 = exce_flushing ? 1'h0 : _GEN_41; // @[IDU.scala 257:28 IDU.scala 258:19]
  wire  _GEN_44 = exce_flushing ? 1'h0 : _GEN_42; // @[IDU.scala 257:28 IDU.scala 259:19]
  ysyx_040978_Controller ctrl ( // @[IDU.scala 53:20]
    .io_inst(ctrl_io_inst),
    .io_operator_auipc(ctrl_io_operator_auipc),
    .io_operator_lui(ctrl_io_operator_lui),
    .io_operator_jal(ctrl_io_operator_jal),
    .io_operator_jalr(ctrl_io_operator_jalr),
    .io_operator_lb(ctrl_io_operator_lb),
    .io_operator_lh(ctrl_io_operator_lh),
    .io_operator_lw(ctrl_io_operator_lw),
    .io_operator_lbu(ctrl_io_operator_lbu),
    .io_operator_lhu(ctrl_io_operator_lhu),
    .io_operator_ld(ctrl_io_operator_ld),
    .io_operator_lwu(ctrl_io_operator_lwu),
    .io_operator_sb(ctrl_io_operator_sb),
    .io_operator_sh(ctrl_io_operator_sh),
    .io_operator_sw(ctrl_io_operator_sw),
    .io_operator_sd(ctrl_io_operator_sd),
    .io_operator_beq(ctrl_io_operator_beq),
    .io_operator_bne(ctrl_io_operator_bne),
    .io_operator_blt(ctrl_io_operator_blt),
    .io_operator_bge(ctrl_io_operator_bge),
    .io_operator_bltu(ctrl_io_operator_bltu),
    .io_operator_bgeu(ctrl_io_operator_bgeu),
    .io_operator_add(ctrl_io_operator_add),
    .io_operator_sub(ctrl_io_operator_sub),
    .io_operator_sll(ctrl_io_operator_sll),
    .io_operator_slt(ctrl_io_operator_slt),
    .io_operator_sltu(ctrl_io_operator_sltu),
    .io_operator_xor(ctrl_io_operator_xor),
    .io_operator_srl(ctrl_io_operator_srl),
    .io_operator_sra(ctrl_io_operator_sra),
    .io_operator_or(ctrl_io_operator_or),
    .io_operator_and(ctrl_io_operator_and),
    .io_operator_mul(ctrl_io_operator_mul),
    .io_operator_mulh(ctrl_io_operator_mulh),
    .io_operator_mulhu(ctrl_io_operator_mulhu),
    .io_operator_mulhsu(ctrl_io_operator_mulhsu),
    .io_operator_div(ctrl_io_operator_div),
    .io_operator_divu(ctrl_io_operator_divu),
    .io_operator_rem(ctrl_io_operator_rem),
    .io_operator_remu(ctrl_io_operator_remu),
    .io_operator_ecall(ctrl_io_operator_ecall),
    .io_operator_mret(ctrl_io_operator_mret),
    .io_operator_fencei(ctrl_io_operator_fencei),
    .io_operator_csr_is_csr(ctrl_io_operator_csr_is_csr),
    .io_operator_csr_csrrw(ctrl_io_operator_csr_csrrw),
    .io_operator_csr_csrrs(ctrl_io_operator_csr_csrrs),
    .io_operator_csr_csrrc(ctrl_io_operator_csr_csrrc),
    .io_operator_csr_csrrwi(ctrl_io_operator_csr_csrrwi),
    .io_operator_csr_csrrsi(ctrl_io_operator_csr_csrrsi),
    .io_operator_csr_csrrci(ctrl_io_operator_csr_csrrci),
    .io_optype_Btype(ctrl_io_optype_Btype),
    .io_optype_Jtype(ctrl_io_optype_Jtype),
    .io_optype_Stype(ctrl_io_optype_Stype),
    .io_optype_Rtype(ctrl_io_optype_Rtype),
    .io_optype_Utype(ctrl_io_optype_Utype),
    .io_optype_Itype(ctrl_io_optype_Itype),
    .io_srcsize_byte(ctrl_io_srcsize_byte),
    .io_srcsize_hword(ctrl_io_srcsize_hword),
    .io_srcsize_word(ctrl_io_srcsize_word),
    .io_srcsize_dword(ctrl_io_srcsize_dword),
    .io_is_load(ctrl_io_is_load),
    .io_is_save(ctrl_io_is_save),
    .io_csr_hit_is_mepc(ctrl_io_csr_hit_is_mepc),
    .io_csr_hit_is_mtvec(ctrl_io_csr_hit_is_mtvec),
    .io_csr_hit_is_mstatus(ctrl_io_csr_hit_is_mstatus),
    .io_csr_hit_is_mie(ctrl_io_csr_hit_is_mie),
    .io_csr_hit_is_mcause(ctrl_io_csr_hit_is_mcause),
    .io_csr_hit_is_mip(ctrl_io_csr_hit_is_mip),
    .io_csr_hit_is_mtime(ctrl_io_csr_hit_is_mtime),
    .io_csr_hit_is_mcycle(ctrl_io_csr_hit_is_mcycle),
    .io_csr_hit_is_mhartid(ctrl_io_csr_hit_is_mhartid)
  );
  ysyx_040978_MduCtrl mdu_ctrl ( // @[IDU.scala 143:32]
    .io_operator_mul(mdu_ctrl_io_operator_mul),
    .io_operator_mulh(mdu_ctrl_io_operator_mulh),
    .io_operator_mulhu(mdu_ctrl_io_operator_mulhu),
    .io_operator_mulhsu(mdu_ctrl_io_operator_mulhsu),
    .io_operator_div(mdu_ctrl_io_operator_div),
    .io_operator_divu(mdu_ctrl_io_operator_divu),
    .io_operator_rem(mdu_ctrl_io_operator_rem),
    .io_operator_remu(mdu_ctrl_io_operator_remu),
    .io_mdu_op_mul_signed(mdu_ctrl_io_mdu_op_mul_signed),
    .io_mdu_op_is_mu(mdu_ctrl_io_mdu_op_is_mu),
    .io_mdu_op_mul_32(mdu_ctrl_io_mdu_op_mul_32),
    .io_mdu_op_div_signed(mdu_ctrl_io_mdu_op_div_signed),
    .io_mdu_op_is_div(mdu_ctrl_io_mdu_op_is_div),
    .io_mdu_op_is_du(mdu_ctrl_io_mdu_op_is_du)
  );
  assign io_regfile_addr1 = io_prev_bits_if2id_inst[19:15]; // @[IDU.scala 64:20]
  assign io_regfile_addr2 = io_prev_bits_if2id_inst[24:20]; // @[IDU.scala 65:20]
  assign io_fwu_optype_Itype = ctrl_io_optype_Itype; // @[IDU.scala 71:14]
  assign io_fwu_src1_addr = io_prev_bits_if2id_inst[19:15]; // @[IDU.scala 75:24]
  assign io_fwu_src2_addr = io_prev_bits_if2id_inst[24:20]; // @[IDU.scala 76:24]
  assign io_fwu_src1_data = io_regfile_data1; // @[IDU.scala 73:17]
  assign io_fwu_src2_data = io_regfile_data2; // @[IDU.scala 74:17]
  assign io_bru_brh = io_next_bits_id2ex_exec | io_next_bits_id2ex_intr ? 1'h0 : _GEN_31; // @[IDU.scala 231:36 IDU.scala 236:15]
  assign io_bru_jal = io_next_bits_id2ex_exec | io_next_bits_id2ex_intr ? 1'h0 : _GEN_30; // @[IDU.scala 231:36 IDU.scala 235:15]
  assign io_bru_jalr = io_next_bits_id2ex_exec | io_next_bits_id2ex_intr | _GEN_29; // @[IDU.scala 231:36 IDU.scala 234:15]
  assign io_bru_pc = io_prev_bits_if2id_pc; // @[IDU.scala 168:12]
  assign io_bru_src1 = io_next_bits_id2ex_exec | io_next_bits_id2ex_intr ? io_csr_out_mtvec : _GEN_27; // @[IDU.scala 231:36 IDU.scala 232:15]
  assign io_bru_src2 = io_next_bits_id2ex_exec | io_next_bits_id2ex_intr ? 64'h0 : _GEN_28; // @[IDU.scala 231:36 IDU.scala 233:15]
  assign io_bru_imm = ctrl_io_operator_jal ? _io_bru_imm_T : _io_bru_imm_T_2; // @[Mux.scala 98:16]
  assign io_prev_ready = ~io_next_ready & ~exce_flushing ? io_next_ready : _GEN_43; // @[IDU.scala 254:40 IDU.scala 255:19]
  assign io_next_valid = ~io_next_ready & ~exce_flushing ? io_prev_valid : _GEN_44; // @[IDU.scala 254:40 IDU.scala 256:19]
  assign io_next_bits_id2ex_alu_src1 = ctrl_io_srcsize_word ? {{32'd0}, io_fwu_fw_src1_data[31:0]} : io_fwu_fw_src1_data
    ; // @[IDU.scala 136:23]
  assign io_next_bits_id2ex_alu_src2 = ctrl_io_srcsize_word ? {{32'd0}, io_next_bits_id2ex_src2[31:0]} :
    io_next_bits_id2ex_src2; // @[IDU.scala 137:23]
  assign io_next_bits_id2ex_salu_src1 = ctrl_io_srcsize_word ? $signed({{32{_io_next_bits_id2ex_salu_src1_T_1[31]}},
    _io_next_bits_id2ex_salu_src1_T_1}) : $signed(io_fwu_fw_src1_data); // @[IDU.scala 138:23]
  assign io_next_bits_id2ex_salu_src2 = ctrl_io_srcsize_word ? $signed({{32{_io_next_bits_id2ex_salu_src2_T_1[31]}},
    _io_next_bits_id2ex_salu_src2_T_1}) : $signed(io_next_bits_id2ex_src2); // @[IDU.scala 139:23]
  assign io_next_bits_id2ex_src1 = _io_next_bits_id2ex_src1_T_3 ? io_fwu_fw_src1_data : _io_next_bits_id2ex_src1_T_5; // @[Mux.scala 98:16]
  assign io_next_bits_id2ex_src2 = _io_next_bits_id2ex_src2_T_1 ? io_fwu_fw_src2_data : _io_next_bits_id2ex_src2_T_3; // @[Mux.scala 98:16]
  assign io_next_bits_id2ex_src3 = ctrl_io_operator_jalr | ctrl_io_optype_Jtype | ctrl_io_optype_Utype ?
    io_prev_bits_if2id_pc : _io_next_bits_id2ex_src3_T_2; // @[IDU.scala 156:18]
  assign io_next_bits_id2ex_operator_auipc = ctrl_io_operator_auipc; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_lui = ctrl_io_operator_lui; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_jal = ctrl_io_operator_jal; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_jalr = ctrl_io_operator_jalr; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sb = ctrl_io_operator_sb; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sh = ctrl_io_operator_sh; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sw = ctrl_io_operator_sw; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sd = ctrl_io_operator_sd; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_add = ctrl_io_operator_add; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sub = ctrl_io_operator_sub; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sll = ctrl_io_operator_sll; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_slt = ctrl_io_operator_slt; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sltu = ctrl_io_operator_sltu; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_xor = ctrl_io_operator_xor; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_srl = ctrl_io_operator_srl; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_sra = ctrl_io_operator_sra; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_or = ctrl_io_operator_or; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_and = ctrl_io_operator_and; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_is_csr = ctrl_io_operator_csr_is_csr; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrw = ctrl_io_operator_csr_csrrw; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrs = ctrl_io_operator_csr_csrrs; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrc = ctrl_io_operator_csr_csrrc; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrwi = ctrl_io_operator_csr_csrrwi; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrsi = ctrl_io_operator_csr_csrrsi; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_operator_csr_csrrci = ctrl_io_operator_csr_csrrci; // @[IDU.scala 102:17]
  assign io_next_bits_id2ex_srcsize_byte = ctrl_io_srcsize_byte; // @[IDU.scala 104:17]
  assign io_next_bits_id2ex_srcsize_hword = ctrl_io_srcsize_hword; // @[IDU.scala 104:17]
  assign io_next_bits_id2ex_srcsize_word = ctrl_io_srcsize_word; // @[IDU.scala 104:17]
  assign io_next_bits_id2ex_srcsize_dword = ctrl_io_srcsize_dword; // @[IDU.scala 104:17]
  assign io_next_bits_id2ex_is_load = ctrl_io_is_load; // @[IDU.scala 105:17]
  assign io_next_bits_id2ex_is_save = ctrl_io_is_save; // @[IDU.scala 106:17]
  assign io_next_bits_id2ex_div_inf = io_next_bits_id2ex_src2 == 64'h0 & (ctrl_io_operator_div | ctrl_io_operator_divu); // @[IDU.scala 141:41]
  assign io_next_bits_id2ex_csr_we = _io_next_bits_id2ex_csr_we_T | _io_next_bits_id2ex_csr_we_T_6; // @[Mux.scala 98:16]
  assign io_next_bits_id2ex_csr_hit_is_mepc = ctrl_io_csr_hit_is_mepc; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mtvec = ctrl_io_csr_hit_is_mtvec; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mstatus = ctrl_io_csr_hit_is_mstatus; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mie = ctrl_io_csr_hit_is_mie; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mcause = ctrl_io_csr_hit_is_mcause; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mip = ctrl_io_csr_hit_is_mip; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mtime = ctrl_io_csr_hit_is_mtime; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mcycle = ctrl_io_csr_hit_is_mcycle; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_csr_hit_is_mhartid = ctrl_io_csr_hit_is_mhartid; // @[IDU.scala 112:17]
  assign io_next_bits_id2ex_mdu_op_mul_signed = mdu_ctrl_io_mdu_op_mul_signed; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_mdu_op_is_mu = mdu_ctrl_io_mdu_op_is_mu; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_mdu_op_mul_32 = mdu_ctrl_io_mdu_op_mul_32; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_mdu_op_div_signed = mdu_ctrl_io_mdu_op_div_signed; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_mdu_op_is_div = mdu_ctrl_io_mdu_op_is_div; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_mdu_op_is_du = mdu_ctrl_io_mdu_op_is_du; // @[IDU.scala 152:14]
  assign io_next_bits_id2ex_zimm = io_prev_bits_if2id_inst[19:15]; // @[IDU.scala 113:24]
  assign io_next_bits_id2ex_intr = io_prev_valid & io_next_ready & _GEN_20; // @[IDU.scala 204:38 IDU.scala 199:16]
  assign io_next_bits_id2ex_exec = io_prev_valid & io_next_ready & _GEN_21; // @[IDU.scala 204:38 IDU.scala 200:16]
  assign io_next_bits_id2ex_mret = io_prev_valid & io_next_ready & _GEN_22; // @[IDU.scala 204:38 IDU.scala 202:16]
  assign io_next_bits_id2ex_exce_code = io_prev_valid & io_next_ready ? _GEN_19 : 4'h0; // @[IDU.scala 204:38 IDU.scala 203:21]
  assign io_next_bits_id2ex_pc = io_prev_bits_if2id_pc; // @[IDU.scala 201:14]
  assign io_next_bits_id2ex_is_iem = ctrl_io_operator_mret | io_next_bits_id2ex_exec | io_next_bits_id2ex_intr; // @[IDU.scala 229:68]
  assign io_next_bits_id2mem_fencei = ctrl_io_operator_fencei; // @[IDU.scala 78:15]
  assign io_next_bits_id2mem_size_byte = ctrl_io_srcsize_byte; // @[IDU.scala 80:13]
  assign io_next_bits_id2mem_size_hword = ctrl_io_srcsize_hword; // @[IDU.scala 80:13]
  assign io_next_bits_id2mem_size_word = ctrl_io_srcsize_word; // @[IDU.scala 80:13]
  assign io_next_bits_id2mem_size_dword = ctrl_io_srcsize_dword; // @[IDU.scala 80:13]
  assign io_next_bits_id2mem_sext_flag = ctrl_io_operator_lb | ctrl_io_operator_lh | ctrl_io_operator_lw |
    ctrl_io_operator_ld & ~(ctrl_io_operator_lbu | ctrl_io_operator_lhu | ctrl_io_operator_lwu); // @[IDU.scala 79:62]
  assign io_next_bits_id2mem_memory_rd_en = ctrl_io_is_load; // @[IDU.scala 82:21]
  assign io_next_bits_id2mem_memory_we_en = ctrl_io_is_save; // @[IDU.scala 81:21]
  assign io_next_bits_id2wb_intr_exce_ret = ctrl_io_operator_mret | io_next_bits_id2ex_exec | io_next_bits_id2ex_intr; // @[IDU.scala 229:68]
  assign io_next_bits_id2wb_fencei = ctrl_io_operator_fencei; // @[IDU.scala 85:14]
  assign io_next_bits_id2wb_wb_sel = ctrl_io_is_load; // @[IDU.scala 86:14]
  assign io_next_bits_id2wb_regfile_we_en = ctrl_io_optype_Utype | ctrl_io_optype_Itype | ctrl_io_optype_Rtype |
    ctrl_io_optype_Jtype | ctrl_io_operator_csr_is_csr; // @[IDU.scala 87:82]
  assign io_next_bits_id2wb_regfile_we_addr = ctrl_io_optype_Btype | ctrl_io_optype_Stype ? 5'h0 :
    io_prev_bits_if2id_inst[11:7]; // @[IDU.scala 88:29]
  assign fenceiing_0 = fenceiing;
  assign ctrl_io_inst = io_prev_bits_if2id_inst; // @[IDU.scala 60:16]
  assign mdu_ctrl_io_operator_mul = ctrl_io_operator_mul; // @[IDU.scala 144:33]
  assign mdu_ctrl_io_operator_mulh = ctrl_io_operator_mulh; // @[IDU.scala 145:33]
  assign mdu_ctrl_io_operator_mulhu = ctrl_io_operator_mulhu; // @[IDU.scala 146:33]
  assign mdu_ctrl_io_operator_mulhsu = ctrl_io_operator_mulhsu; // @[IDU.scala 147:33]
  assign mdu_ctrl_io_operator_div = ~_io_next_bits_id2ex_div_inf_T & ctrl_io_operator_div; // @[IDU.scala 148:50]
  assign mdu_ctrl_io_operator_divu = _mdu_ctrl_io_operator_div_T & ctrl_io_operator_divu; // @[IDU.scala 149:50]
  assign mdu_ctrl_io_operator_rem = ctrl_io_operator_rem; // @[IDU.scala 150:33]
  assign mdu_ctrl_io_operator_remu = ctrl_io_operator_remu; // @[IDU.scala 151:33]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 184:26]
      fenceiing <= 1'h0; // @[IDU.scala 184:26]
    end else if (wb_fencei_0 & io_next_ready) begin // @[IDU.scala 187:36]
      fenceiing <= 1'h0; // @[IDU.scala 188:15]
    end else begin
      fenceiing <= _GEN_0;
    end
    if (reset) begin // @[IDU.scala 197:38]
      exce_flushing <= 1'h0; // @[IDU.scala 197:38]
    end else if (wb_intr_exce_ret_0 & io_next_ready) begin // @[IDU.scala 251:43]
      exce_flushing <= 1'h0; // @[IDU.scala 251:59]
    end else begin
      exce_flushing <= _GEN_37;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fenceiing = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  exce_flushing = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_EXReg(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [63:0] io_prev_bits_id2ex_alu_src1,
  input  [63:0] io_prev_bits_id2ex_alu_src2,
  input  [63:0] io_prev_bits_id2ex_salu_src1,
  input  [63:0] io_prev_bits_id2ex_salu_src2,
  input  [63:0] io_prev_bits_id2ex_src1,
  input  [63:0] io_prev_bits_id2ex_src2,
  input  [63:0] io_prev_bits_id2ex_src3,
  input         io_prev_bits_id2ex_operator_auipc,
  input         io_prev_bits_id2ex_operator_lui,
  input         io_prev_bits_id2ex_operator_jal,
  input         io_prev_bits_id2ex_operator_jalr,
  input         io_prev_bits_id2ex_operator_sb,
  input         io_prev_bits_id2ex_operator_sh,
  input         io_prev_bits_id2ex_operator_sw,
  input         io_prev_bits_id2ex_operator_sd,
  input         io_prev_bits_id2ex_operator_add,
  input         io_prev_bits_id2ex_operator_sub,
  input         io_prev_bits_id2ex_operator_sll,
  input         io_prev_bits_id2ex_operator_slt,
  input         io_prev_bits_id2ex_operator_sltu,
  input         io_prev_bits_id2ex_operator_xor,
  input         io_prev_bits_id2ex_operator_srl,
  input         io_prev_bits_id2ex_operator_sra,
  input         io_prev_bits_id2ex_operator_or,
  input         io_prev_bits_id2ex_operator_and,
  input         io_prev_bits_id2ex_operator_csr_is_csr,
  input         io_prev_bits_id2ex_operator_csr_csrrw,
  input         io_prev_bits_id2ex_operator_csr_csrrs,
  input         io_prev_bits_id2ex_operator_csr_csrrc,
  input         io_prev_bits_id2ex_operator_csr_csrrwi,
  input         io_prev_bits_id2ex_operator_csr_csrrsi,
  input         io_prev_bits_id2ex_operator_csr_csrrci,
  input         io_prev_bits_id2ex_srcsize_byte,
  input         io_prev_bits_id2ex_srcsize_hword,
  input         io_prev_bits_id2ex_srcsize_word,
  input         io_prev_bits_id2ex_srcsize_dword,
  input         io_prev_bits_id2ex_is_load,
  input         io_prev_bits_id2ex_is_save,
  input         io_prev_bits_id2ex_div_inf,
  input         io_prev_bits_id2ex_csr_we,
  input         io_prev_bits_id2ex_csr_hit_is_mepc,
  input         io_prev_bits_id2ex_csr_hit_is_mtvec,
  input         io_prev_bits_id2ex_csr_hit_is_mstatus,
  input         io_prev_bits_id2ex_csr_hit_is_mie,
  input         io_prev_bits_id2ex_csr_hit_is_mcause,
  input         io_prev_bits_id2ex_csr_hit_is_mip,
  input         io_prev_bits_id2ex_csr_hit_is_mtime,
  input         io_prev_bits_id2ex_csr_hit_is_mcycle,
  input         io_prev_bits_id2ex_csr_hit_is_mhartid,
  input         io_prev_bits_id2ex_mdu_op_mul_signed,
  input         io_prev_bits_id2ex_mdu_op_is_mu,
  input         io_prev_bits_id2ex_mdu_op_mul_32,
  input  [1:0]  io_prev_bits_id2ex_mdu_op_div_signed,
  input         io_prev_bits_id2ex_mdu_op_is_div,
  input         io_prev_bits_id2ex_mdu_op_is_du,
  input  [4:0]  io_prev_bits_id2ex_zimm,
  input         io_prev_bits_id2ex_intr,
  input         io_prev_bits_id2ex_exec,
  input         io_prev_bits_id2ex_mret,
  input  [3:0]  io_prev_bits_id2ex_exce_code,
  input  [63:0] io_prev_bits_id2ex_pc,
  input         io_prev_bits_id2ex_is_iem,
  input         io_prev_bits_id2mem_fencei,
  input         io_prev_bits_id2mem_size_byte,
  input         io_prev_bits_id2mem_size_hword,
  input         io_prev_bits_id2mem_size_word,
  input         io_prev_bits_id2mem_size_dword,
  input         io_prev_bits_id2mem_sext_flag,
  input         io_prev_bits_id2mem_memory_rd_en,
  input         io_prev_bits_id2mem_memory_we_en,
  input         io_prev_bits_id2wb_intr_exce_ret,
  input         io_prev_bits_id2wb_fencei,
  input         io_prev_bits_id2wb_wb_sel,
  input         io_prev_bits_id2wb_regfile_we_en,
  input  [4:0]  io_prev_bits_id2wb_regfile_we_addr,
  input         io_next_ready,
  output        io_next_valid,
  output [63:0] io_next_bits_id2ex_alu_src1,
  output [63:0] io_next_bits_id2ex_alu_src2,
  output [63:0] io_next_bits_id2ex_salu_src1,
  output [63:0] io_next_bits_id2ex_salu_src2,
  output [63:0] io_next_bits_id2ex_src1,
  output [63:0] io_next_bits_id2ex_src2,
  output [63:0] io_next_bits_id2ex_src3,
  output        io_next_bits_id2ex_operator_auipc,
  output        io_next_bits_id2ex_operator_lui,
  output        io_next_bits_id2ex_operator_jal,
  output        io_next_bits_id2ex_operator_jalr,
  output        io_next_bits_id2ex_operator_sb,
  output        io_next_bits_id2ex_operator_sh,
  output        io_next_bits_id2ex_operator_sw,
  output        io_next_bits_id2ex_operator_sd,
  output        io_next_bits_id2ex_operator_add,
  output        io_next_bits_id2ex_operator_sub,
  output        io_next_bits_id2ex_operator_sll,
  output        io_next_bits_id2ex_operator_slt,
  output        io_next_bits_id2ex_operator_sltu,
  output        io_next_bits_id2ex_operator_xor,
  output        io_next_bits_id2ex_operator_srl,
  output        io_next_bits_id2ex_operator_sra,
  output        io_next_bits_id2ex_operator_or,
  output        io_next_bits_id2ex_operator_and,
  output        io_next_bits_id2ex_operator_csr_is_csr,
  output        io_next_bits_id2ex_operator_csr_csrrw,
  output        io_next_bits_id2ex_operator_csr_csrrs,
  output        io_next_bits_id2ex_operator_csr_csrrc,
  output        io_next_bits_id2ex_operator_csr_csrrwi,
  output        io_next_bits_id2ex_operator_csr_csrrsi,
  output        io_next_bits_id2ex_operator_csr_csrrci,
  output        io_next_bits_id2ex_srcsize_byte,
  output        io_next_bits_id2ex_srcsize_hword,
  output        io_next_bits_id2ex_srcsize_word,
  output        io_next_bits_id2ex_srcsize_dword,
  output        io_next_bits_id2ex_is_load,
  output        io_next_bits_id2ex_is_save,
  output        io_next_bits_id2ex_div_inf,
  output        io_next_bits_id2ex_csr_we,
  output        io_next_bits_id2ex_csr_hit_is_mepc,
  output        io_next_bits_id2ex_csr_hit_is_mtvec,
  output        io_next_bits_id2ex_csr_hit_is_mstatus,
  output        io_next_bits_id2ex_csr_hit_is_mie,
  output        io_next_bits_id2ex_csr_hit_is_mcause,
  output        io_next_bits_id2ex_csr_hit_is_mip,
  output        io_next_bits_id2ex_csr_hit_is_mtime,
  output        io_next_bits_id2ex_csr_hit_is_mcycle,
  output        io_next_bits_id2ex_csr_hit_is_mhartid,
  output        io_next_bits_id2ex_mdu_op_mul_signed,
  output        io_next_bits_id2ex_mdu_op_is_mu,
  output        io_next_bits_id2ex_mdu_op_mul_32,
  output [1:0]  io_next_bits_id2ex_mdu_op_div_signed,
  output        io_next_bits_id2ex_mdu_op_is_div,
  output        io_next_bits_id2ex_mdu_op_is_du,
  output [4:0]  io_next_bits_id2ex_zimm,
  output        io_next_bits_id2ex_intr,
  output        io_next_bits_id2ex_exec,
  output        io_next_bits_id2ex_mret,
  output [3:0]  io_next_bits_id2ex_exce_code,
  output [63:0] io_next_bits_id2ex_pc,
  output        io_next_bits_id2ex_is_iem,
  output        io_next_bits_id2mem_fencei,
  output        io_next_bits_id2mem_size_byte,
  output        io_next_bits_id2mem_size_hword,
  output        io_next_bits_id2mem_size_word,
  output        io_next_bits_id2mem_size_dword,
  output        io_next_bits_id2mem_sext_flag,
  output        io_next_bits_id2mem_memory_rd_en,
  output        io_next_bits_id2mem_memory_we_en,
  output        io_next_bits_id2wb_intr_exce_ret,
  output        io_next_bits_id2wb_fencei,
  output        io_next_bits_id2wb_wb_sel,
  output        io_next_bits_id2wb_regfile_we_en,
  output [4:0]  io_next_bits_id2wb_regfile_we_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
`endif // RANDOMIZE_REG_INIT
  reg  io_next_valid_r; // @[Reg.scala 27:20]
  wire  data_id2ex_operator_auipc = io_prev_valid & io_prev_bits_id2ex_operator_auipc; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_lui = io_prev_valid & io_prev_bits_id2ex_operator_lui; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_jal = io_prev_valid & io_prev_bits_id2ex_operator_jal; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_jalr = io_prev_valid & io_prev_bits_id2ex_operator_jalr; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sb = io_prev_valid & io_prev_bits_id2ex_operator_sb; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sh = io_prev_valid & io_prev_bits_id2ex_operator_sh; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sw = io_prev_valid & io_prev_bits_id2ex_operator_sw; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sd = io_prev_valid & io_prev_bits_id2ex_operator_sd; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_add = io_prev_valid & io_prev_bits_id2ex_operator_add; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sub = io_prev_valid & io_prev_bits_id2ex_operator_sub; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sll = io_prev_valid & io_prev_bits_id2ex_operator_sll; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_slt = io_prev_valid & io_prev_bits_id2ex_operator_slt; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sltu = io_prev_valid & io_prev_bits_id2ex_operator_sltu; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_xor = io_prev_valid & io_prev_bits_id2ex_operator_xor; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_srl = io_prev_valid & io_prev_bits_id2ex_operator_srl; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_sra = io_prev_valid & io_prev_bits_id2ex_operator_sra; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_or = io_prev_valid & io_prev_bits_id2ex_operator_or; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_and = io_prev_valid & io_prev_bits_id2ex_operator_and; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_is_csr = io_prev_valid & io_prev_bits_id2ex_operator_csr_is_csr; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrw = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrs = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrc = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrwi = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrsi = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 21:17]
  wire  data_id2ex_operator_csr_csrrci = io_prev_valid & io_prev_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 21:17]
  wire  data_id2ex_srcsize_byte = io_prev_valid & io_prev_bits_id2ex_srcsize_byte; // @[EXU.scala 21:17]
  wire  data_id2ex_srcsize_hword = io_prev_valid & io_prev_bits_id2ex_srcsize_hword; // @[EXU.scala 21:17]
  wire  data_id2ex_srcsize_word = io_prev_valid & io_prev_bits_id2ex_srcsize_word; // @[EXU.scala 21:17]
  wire  data_id2ex_srcsize_dword = io_prev_valid & io_prev_bits_id2ex_srcsize_dword; // @[EXU.scala 21:17]
  wire  data_id2ex_is_load = io_prev_valid & io_prev_bits_id2ex_is_load; // @[EXU.scala 21:17]
  wire  data_id2ex_is_save = io_prev_valid & io_prev_bits_id2ex_is_save; // @[EXU.scala 21:17]
  wire  data_id2ex_div_inf = io_prev_valid & io_prev_bits_id2ex_div_inf; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_we = io_prev_valid & io_prev_bits_id2ex_csr_we; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mepc = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mtvec = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mstatus = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mie = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mcause = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mip = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mtime = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mcycle = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 21:17]
  wire  data_id2ex_csr_hit_is_mhartid = io_prev_valid & io_prev_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 21:17]
  wire  data_id2ex_mdu_op_mul_signed = io_prev_valid & io_prev_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 21:17]
  wire  data_id2ex_mdu_op_is_mu = io_prev_valid & io_prev_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 21:17]
  wire  data_id2ex_mdu_op_mul_32 = io_prev_valid & io_prev_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 21:17]
  wire  data_id2ex_mdu_op_is_div = io_prev_valid & io_prev_bits_id2ex_mdu_op_is_div; // @[EXU.scala 21:17]
  wire  data_id2ex_mdu_op_is_du = io_prev_valid & io_prev_bits_id2ex_mdu_op_is_du; // @[EXU.scala 21:17]
  wire  data_id2ex_intr = io_prev_valid & io_prev_bits_id2ex_intr; // @[EXU.scala 21:17]
  wire  data_id2ex_exec = io_prev_valid & io_prev_bits_id2ex_exec; // @[EXU.scala 21:17]
  wire  data_id2ex_mret = io_prev_valid & io_prev_bits_id2ex_mret; // @[EXU.scala 21:17]
  wire  data_id2ex_is_iem = io_prev_valid & io_prev_bits_id2ex_is_iem; // @[EXU.scala 21:17]
  wire  data_id2mem_fencei = io_prev_valid & io_prev_bits_id2mem_fencei; // @[EXU.scala 21:17]
  wire  data_id2mem_size_byte = io_prev_valid & io_prev_bits_id2mem_size_byte; // @[EXU.scala 21:17]
  wire  data_id2mem_size_hword = io_prev_valid & io_prev_bits_id2mem_size_hword; // @[EXU.scala 21:17]
  wire  data_id2mem_size_word = io_prev_valid & io_prev_bits_id2mem_size_word; // @[EXU.scala 21:17]
  wire  data_id2mem_size_dword = io_prev_valid & io_prev_bits_id2mem_size_dword; // @[EXU.scala 21:17]
  wire  data_id2mem_sext_flag = io_prev_valid & io_prev_bits_id2mem_sext_flag; // @[EXU.scala 21:17]
  wire  data_id2mem_memory_rd_en = io_prev_valid & io_prev_bits_id2mem_memory_rd_en; // @[EXU.scala 21:17]
  wire  data_id2mem_memory_we_en = io_prev_valid & io_prev_bits_id2mem_memory_we_en; // @[EXU.scala 21:17]
  wire  data_id2wb_intr_exce_ret = io_prev_valid & io_prev_bits_id2wb_intr_exce_ret; // @[EXU.scala 21:17]
  wire  data_id2wb_fencei = io_prev_valid & io_prev_bits_id2wb_fencei; // @[EXU.scala 21:17]
  wire  data_id2wb_wb_sel = io_prev_valid & io_prev_bits_id2wb_wb_sel; // @[EXU.scala 21:17]
  wire  data_id2wb_regfile_we_en = io_prev_valid & io_prev_bits_id2wb_regfile_we_en; // @[EXU.scala 21:17]
  reg [63:0] reg_id2ex_alu_src1; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_alu_src2; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_salu_src1; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_salu_src2; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_src1; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_src2; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_src3; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_auipc; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_lui; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_jal; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_jalr; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sb; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sh; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sw; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sd; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_add; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sub; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sll; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_slt; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sltu; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_xor; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_srl; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_sra; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_or; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_and; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_is_csr; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrw; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrs; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrc; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrwi; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrsi; // @[Reg.scala 27:20]
  reg  reg_id2ex_operator_csr_csrrci; // @[Reg.scala 27:20]
  reg  reg_id2ex_srcsize_byte; // @[Reg.scala 27:20]
  reg  reg_id2ex_srcsize_hword; // @[Reg.scala 27:20]
  reg  reg_id2ex_srcsize_word; // @[Reg.scala 27:20]
  reg  reg_id2ex_srcsize_dword; // @[Reg.scala 27:20]
  reg  reg_id2ex_is_load; // @[Reg.scala 27:20]
  reg  reg_id2ex_is_save; // @[Reg.scala 27:20]
  reg  reg_id2ex_div_inf; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_we; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mepc; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mtvec; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mstatus; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mie; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mcause; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mip; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mtime; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mcycle; // @[Reg.scala 27:20]
  reg  reg_id2ex_csr_hit_is_mhartid; // @[Reg.scala 27:20]
  reg  reg_id2ex_mdu_op_mul_signed; // @[Reg.scala 27:20]
  reg  reg_id2ex_mdu_op_is_mu; // @[Reg.scala 27:20]
  reg  reg_id2ex_mdu_op_mul_32; // @[Reg.scala 27:20]
  reg [1:0] reg_id2ex_mdu_op_div_signed; // @[Reg.scala 27:20]
  reg  reg_id2ex_mdu_op_is_div; // @[Reg.scala 27:20]
  reg  reg_id2ex_mdu_op_is_du; // @[Reg.scala 27:20]
  reg [4:0] reg_id2ex_zimm; // @[Reg.scala 27:20]
  reg  reg_id2ex_intr; // @[Reg.scala 27:20]
  reg  reg_id2ex_exec; // @[Reg.scala 27:20]
  reg  reg_id2ex_mret; // @[Reg.scala 27:20]
  reg [3:0] reg_id2ex_exce_code; // @[Reg.scala 27:20]
  reg [63:0] reg_id2ex_pc; // @[Reg.scala 27:20]
  reg  reg_id2ex_is_iem; // @[Reg.scala 27:20]
  reg  reg_id2mem_fencei; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_byte; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_hword; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_word; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_dword; // @[Reg.scala 27:20]
  reg  reg_id2mem_sext_flag; // @[Reg.scala 27:20]
  reg  reg_id2mem_memory_rd_en; // @[Reg.scala 27:20]
  reg  reg_id2mem_memory_we_en; // @[Reg.scala 27:20]
  reg  reg_id2wb_intr_exce_ret; // @[Reg.scala 27:20]
  reg  reg_id2wb_fencei; // @[Reg.scala 27:20]
  reg  reg_id2wb_wb_sel; // @[Reg.scala 27:20]
  reg  reg_id2wb_regfile_we_en; // @[Reg.scala 27:20]
  reg [4:0] reg_id2wb_regfile_we_addr; // @[Reg.scala 27:20]
  assign io_prev_ready = io_next_ready; // @[EXU.scala 17:11]
  assign io_next_valid = io_next_valid_r; // @[EXU.scala 19:11]
  assign io_next_bits_id2ex_alu_src1 = reg_id2ex_alu_src1; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_alu_src2 = reg_id2ex_alu_src2; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_salu_src1 = reg_id2ex_salu_src1; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_salu_src2 = reg_id2ex_salu_src2; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_src1 = reg_id2ex_src1; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_src2 = reg_id2ex_src2; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_src3 = reg_id2ex_src3; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_auipc = reg_id2ex_operator_auipc; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_lui = reg_id2ex_operator_lui; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_jal = reg_id2ex_operator_jal; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_jalr = reg_id2ex_operator_jalr; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sb = reg_id2ex_operator_sb; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sh = reg_id2ex_operator_sh; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sw = reg_id2ex_operator_sw; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sd = reg_id2ex_operator_sd; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_add = reg_id2ex_operator_add; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sub = reg_id2ex_operator_sub; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sll = reg_id2ex_operator_sll; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_slt = reg_id2ex_operator_slt; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sltu = reg_id2ex_operator_sltu; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_xor = reg_id2ex_operator_xor; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_srl = reg_id2ex_operator_srl; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_sra = reg_id2ex_operator_sra; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_or = reg_id2ex_operator_or; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_and = reg_id2ex_operator_and; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_is_csr = reg_id2ex_operator_csr_is_csr; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrw = reg_id2ex_operator_csr_csrrw; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrs = reg_id2ex_operator_csr_csrrs; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrc = reg_id2ex_operator_csr_csrrc; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrwi = reg_id2ex_operator_csr_csrrwi; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrsi = reg_id2ex_operator_csr_csrrsi; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_operator_csr_csrrci = reg_id2ex_operator_csr_csrrci; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_srcsize_byte = reg_id2ex_srcsize_byte; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_srcsize_hword = reg_id2ex_srcsize_hword; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_srcsize_word = reg_id2ex_srcsize_word; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_srcsize_dword = reg_id2ex_srcsize_dword; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_is_load = reg_id2ex_is_load; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_is_save = reg_id2ex_is_save; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_div_inf = reg_id2ex_div_inf; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_we = reg_id2ex_csr_we; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mepc = reg_id2ex_csr_hit_is_mepc; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mtvec = reg_id2ex_csr_hit_is_mtvec; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mstatus = reg_id2ex_csr_hit_is_mstatus; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mie = reg_id2ex_csr_hit_is_mie; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mcause = reg_id2ex_csr_hit_is_mcause; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mip = reg_id2ex_csr_hit_is_mip; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mtime = reg_id2ex_csr_hit_is_mtime; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mcycle = reg_id2ex_csr_hit_is_mcycle; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_csr_hit_is_mhartid = reg_id2ex_csr_hit_is_mhartid; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_mul_signed = reg_id2ex_mdu_op_mul_signed; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_is_mu = reg_id2ex_mdu_op_is_mu; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_mul_32 = reg_id2ex_mdu_op_mul_32; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_div_signed = reg_id2ex_mdu_op_div_signed; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_is_div = reg_id2ex_mdu_op_is_div; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mdu_op_is_du = reg_id2ex_mdu_op_is_du; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_zimm = reg_id2ex_zimm; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_intr = reg_id2ex_intr; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_exec = reg_id2ex_exec; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_mret = reg_id2ex_mret; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_exce_code = reg_id2ex_exce_code; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_pc = reg_id2ex_pc; // @[EXU.scala 23:12]
  assign io_next_bits_id2ex_is_iem = reg_id2ex_is_iem; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_fencei = reg_id2mem_fencei; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_size_byte = reg_id2mem_size_byte; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_size_hword = reg_id2mem_size_hword; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_size_word = reg_id2mem_size_word; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_size_dword = reg_id2mem_size_dword; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_sext_flag = reg_id2mem_sext_flag; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_memory_rd_en = reg_id2mem_memory_rd_en; // @[EXU.scala 23:12]
  assign io_next_bits_id2mem_memory_we_en = reg_id2mem_memory_we_en; // @[EXU.scala 23:12]
  assign io_next_bits_id2wb_intr_exce_ret = reg_id2wb_intr_exce_ret; // @[EXU.scala 23:12]
  assign io_next_bits_id2wb_fencei = reg_id2wb_fencei; // @[EXU.scala 23:12]
  assign io_next_bits_id2wb_wb_sel = reg_id2wb_wb_sel; // @[EXU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_en = reg_id2wb_regfile_we_en; // @[EXU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_addr = reg_id2wb_regfile_we_addr; // @[EXU.scala 23:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      io_next_valid_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      io_next_valid_r <= io_prev_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_alu_src1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_alu_src1 <= io_prev_bits_id2ex_alu_src1;
      end else begin
        reg_id2ex_alu_src1 <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_alu_src2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_alu_src2 <= io_prev_bits_id2ex_alu_src2;
      end else begin
        reg_id2ex_alu_src2 <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_salu_src1 <= 64'sh0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_salu_src1 <= io_prev_bits_id2ex_salu_src1;
      end else begin
        reg_id2ex_salu_src1 <= 64'sh0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_salu_src2 <= 64'sh0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_salu_src2 <= io_prev_bits_id2ex_salu_src2;
      end else begin
        reg_id2ex_salu_src2 <= 64'sh0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_src1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_src1 <= io_prev_bits_id2ex_src1;
      end else begin
        reg_id2ex_src1 <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_src2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_src2 <= io_prev_bits_id2ex_src2;
      end else begin
        reg_id2ex_src2 <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_src3 <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_src3 <= io_prev_bits_id2ex_src3;
      end else begin
        reg_id2ex_src3 <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_auipc <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_auipc <= data_id2ex_operator_auipc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_lui <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_lui <= data_id2ex_operator_lui; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_jal <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_jal <= data_id2ex_operator_jal; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_jalr <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_jalr <= data_id2ex_operator_jalr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sb <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sb <= data_id2ex_operator_sb; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sh <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sh <= data_id2ex_operator_sh; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sw <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sw <= data_id2ex_operator_sw; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sd <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sd <= data_id2ex_operator_sd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_add <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_add <= data_id2ex_operator_add; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sub <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sub <= data_id2ex_operator_sub; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sll <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sll <= data_id2ex_operator_sll; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_slt <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_slt <= data_id2ex_operator_slt; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sltu <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sltu <= data_id2ex_operator_sltu; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_xor <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_xor <= data_id2ex_operator_xor; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_srl <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_srl <= data_id2ex_operator_srl; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_sra <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_sra <= data_id2ex_operator_sra; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_or <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_or <= data_id2ex_operator_or; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_and <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_and <= data_id2ex_operator_and; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_is_csr <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_is_csr <= data_id2ex_operator_csr_is_csr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrw <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrw <= data_id2ex_operator_csr_csrrw; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrs <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrs <= data_id2ex_operator_csr_csrrs; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrc <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrc <= data_id2ex_operator_csr_csrrc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrwi <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrwi <= data_id2ex_operator_csr_csrrwi; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrsi <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrsi <= data_id2ex_operator_csr_csrrsi; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_operator_csr_csrrci <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_operator_csr_csrrci <= data_id2ex_operator_csr_csrrci; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_srcsize_byte <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_srcsize_byte <= data_id2ex_srcsize_byte; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_srcsize_hword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_srcsize_hword <= data_id2ex_srcsize_hword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_srcsize_word <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_srcsize_word <= data_id2ex_srcsize_word; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_srcsize_dword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_srcsize_dword <= data_id2ex_srcsize_dword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_is_load <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_is_load <= data_id2ex_is_load; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_is_save <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_is_save <= data_id2ex_is_save; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_div_inf <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_div_inf <= data_id2ex_div_inf; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_we <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_we <= data_id2ex_csr_we; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mepc <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mepc <= data_id2ex_csr_hit_is_mepc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mtvec <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mtvec <= data_id2ex_csr_hit_is_mtvec; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mstatus <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mstatus <= data_id2ex_csr_hit_is_mstatus; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mie <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mie <= data_id2ex_csr_hit_is_mie; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mcause <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mcause <= data_id2ex_csr_hit_is_mcause; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mip <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mip <= data_id2ex_csr_hit_is_mip; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mtime <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mtime <= data_id2ex_csr_hit_is_mtime; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mcycle <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mcycle <= data_id2ex_csr_hit_is_mcycle; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_csr_hit_is_mhartid <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_csr_hit_is_mhartid <= data_id2ex_csr_hit_is_mhartid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_mul_signed <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mdu_op_mul_signed <= data_id2ex_mdu_op_mul_signed; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_is_mu <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mdu_op_is_mu <= data_id2ex_mdu_op_is_mu; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_mul_32 <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mdu_op_mul_32 <= data_id2ex_mdu_op_mul_32; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_div_signed <= 2'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_mdu_op_div_signed <= io_prev_bits_id2ex_mdu_op_div_signed;
      end else begin
        reg_id2ex_mdu_op_div_signed <= 2'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_is_div <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mdu_op_is_div <= data_id2ex_mdu_op_is_div; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mdu_op_is_du <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mdu_op_is_du <= data_id2ex_mdu_op_is_du; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_zimm <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_zimm <= io_prev_bits_id2ex_zimm;
      end else begin
        reg_id2ex_zimm <= 5'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_intr <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_intr <= data_id2ex_intr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_exec <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_exec <= data_id2ex_exec; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_mret <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_mret <= data_id2ex_mret; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_exce_code <= 4'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_exce_code <= io_prev_bits_id2ex_exce_code;
      end else begin
        reg_id2ex_exce_code <= 4'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_pc <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2ex_pc <= io_prev_bits_id2ex_pc;
      end else begin
        reg_id2ex_pc <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2ex_is_iem <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2ex_is_iem <= data_id2ex_is_iem; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_fencei <= data_id2mem_fencei; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_byte <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_byte <= data_id2mem_size_byte; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_hword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_hword <= data_id2mem_size_hword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_word <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_word <= data_id2mem_size_word; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_dword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_dword <= data_id2mem_size_dword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_sext_flag <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_sext_flag <= data_id2mem_sext_flag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_memory_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_memory_rd_en <= data_id2mem_memory_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_memory_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_memory_we_en <= data_id2mem_memory_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_intr_exce_ret <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_intr_exce_ret <= data_id2wb_intr_exce_ret; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_fencei <= data_id2wb_fencei; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_wb_sel <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_wb_sel <= data_id2wb_wb_sel; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_regfile_we_en <= data_id2wb_regfile_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[EXU.scala 21:17]
        reg_id2wb_regfile_we_addr <= io_prev_bits_id2wb_regfile_we_addr;
      end else begin
        reg_id2wb_regfile_we_addr <= 5'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_next_valid_r = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  reg_id2ex_alu_src1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_id2ex_alu_src2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_id2ex_salu_src1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  reg_id2ex_salu_src2 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_id2ex_src1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_id2ex_src2 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_id2ex_src3 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  reg_id2ex_operator_auipc = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  reg_id2ex_operator_lui = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_id2ex_operator_jal = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_id2ex_operator_jalr = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reg_id2ex_operator_sb = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  reg_id2ex_operator_sh = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  reg_id2ex_operator_sw = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_id2ex_operator_sd = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  reg_id2ex_operator_add = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_id2ex_operator_sub = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reg_id2ex_operator_sll = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reg_id2ex_operator_slt = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  reg_id2ex_operator_sltu = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  reg_id2ex_operator_xor = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  reg_id2ex_operator_srl = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  reg_id2ex_operator_sra = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  reg_id2ex_operator_or = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  reg_id2ex_operator_and = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  reg_id2ex_operator_csr_is_csr = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrw = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrs = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrc = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrwi = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrsi = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  reg_id2ex_operator_csr_csrrci = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  reg_id2ex_srcsize_byte = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  reg_id2ex_srcsize_hword = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  reg_id2ex_srcsize_word = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  reg_id2ex_srcsize_dword = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  reg_id2ex_is_load = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  reg_id2ex_is_save = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  reg_id2ex_div_inf = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  reg_id2ex_csr_we = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mepc = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mtvec = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mstatus = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mie = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mcause = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mip = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mtime = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mcycle = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  reg_id2ex_csr_hit_is_mhartid = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  reg_id2ex_mdu_op_mul_signed = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  reg_id2ex_mdu_op_is_mu = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  reg_id2ex_mdu_op_mul_32 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  reg_id2ex_mdu_op_div_signed = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  reg_id2ex_mdu_op_is_div = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  reg_id2ex_mdu_op_is_du = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  reg_id2ex_zimm = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  reg_id2ex_intr = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  reg_id2ex_exec = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  reg_id2ex_mret = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  reg_id2ex_exce_code = _RAND_60[3:0];
  _RAND_61 = {2{`RANDOM}};
  reg_id2ex_pc = _RAND_61[63:0];
  _RAND_62 = {1{`RANDOM}};
  reg_id2ex_is_iem = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  reg_id2mem_fencei = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  reg_id2mem_size_byte = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  reg_id2mem_size_hword = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  reg_id2mem_size_word = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  reg_id2mem_size_dword = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  reg_id2mem_sext_flag = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  reg_id2mem_memory_rd_en = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  reg_id2mem_memory_we_en = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  reg_id2wb_intr_exce_ret = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  reg_id2wb_fencei = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  reg_id2wb_wb_sel = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  reg_id2wb_regfile_we_en = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  reg_id2wb_regfile_we_addr = _RAND_75[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_ChiselMDU(
  input         clock,
  input         reset,
  input         io_mdu_op_mul_signed,
  input         io_mdu_op_is_mu,
  input         io_mdu_op_mul_32,
  input  [1:0]  io_mdu_op_div_signed,
  input         io_mdu_op_is_div,
  input         io_mdu_op_is_du,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  output [63:0] io_result,
  output        io_ready
);
  wire  muler_clock; // @[MDU.scala 197:29]
  wire  muler_reset; // @[MDU.scala 197:29]
  wire  muler_in_valid; // @[MDU.scala 197:29]
  wire [1:0] muler_mul_signed; // @[MDU.scala 197:29]
  wire [63:0] muler_multiplicand; // @[MDU.scala 197:29]
  wire [63:0] muler_multiplier; // @[MDU.scala 197:29]
  wire  muler_out_valid; // @[MDU.scala 197:29]
  wire [63:0] muler_result_hi; // @[MDU.scala 197:29]
  wire [63:0] muler_result_lo; // @[MDU.scala 197:29]
  wire  diver_clock; // @[MDU.scala 198:29]
  wire  diver_reset; // @[MDU.scala 198:29]
  wire  diver_in_valid; // @[MDU.scala 198:29]
  wire  diver_div_signed; // @[MDU.scala 198:29]
  wire [63:0] diver_dividend; // @[MDU.scala 198:29]
  wire [63:0] diver_divisor; // @[MDU.scala 198:29]
  wire  diver_out_valid; // @[MDU.scala 198:29]
  wire [63:0] diver_quotient; // @[MDU.scala 198:29]
  wire [63:0] diver_remainder; // @[MDU.scala 198:29]
  wire [63:0] diver_res = io_mdu_op_is_div ? diver_quotient : diver_remainder; // @[MDU.scala 202:30]
  wire [63:0] muler_res = io_mdu_op_mul_32 ? muler_result_lo : muler_result_hi; // @[MDU.scala 211:30]
  ysyx_040978_muler muler ( // @[MDU.scala 197:29]
    .clock(muler_clock),
    .reset(muler_reset),
    .in_valid(muler_in_valid),
    .mul_signed(muler_mul_signed),
    .multiplicand(muler_multiplicand),
    .multiplier(muler_multiplier),
    .out_valid(muler_out_valid),
    .result_hi(muler_result_hi),
    .result_lo(muler_result_lo)
  );
  ysyx_040978_diver diver ( // @[MDU.scala 198:29]
    .clock(diver_clock),
    .reset(diver_reset),
    .in_valid(diver_in_valid),
    .div_signed(diver_div_signed),
    .dividend(diver_dividend),
    .divisor(diver_divisor),
    .out_valid(diver_out_valid),
    .quotient(diver_quotient),
    .remainder(diver_remainder)
  );
  assign io_result = io_mdu_op_is_du ? diver_res : muler_res; // @[MDU.scala 218:19]
  assign io_ready = muler_out_valid | diver_out_valid | ~(io_mdu_op_is_du | io_mdu_op_is_mu); // @[MDU.scala 219:41]
  assign muler_clock = clock; // @[MDU.scala 209:18]
  assign muler_reset = reset; // @[MDU.scala 210:18]
  assign muler_in_valid = io_mdu_op_is_mu & ~muler_out_valid; // @[MDU.scala 213:37]
  assign muler_mul_signed = {{1'd0}, io_mdu_op_mul_signed}; // @[MDU.scala 214:23]
  assign muler_multiplicand = io_src1; // @[MDU.scala 215:25]
  assign muler_multiplier = io_src2; // @[MDU.scala 216:23]
  assign diver_clock = clock; // @[MDU.scala 200:18]
  assign diver_reset = reset; // @[MDU.scala 201:18]
  assign diver_in_valid = io_mdu_op_is_du & ~diver_out_valid; // @[MDU.scala 204:37]
  assign diver_div_signed = io_mdu_op_div_signed[0]; // @[MDU.scala 205:23]
  assign diver_dividend = io_src1; // @[MDU.scala 206:21]
  assign diver_divisor = io_src2; // @[MDU.scala 207:20]
endmodule
module ysyx_040978_MDU(
  input         clock,
  input         reset,
  input         io_mdu_op_mul_signed,
  input         io_mdu_op_is_mu,
  input         io_mdu_op_mul_32,
  input  [1:0]  io_mdu_op_div_signed,
  input         io_mdu_op_is_div,
  input         io_mdu_op_is_du,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  output [63:0] io_result,
  output        io_ready
);
  wire  mdu_clock; // @[MDU.scala 105:21]
  wire  mdu_reset; // @[MDU.scala 105:21]
  wire  mdu_io_mdu_op_mul_signed; // @[MDU.scala 105:21]
  wire  mdu_io_mdu_op_is_mu; // @[MDU.scala 105:21]
  wire  mdu_io_mdu_op_mul_32; // @[MDU.scala 105:21]
  wire [1:0] mdu_io_mdu_op_div_signed; // @[MDU.scala 105:21]
  wire  mdu_io_mdu_op_is_div; // @[MDU.scala 105:21]
  wire  mdu_io_mdu_op_is_du; // @[MDU.scala 105:21]
  wire [63:0] mdu_io_src1; // @[MDU.scala 105:21]
  wire [63:0] mdu_io_src2; // @[MDU.scala 105:21]
  wire [63:0] mdu_io_result; // @[MDU.scala 105:21]
  wire  mdu_io_ready; // @[MDU.scala 105:21]
  ysyx_040978_ChiselMDU mdu ( // @[MDU.scala 105:21]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_mdu_op_mul_signed(mdu_io_mdu_op_mul_signed),
    .io_mdu_op_is_mu(mdu_io_mdu_op_is_mu),
    .io_mdu_op_mul_32(mdu_io_mdu_op_mul_32),
    .io_mdu_op_div_signed(mdu_io_mdu_op_div_signed),
    .io_mdu_op_is_div(mdu_io_mdu_op_is_div),
    .io_mdu_op_is_du(mdu_io_mdu_op_is_du),
    .io_src1(mdu_io_src1),
    .io_src2(mdu_io_src2),
    .io_result(mdu_io_result),
    .io_ready(mdu_io_ready)
  );
  assign io_result = mdu_io_result; // @[MDU.scala 106:12]
  assign io_ready = mdu_io_ready; // @[MDU.scala 106:12]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_mdu_op_mul_signed = io_mdu_op_mul_signed; // @[MDU.scala 106:12]
  assign mdu_io_mdu_op_is_mu = io_mdu_op_is_mu; // @[MDU.scala 106:12]
  assign mdu_io_mdu_op_mul_32 = io_mdu_op_mul_32; // @[MDU.scala 106:12]
  assign mdu_io_mdu_op_div_signed = io_mdu_op_div_signed; // @[MDU.scala 106:12]
  assign mdu_io_mdu_op_is_div = io_mdu_op_is_div; // @[MDU.scala 106:12]
  assign mdu_io_mdu_op_is_du = io_mdu_op_is_du; // @[MDU.scala 106:12]
  assign mdu_io_src1 = io_src1; // @[MDU.scala 106:12]
  assign mdu_io_src2 = io_src2; // @[MDU.scala 106:12]
endmodule
module ysyx_040978_CSRU(
  input         clock,
  input         reset,
  input         io_exu_csr_we,
  input         io_exu_csr_hit_is_mepc,
  input         io_exu_csr_hit_is_mtvec,
  input         io_exu_csr_hit_is_mstatus,
  input         io_exu_csr_hit_is_mie,
  input         io_exu_csr_hit_is_mcause,
  input         io_exu_csr_hit_is_mip,
  input         io_exu_csr_hit_is_mtime,
  input         io_exu_csr_hit_is_mcycle,
  input         io_exu_csr_hit_is_mhartid,
  input  [63:0] io_exu_rs1_data,
  input  [63:0] io_exu_zimm,
  input         io_exu_operator_csrrw,
  input         io_exu_operator_csrrs,
  input         io_exu_operator_csrrc,
  input         io_exu_operator_csrrwi,
  input         io_exu_operator_csrrsi,
  input         io_exu_operator_csrrci,
  output [63:0] io_exu_result,
  input         io_exu_intr,
  input         io_exu_exec,
  input         io_exu_mret,
  input  [3:0]  io_exu_exce_code,
  input  [63:0] io_exu_pc,
  output [63:0] io_ctrl_out_mepc,
  output [63:0] io_ctrl_out_mtvec,
  output        io_ctrl_out_mie,
  output        io_ctrl_out_mtie,
  output        io_ctrl_out_msie,
  output        io_ctrl_out_meie,
  output        io_ctrl_out_mtip,
  output        io_ctrl_out_msip,
  output        io_ctrl_out_meip,
  input         io_sb_clint_msip,
  input         io_sb_clint_mtip,
  input  [63:0] io_sb_clint_mtime,
  input         io_sb_meip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mcycle; // @[CSRU.scala 182:31]
  reg [63:0] mcause; // @[CSRU.scala 151:31]
  reg [63:0] mie; // @[CSRU.scala 141:28]
  reg [63:0] mstatus; // @[CSRU.scala 116:32]
  reg [63:0] mtvec; // @[CSRU.scala 104:30]
  reg [63:0] mepc; // @[CSRU.scala 94:29]
  wire [63:0] _GEN_0 = io_exu_csr_hit_is_mepc ? mepc : 64'h0; // @[CSRU.scala 96:29 CSRU.scala 96:41]
  wire [63:0] _GEN_3 = io_exu_csr_hit_is_mtvec ? mtvec : _GEN_0; // @[CSRU.scala 106:29 CSRU.scala 106:41]
  wire [63:0] _GEN_5 = io_exu_csr_hit_is_mstatus ? mstatus : _GEN_3; // @[CSRU.scala 123:31 CSRU.scala 123:43]
  wire [63:0] _GEN_15 = io_exu_csr_hit_is_mie ? mie : _GEN_5; // @[CSRU.scala 143:27 CSRU.scala 143:39]
  wire [63:0] _GEN_17 = io_exu_csr_hit_is_mcause ? mcause : _GEN_15; // @[CSRU.scala 153:22 CSRU.scala 153:34]
  wire [63:0] _GEN_20 = io_exu_csr_hit_is_mip ? 64'h0 : _GEN_17; // @[CSRU.scala 166:18 CSRU.scala 166:30]
  wire [63:0] _GEN_21 = io_exu_csr_hit_is_mtime ? io_sb_clint_mtime : _GEN_20; // @[CSRU.scala 178:19 CSRU.scala 178:31]
  wire [63:0] _GEN_22 = io_exu_csr_hit_is_mcycle ? mcycle : _GEN_21; // @[CSRU.scala 185:20 CSRU.scala 185:32]
  wire [63:0] csr_rdata = io_exu_csr_hit_is_mhartid ? 64'h0 : _GEN_22; // @[CSRU.scala 189:27 CSRU.scala 189:39]
  wire [63:0] _csr_wdata_T = csr_rdata | io_exu_rs1_data; // @[CSRU.scala 83:26]
  wire [63:0] _csr_wdata_T_1 = ~io_exu_rs1_data; // @[CSRU.scala 84:29]
  wire [63:0] _csr_wdata_T_2 = csr_rdata & _csr_wdata_T_1; // @[CSRU.scala 84:26]
  wire [58:0] csr_wdata_hi = csr_rdata[63:5]; // @[CSRU.scala 86:28]
  wire [4:0] csr_wdata_lo = csr_rdata[4:0] | io_exu_zimm[4:0]; // @[CSRU.scala 86:52]
  wire [63:0] _csr_wdata_T_5 = {csr_wdata_hi,csr_wdata_lo}; // @[Cat.scala 30:58]
  wire [4:0] _csr_wdata_T_8 = ~io_exu_zimm[4:0]; // @[CSRU.scala 87:55]
  wire [4:0] csr_wdata_lo_1 = csr_rdata[4:0] & _csr_wdata_T_8; // @[CSRU.scala 87:52]
  wire [63:0] _csr_wdata_T_9 = {csr_wdata_hi,csr_wdata_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _csr_wdata_T_10 = io_exu_operator_csrrci ? _csr_wdata_T_9 : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _csr_wdata_T_11 = io_exu_operator_csrrsi ? _csr_wdata_T_5 : _csr_wdata_T_10; // @[Mux.scala 98:16]
  wire [63:0] _csr_wdata_T_12 = io_exu_operator_csrrwi ? io_exu_zimm : _csr_wdata_T_11; // @[Mux.scala 98:16]
  wire [63:0] _csr_wdata_T_13 = io_exu_operator_csrrc ? _csr_wdata_T_2 : _csr_wdata_T_12; // @[Mux.scala 98:16]
  wire [63:0] _csr_wdata_T_14 = io_exu_operator_csrrs ? _csr_wdata_T : _csr_wdata_T_13; // @[Mux.scala 98:16]
  wire [63:0] csr_wdata = io_exu_operator_csrrw ? io_exu_rs1_data : _csr_wdata_T_14; // @[Mux.scala 98:16]
  wire  _T_1 = io_exu_intr | io_exu_exec; // @[CSRU.scala 99:24]
  wire [61:0] mtvec_hi = csr_wdata[63:2]; // @[CSRU.scala 107:53]
  wire [63:0] _mtvec_T = {mtvec_hi,2'h0}; // @[Cat.scala 30:58]
  wire [1:0] mstatus_in_hi_hi_lo = mstatus[12:11]; // @[CSRU.scala 119:29]
  wire [50:0] mstatus_in_hi_hi_hi = mstatus[63:13]; // @[CSRU.scala 120:28]
  wire [2:0] mstatus_in_hi_lo_hi = mstatus[10:8]; // @[CSRU.scala 120:61]
  wire [2:0] mstatus_in_lo_hi_hi = mstatus[6:4]; // @[CSRU.scala 120:94]
  wire [2:0] mstatus_in_lo_lo = mstatus[2:0]; // @[CSRU.scala 120:125]
  wire  _T_3 = io_exu_csr_hit_is_mstatus & io_exu_csr_we; // @[CSRU.scala 124:21]
  wire  _GEN_6 = io_exu_mret ? mstatus[7] : mstatus[3]; // @[CSRU.scala 134:24 CSRU.scala 135:22 CSRU.scala 117:19]
  wire  _GEN_8 = _T_1 ? 1'h0 : _GEN_6; // @[CSRU.scala 130:36 CSRU.scala 132:20]
  wire  _GEN_11 = _T_3 & _T_1 ? 1'h0 : _GEN_8; // @[CSRU.scala 126:62 CSRU.scala 129:19]
  wire  mstatus_in_lo_hi_lo = io_exu_csr_hit_is_mstatus & io_exu_csr_we & ~_T_1 ? mstatus[3] : _GEN_11; // @[CSRU.scala 124:56 CSRU.scala 117:19]
  wire  _GEN_7 = _T_1 ? mstatus[3] : mstatus[7]; // @[CSRU.scala 130:36 CSRU.scala 131:21 CSRU.scala 118:19]
  wire  _GEN_10 = _T_3 & _T_1 ? mstatus[3] : _GEN_7; // @[CSRU.scala 126:62 CSRU.scala 128:20]
  wire  mstatus_in_hi_lo_lo = io_exu_csr_hit_is_mstatus & io_exu_csr_we & ~_T_1 ? mstatus[7] : _GEN_10; // @[CSRU.scala 124:56 CSRU.scala 118:19]
  wire [63:0] _mstatus_in_T = {mstatus_in_hi_hi_hi,mstatus_in_hi_hi_lo,mstatus_in_hi_lo_hi,mstatus_in_hi_lo_lo,
    mstatus_in_lo_hi_hi,mstatus_in_lo_hi_lo,mstatus_in_lo_lo}; // @[Cat.scala 30:58]
  wire [31:0] mstatus_in_hi_1 = mstatus[63:32]; // @[CSRU.scala 125:30]
  wire [31:0] mstatus_in_lo_1 = csr_wdata[31:0]; // @[CSRU.scala 125:49]
  wire [63:0] _mstatus_in_T_1 = {mstatus_in_hi_1,mstatus_in_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _mcause_T = {60'h800000000000000,io_exu_exce_code}; // @[Cat.scala 30:58]
  wire [63:0] _mcause_T_1 = {60'h0,io_exu_exce_code}; // @[Cat.scala 30:58]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[CSRU.scala 184:20]
  assign io_exu_result = io_exu_csr_hit_is_mhartid ? 64'h0 : _GEN_22; // @[CSRU.scala 189:27 CSRU.scala 189:39]
  assign io_ctrl_out_mepc = mepc; // @[CSRU.scala 100:15]
  assign io_ctrl_out_mtvec = mtvec; // @[CSRU.scala 108:16]
  assign io_ctrl_out_mie = mstatus[3]; // @[CSRU.scala 137:24]
  assign io_ctrl_out_mtie = mie[7]; // @[CSRU.scala 146:21]
  assign io_ctrl_out_msie = mie[3]; // @[CSRU.scala 145:21]
  assign io_ctrl_out_meie = mie[11]; // @[CSRU.scala 147:21]
  assign io_ctrl_out_mtip = io_sb_clint_mtip; // @[CSRU.scala 171:15]
  assign io_ctrl_out_msip = io_sb_clint_msip; // @[CSRU.scala 170:15]
  assign io_ctrl_out_meip = io_sb_meip; // @[CSRU.scala 172:15]
  always @(posedge clock) begin
    if (reset) begin // @[CSRU.scala 182:31]
      mcycle <= 64'h0; // @[CSRU.scala 182:31]
    end else begin
      mcycle <= _mcycle_T_1; // @[CSRU.scala 184:10]
    end
    if (reset) begin // @[CSRU.scala 151:31]
      mcause <= 64'h0; // @[CSRU.scala 151:31]
    end else if (io_exu_intr) begin // @[CSRU.scala 154:22]
      mcause <= _mcause_T; // @[CSRU.scala 154:31]
    end else if (io_exu_exec) begin // @[CSRU.scala 155:24]
      mcause <= _mcause_T_1; // @[CSRU.scala 155:33]
    end
    if (reset) begin // @[CSRU.scala 141:28]
      mie <= 64'h0; // @[CSRU.scala 141:28]
    end else if (io_exu_csr_hit_is_mie & io_exu_csr_we) begin // @[CSRU.scala 144:27]
      if (io_exu_operator_csrrw) begin // @[Mux.scala 98:16]
        mie <= io_exu_rs1_data;
      end else if (io_exu_operator_csrrs) begin // @[Mux.scala 98:16]
        mie <= _csr_wdata_T;
      end else begin
        mie <= _csr_wdata_T_13;
      end
    end
    if (reset) begin // @[CSRU.scala 116:32]
      mstatus <= 64'ha00000000; // @[CSRU.scala 116:32]
    end else if (io_exu_csr_hit_is_mstatus & io_exu_csr_we & ~_T_1) begin // @[CSRU.scala 124:56]
      mstatus <= _mstatus_in_T_1; // @[CSRU.scala 125:16]
    end else if (_T_3 & _T_1) begin // @[CSRU.scala 126:62]
      mstatus <= _mstatus_in_T_1; // @[CSRU.scala 127:16]
    end else begin
      mstatus <= _mstatus_in_T; // @[CSRU.scala 120:14]
    end
    if (reset) begin // @[CSRU.scala 104:30]
      mtvec <= 64'h0; // @[CSRU.scala 104:30]
    end else if (io_exu_csr_hit_is_mtvec & io_exu_csr_we) begin // @[CSRU.scala 107:29]
      mtvec <= _mtvec_T; // @[CSRU.scala 107:37]
    end
    if (reset) begin // @[CSRU.scala 94:29]
      mepc <= 64'h0; // @[CSRU.scala 94:29]
    end else if (io_exu_csr_hit_is_mepc & io_exu_csr_we) begin // @[CSRU.scala 98:30]
      if (io_exu_operator_csrrw) begin // @[Mux.scala 98:16]
        mepc <= io_exu_rs1_data;
      end else if (io_exu_operator_csrrs) begin // @[Mux.scala 98:16]
        mepc <= _csr_wdata_T;
      end else begin
        mepc <= _csr_wdata_T_13;
      end
    end else if (io_exu_intr | io_exu_exec) begin // @[CSRU.scala 99:36]
      mepc <= io_exu_pc; // @[CSRU.scala 99:43]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mcycle = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcause = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mie = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatus = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtvec = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mepc = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_EXU(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [63:0] io_prev_bits_id2ex_alu_src1,
  input  [63:0] io_prev_bits_id2ex_alu_src2,
  input  [63:0] io_prev_bits_id2ex_salu_src1,
  input  [63:0] io_prev_bits_id2ex_salu_src2,
  input  [63:0] io_prev_bits_id2ex_src1,
  input  [63:0] io_prev_bits_id2ex_src2,
  input  [63:0] io_prev_bits_id2ex_src3,
  input         io_prev_bits_id2ex_operator_auipc,
  input         io_prev_bits_id2ex_operator_lui,
  input         io_prev_bits_id2ex_operator_jal,
  input         io_prev_bits_id2ex_operator_jalr,
  input         io_prev_bits_id2ex_operator_sb,
  input         io_prev_bits_id2ex_operator_sh,
  input         io_prev_bits_id2ex_operator_sw,
  input         io_prev_bits_id2ex_operator_sd,
  input         io_prev_bits_id2ex_operator_add,
  input         io_prev_bits_id2ex_operator_sub,
  input         io_prev_bits_id2ex_operator_sll,
  input         io_prev_bits_id2ex_operator_slt,
  input         io_prev_bits_id2ex_operator_sltu,
  input         io_prev_bits_id2ex_operator_xor,
  input         io_prev_bits_id2ex_operator_srl,
  input         io_prev_bits_id2ex_operator_sra,
  input         io_prev_bits_id2ex_operator_or,
  input         io_prev_bits_id2ex_operator_and,
  input         io_prev_bits_id2ex_operator_csr_is_csr,
  input         io_prev_bits_id2ex_operator_csr_csrrw,
  input         io_prev_bits_id2ex_operator_csr_csrrs,
  input         io_prev_bits_id2ex_operator_csr_csrrc,
  input         io_prev_bits_id2ex_operator_csr_csrrwi,
  input         io_prev_bits_id2ex_operator_csr_csrrsi,
  input         io_prev_bits_id2ex_operator_csr_csrrci,
  input         io_prev_bits_id2ex_srcsize_byte,
  input         io_prev_bits_id2ex_srcsize_hword,
  input         io_prev_bits_id2ex_srcsize_word,
  input         io_prev_bits_id2ex_srcsize_dword,
  input         io_prev_bits_id2ex_is_load,
  input         io_prev_bits_id2ex_is_save,
  input         io_prev_bits_id2ex_div_inf,
  input         io_prev_bits_id2ex_csr_we,
  input         io_prev_bits_id2ex_csr_hit_is_mepc,
  input         io_prev_bits_id2ex_csr_hit_is_mtvec,
  input         io_prev_bits_id2ex_csr_hit_is_mstatus,
  input         io_prev_bits_id2ex_csr_hit_is_mie,
  input         io_prev_bits_id2ex_csr_hit_is_mcause,
  input         io_prev_bits_id2ex_csr_hit_is_mip,
  input         io_prev_bits_id2ex_csr_hit_is_mtime,
  input         io_prev_bits_id2ex_csr_hit_is_mcycle,
  input         io_prev_bits_id2ex_csr_hit_is_mhartid,
  input         io_prev_bits_id2ex_mdu_op_mul_signed,
  input         io_prev_bits_id2ex_mdu_op_is_mu,
  input         io_prev_bits_id2ex_mdu_op_mul_32,
  input  [1:0]  io_prev_bits_id2ex_mdu_op_div_signed,
  input         io_prev_bits_id2ex_mdu_op_is_div,
  input         io_prev_bits_id2ex_mdu_op_is_du,
  input  [4:0]  io_prev_bits_id2ex_zimm,
  input         io_prev_bits_id2ex_intr,
  input         io_prev_bits_id2ex_exec,
  input         io_prev_bits_id2ex_mret,
  input  [3:0]  io_prev_bits_id2ex_exce_code,
  input  [63:0] io_prev_bits_id2ex_pc,
  input         io_prev_bits_id2ex_is_iem,
  input         io_prev_bits_id2mem_fencei,
  input         io_prev_bits_id2mem_size_byte,
  input         io_prev_bits_id2mem_size_hword,
  input         io_prev_bits_id2mem_size_word,
  input         io_prev_bits_id2mem_size_dword,
  input         io_prev_bits_id2mem_sext_flag,
  input         io_prev_bits_id2mem_memory_rd_en,
  input         io_prev_bits_id2mem_memory_we_en,
  input         io_prev_bits_id2wb_intr_exce_ret,
  input         io_prev_bits_id2wb_fencei,
  input         io_prev_bits_id2wb_wb_sel,
  input         io_prev_bits_id2wb_regfile_we_en,
  input  [4:0]  io_prev_bits_id2wb_regfile_we_addr,
  input         io_next_ready,
  output        io_next_valid,
  output        io_next_bits_id2mem_fencei,
  output        io_next_bits_id2mem_size_byte,
  output        io_next_bits_id2mem_size_hword,
  output        io_next_bits_id2mem_size_word,
  output        io_next_bits_id2mem_size_dword,
  output        io_next_bits_id2mem_sext_flag,
  output        io_next_bits_id2mem_memory_rd_en,
  output        io_next_bits_id2mem_memory_we_en,
  output        io_next_bits_id2wb_intr_exce_ret,
  output        io_next_bits_id2wb_fencei,
  output        io_next_bits_id2wb_wb_sel,
  output        io_next_bits_id2wb_regfile_we_en,
  output [4:0]  io_next_bits_id2wb_regfile_we_addr,
  output [38:0] io_next_bits_ex2mem_addr,
  output [63:0] io_next_bits_ex2mem_we_data,
  output [7:0]  io_next_bits_ex2mem_we_mask,
  output [63:0] io_next_bits_ex2wb_result_data,
  output [63:0] io_csr2ctrl_out_mepc,
  output [63:0] io_csr2ctrl_out_mtvec,
  output        io_csr2ctrl_out_mie,
  output        io_csr2ctrl_out_mtie,
  output        io_csr2ctrl_out_msie,
  output        io_csr2ctrl_out_meie,
  output        io_csr2ctrl_out_mtip,
  output        io_csr2ctrl_out_msip,
  output        io_csr2ctrl_out_meip,
  input         io_sb_clint_msip,
  input         io_sb_clint_mtip,
  input  [63:0] io_sb_clint_mtime,
  input         io_sb_meip
);
  wire  mdu_clock; // @[EXU.scala 57:27]
  wire  mdu_reset; // @[EXU.scala 57:27]
  wire  mdu_io_mdu_op_mul_signed; // @[EXU.scala 57:27]
  wire  mdu_io_mdu_op_is_mu; // @[EXU.scala 57:27]
  wire  mdu_io_mdu_op_mul_32; // @[EXU.scala 57:27]
  wire [1:0] mdu_io_mdu_op_div_signed; // @[EXU.scala 57:27]
  wire  mdu_io_mdu_op_is_div; // @[EXU.scala 57:27]
  wire  mdu_io_mdu_op_is_du; // @[EXU.scala 57:27]
  wire [63:0] mdu_io_src1; // @[EXU.scala 57:27]
  wire [63:0] mdu_io_src2; // @[EXU.scala 57:27]
  wire [63:0] mdu_io_result; // @[EXU.scala 57:27]
  wire  mdu_io_ready; // @[EXU.scala 57:27]
  wire  csru_clock; // @[EXU.scala 116:28]
  wire  csru_reset; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_we; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mepc; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mtvec; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mstatus; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mie; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mcause; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mip; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mtime; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mcycle; // @[EXU.scala 116:28]
  wire  csru_io_exu_csr_hit_is_mhartid; // @[EXU.scala 116:28]
  wire [63:0] csru_io_exu_rs1_data; // @[EXU.scala 116:28]
  wire [63:0] csru_io_exu_zimm; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrw; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrs; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrc; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrwi; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrsi; // @[EXU.scala 116:28]
  wire  csru_io_exu_operator_csrrci; // @[EXU.scala 116:28]
  wire [63:0] csru_io_exu_result; // @[EXU.scala 116:28]
  wire  csru_io_exu_intr; // @[EXU.scala 116:28]
  wire  csru_io_exu_exec; // @[EXU.scala 116:28]
  wire  csru_io_exu_mret; // @[EXU.scala 116:28]
  wire [3:0] csru_io_exu_exce_code; // @[EXU.scala 116:28]
  wire [63:0] csru_io_exu_pc; // @[EXU.scala 116:28]
  wire [63:0] csru_io_ctrl_out_mepc; // @[EXU.scala 116:28]
  wire [63:0] csru_io_ctrl_out_mtvec; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_mie; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_mtie; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_msie; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_meie; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_mtip; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_msip; // @[EXU.scala 116:28]
  wire  csru_io_ctrl_out_meip; // @[EXU.scala 116:28]
  wire  csru_io_sb_clint_msip; // @[EXU.scala 116:28]
  wire  csru_io_sb_clint_mtip; // @[EXU.scala 116:28]
  wire [63:0] csru_io_sb_clint_mtime; // @[EXU.scala 116:28]
  wire  csru_io_sb_meip; // @[EXU.scala 116:28]
  wire [5:0] shift_src2 = io_prev_bits_id2ex_srcsize_word ? {{1'd0}, io_prev_bits_id2ex_src2[4:0]} :
    io_prev_bits_id2ex_src2[5:0]; // @[EXU.scala 55:31]
  wire [63:0] mdu_result = io_prev_bits_id2ex_div_inf ? 64'hffffffffffffffff : mdu_io_result; // @[EXU.scala 60:31]
  wire [126:0] _GEN_22 = {{63'd0}, io_prev_bits_id2ex_alu_src1}; // @[EXU.scala 65:28]
  wire [126:0] _result_sll_T = _GEN_22 << shift_src2; // @[EXU.scala 65:28]
  wire [63:0] result_srl = io_prev_bits_id2ex_alu_src1 >> shift_src2; // @[EXU.scala 67:27]
  wire [63:0] add_src1_src3 = io_prev_bits_id2ex_src1 + io_prev_bits_id2ex_src3; // @[EXU.scala 70:36]
  wire  _result_T = io_prev_bits_id2ex_operator_jal | io_prev_bits_id2ex_operator_jalr; // @[EXU.scala 75:21]
  wire [63:0] _result_T_2 = 64'h4 + io_prev_bits_id2ex_src3; // @[EXU.scala 75:46]
  wire [63:0] _result_T_4 = io_prev_bits_id2ex_alu_src1 - io_prev_bits_id2ex_alu_src2; // @[EXU.scala 80:38]
  wire [63:0] _result_T_6 = io_prev_bits_id2ex_alu_src1 + io_prev_bits_id2ex_alu_src2; // @[EXU.scala 81:38]
  wire [63:0] _result_T_7 = io_prev_bits_id2ex_alu_src1 ^ io_prev_bits_id2ex_alu_src2; // @[EXU.scala 82:38]
  wire [63:0] _result_T_8 = io_prev_bits_id2ex_alu_src1 | io_prev_bits_id2ex_alu_src2; // @[EXU.scala 83:38]
  wire [63:0] _result_T_9 = io_prev_bits_id2ex_alu_src1 & io_prev_bits_id2ex_alu_src2; // @[EXU.scala 84:38]
  wire  _result_T_10 = $signed(io_prev_bits_id2ex_salu_src1) < $signed(io_prev_bits_id2ex_salu_src2); // @[EXU.scala 85:39]
  wire  _result_T_11 = io_prev_bits_id2ex_alu_src1 < io_prev_bits_id2ex_alu_src2; // @[EXU.scala 86:38]
  wire [63:0] _result_T_12 = $signed(io_prev_bits_id2ex_salu_src1) >>> shift_src2; // @[EXU.scala 89:39]
  wire [63:0] _result_T_13 = io_prev_bits_id2ex_operator_sra ? _result_T_12 : mdu_result; // @[Mux.scala 98:16]
  wire [63:0] _result_T_14 = io_prev_bits_id2ex_operator_srl ? result_srl : _result_T_13; // @[Mux.scala 98:16]
  wire [63:0] result_sll = _result_sll_T[63:0]; // @[EXU.scala 64:32 EXU.scala 65:14]
  wire [63:0] _result_T_15 = io_prev_bits_id2ex_operator_sll ? result_sll : _result_T_14; // @[Mux.scala 98:16]
  wire [63:0] _result_T_16 = io_prev_bits_id2ex_operator_sltu ? {{63'd0}, _result_T_11} : _result_T_15; // @[Mux.scala 98:16]
  wire [63:0] _result_T_17 = io_prev_bits_id2ex_operator_slt ? {{63'd0}, _result_T_10} : _result_T_16; // @[Mux.scala 98:16]
  wire [63:0] _result_T_18 = io_prev_bits_id2ex_operator_and ? _result_T_9 : _result_T_17; // @[Mux.scala 98:16]
  wire [63:0] _result_T_19 = io_prev_bits_id2ex_operator_or ? _result_T_8 : _result_T_18; // @[Mux.scala 98:16]
  wire [63:0] _result_T_20 = io_prev_bits_id2ex_operator_xor ? _result_T_7 : _result_T_19; // @[Mux.scala 98:16]
  wire [63:0] _result_T_21 = io_prev_bits_id2ex_operator_add ? _result_T_6 : _result_T_20; // @[Mux.scala 98:16]
  wire [63:0] _result_T_22 = io_prev_bits_id2ex_operator_sub ? _result_T_4 : _result_T_21; // @[Mux.scala 98:16]
  wire [63:0] _result_T_23 = io_prev_bits_id2ex_operator_sd ? io_prev_bits_id2ex_src2 : _result_T_22; // @[Mux.scala 98:16]
  wire [63:0] _result_T_24 = io_prev_bits_id2ex_operator_sw ? io_prev_bits_id2ex_src2 : _result_T_23; // @[Mux.scala 98:16]
  wire [63:0] _result_T_25 = io_prev_bits_id2ex_operator_sh ? io_prev_bits_id2ex_src2 : _result_T_24; // @[Mux.scala 98:16]
  wire [63:0] _result_T_26 = io_prev_bits_id2ex_operator_sb ? io_prev_bits_id2ex_src2 : _result_T_25; // @[Mux.scala 98:16]
  wire [63:0] _result_T_27 = _result_T ? _result_T_2 : _result_T_26; // @[Mux.scala 98:16]
  wire [63:0] _result_T_28 = io_prev_bits_id2ex_operator_lui ? io_prev_bits_id2ex_src1 : _result_T_27; // @[Mux.scala 98:16]
  wire [63:0] result = io_prev_bits_id2ex_operator_auipc ? add_src1_src3 : _result_T_28; // @[Mux.scala 98:16]
  wire [7:0] _result_out_signed_T_1 = result[7:0]; // @[EXU.scala 95:29]
  wire [15:0] _result_out_signed_T_3 = result[15:0]; // @[EXU.scala 96:30]
  wire [31:0] _result_out_signed_T_5 = result[31:0]; // @[EXU.scala 97:30]
  wire [63:0] _result_out_signed_T_7 = io_prev_bits_id2ex_operator_auipc ? add_src1_src3 : _result_T_28; // @[EXU.scala 98:30]
  wire [63:0] _result_out_signed_T_8 = io_prev_bits_id2ex_srcsize_dword ? $signed(_result_out_signed_T_7) : $signed(64'sh0
    ); // @[Mux.scala 98:16]
  wire [63:0] _result_out_signed_T_9 = io_prev_bits_id2ex_srcsize_word ? $signed({{32{_result_out_signed_T_5[31]}},
    _result_out_signed_T_5}) : $signed(_result_out_signed_T_8); // @[Mux.scala 98:16]
  wire [63:0] _result_out_signed_T_10 = io_prev_bits_id2ex_srcsize_hword ? $signed({{48{_result_out_signed_T_3[15]}},
    _result_out_signed_T_3}) : $signed(_result_out_signed_T_9); // @[Mux.scala 98:16]
  wire [63:0] _result_out_T = io_prev_bits_id2ex_srcsize_byte ? $signed({{56{_result_out_signed_T_1[7]}},
    _result_out_signed_T_1}) : $signed(_result_out_signed_T_10); // @[EXU.scala 101:65]
  wire [63:0] result_out = io_prev_bits_id2ex_srcsize_dword ? result : _result_out_T; // @[EXU.scala 101:31]
  wire [38:0] _io_next_bits_ex2mem_addr_T_4 = io_prev_bits_id2ex_src1[38:0] + io_prev_bits_id2ex_src2[38:0]; // @[EXU.scala 105:32]
  wire [38:0] _io_next_bits_ex2mem_addr_T_5 = io_prev_bits_id2ex_is_load ? _io_next_bits_ex2mem_addr_T_4 : 39'h0; // @[Mux.scala 98:16]
  wire [38:0] _io_next_bits_ex2mem_addr_T_6 = io_prev_bits_id2ex_is_save ? add_src1_src3[38:0] :
    _io_next_bits_ex2mem_addr_T_5; // @[Mux.scala 98:16]
  wire [7:0] _io_next_bits_ex2mem_we_mask_T = io_prev_bits_id2ex_srcsize_dword ? 8'hff : 8'h0; // @[Mux.scala 98:16]
  wire [7:0] _io_next_bits_ex2mem_we_mask_T_1 = io_prev_bits_id2ex_srcsize_word ? 8'hf : _io_next_bits_ex2mem_we_mask_T; // @[Mux.scala 98:16]
  wire [7:0] _io_next_bits_ex2mem_we_mask_T_2 = io_prev_bits_id2ex_srcsize_hword ? 8'h3 :
    _io_next_bits_ex2mem_we_mask_T_1; // @[Mux.scala 98:16]
  wire [7:0] _io_next_bits_ex2mem_we_mask_T_3 = io_prev_bits_id2ex_srcsize_byte ? 8'h1 :
    _io_next_bits_ex2mem_we_mask_T_2; // @[Mux.scala 98:16]
  wire [63:0] _GEN_0 = io_prev_bits_id2ex_operator_csr_is_csr ? csru_io_exu_result : result_out; // @[EXU.scala 131:28 EXU.scala 131:46 EXU.scala 114:19]
  ysyx_040978_MDU mdu ( // @[EXU.scala 57:27]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_mdu_op_mul_signed(mdu_io_mdu_op_mul_signed),
    .io_mdu_op_is_mu(mdu_io_mdu_op_is_mu),
    .io_mdu_op_mul_32(mdu_io_mdu_op_mul_32),
    .io_mdu_op_div_signed(mdu_io_mdu_op_div_signed),
    .io_mdu_op_is_div(mdu_io_mdu_op_is_div),
    .io_mdu_op_is_du(mdu_io_mdu_op_is_du),
    .io_src1(mdu_io_src1),
    .io_src2(mdu_io_src2),
    .io_result(mdu_io_result),
    .io_ready(mdu_io_ready)
  );
  ysyx_040978_CSRU csru ( // @[EXU.scala 116:28]
    .clock(csru_clock),
    .reset(csru_reset),
    .io_exu_csr_we(csru_io_exu_csr_we),
    .io_exu_csr_hit_is_mepc(csru_io_exu_csr_hit_is_mepc),
    .io_exu_csr_hit_is_mtvec(csru_io_exu_csr_hit_is_mtvec),
    .io_exu_csr_hit_is_mstatus(csru_io_exu_csr_hit_is_mstatus),
    .io_exu_csr_hit_is_mie(csru_io_exu_csr_hit_is_mie),
    .io_exu_csr_hit_is_mcause(csru_io_exu_csr_hit_is_mcause),
    .io_exu_csr_hit_is_mip(csru_io_exu_csr_hit_is_mip),
    .io_exu_csr_hit_is_mtime(csru_io_exu_csr_hit_is_mtime),
    .io_exu_csr_hit_is_mcycle(csru_io_exu_csr_hit_is_mcycle),
    .io_exu_csr_hit_is_mhartid(csru_io_exu_csr_hit_is_mhartid),
    .io_exu_rs1_data(csru_io_exu_rs1_data),
    .io_exu_zimm(csru_io_exu_zimm),
    .io_exu_operator_csrrw(csru_io_exu_operator_csrrw),
    .io_exu_operator_csrrs(csru_io_exu_operator_csrrs),
    .io_exu_operator_csrrc(csru_io_exu_operator_csrrc),
    .io_exu_operator_csrrwi(csru_io_exu_operator_csrrwi),
    .io_exu_operator_csrrsi(csru_io_exu_operator_csrrsi),
    .io_exu_operator_csrrci(csru_io_exu_operator_csrrci),
    .io_exu_result(csru_io_exu_result),
    .io_exu_intr(csru_io_exu_intr),
    .io_exu_exec(csru_io_exu_exec),
    .io_exu_mret(csru_io_exu_mret),
    .io_exu_exce_code(csru_io_exu_exce_code),
    .io_exu_pc(csru_io_exu_pc),
    .io_ctrl_out_mepc(csru_io_ctrl_out_mepc),
    .io_ctrl_out_mtvec(csru_io_ctrl_out_mtvec),
    .io_ctrl_out_mie(csru_io_ctrl_out_mie),
    .io_ctrl_out_mtie(csru_io_ctrl_out_mtie),
    .io_ctrl_out_msie(csru_io_ctrl_out_msie),
    .io_ctrl_out_meie(csru_io_ctrl_out_meie),
    .io_ctrl_out_mtip(csru_io_ctrl_out_mtip),
    .io_ctrl_out_msip(csru_io_ctrl_out_msip),
    .io_ctrl_out_meip(csru_io_ctrl_out_meip),
    .io_sb_clint_msip(csru_io_sb_clint_msip),
    .io_sb_clint_mtip(csru_io_sb_clint_mtip),
    .io_sb_clint_mtime(csru_io_sb_clint_mtime),
    .io_sb_meip(csru_io_sb_meip)
  );
  assign io_prev_ready = io_next_ready & mdu_io_ready; // @[EXU.scala 137:34]
  assign io_next_valid = io_prev_valid & mdu_io_ready; // @[EXU.scala 138:34]
  assign io_next_bits_id2mem_fencei = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_fencei; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_size_byte = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_size_byte; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_size_hword = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_size_hword; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_size_word = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_size_word; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_size_dword = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_size_dword; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_sext_flag = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_sext_flag; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_memory_rd_en = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_memory_rd_en; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2mem_memory_we_en = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2mem_memory_we_en; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 34:23]
  assign io_next_bits_id2wb_intr_exce_ret = io_prev_bits_id2wb_intr_exce_ret; // @[EXU.scala 132:19 EXU.scala 134:38 EXU.scala 33:22]
  assign io_next_bits_id2wb_fencei = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2wb_fencei; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 33:22]
  assign io_next_bits_id2wb_wb_sel = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2wb_wb_sel; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 33:22]
  assign io_next_bits_id2wb_regfile_we_en = io_prev_bits_id2ex_is_iem ? 1'h0 : io_prev_bits_id2wb_regfile_we_en; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 33:22]
  assign io_next_bits_id2wb_regfile_we_addr = io_prev_bits_id2ex_is_iem ? 5'h0 : io_prev_bits_id2wb_regfile_we_addr; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 33:22]
  assign io_next_bits_ex2mem_addr = io_prev_bits_id2ex_is_iem ? 39'h0 : _io_next_bits_ex2mem_addr_T_6; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 103:13]
  assign io_next_bits_ex2mem_we_data = io_prev_bits_id2ex_is_iem ? 64'h0 : result_out; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 107:16]
  assign io_next_bits_ex2mem_we_mask = io_prev_bits_id2ex_is_iem ? 8'h0 : _io_next_bits_ex2mem_we_mask_T_3; // @[EXU.scala 132:19 EXU.scala 133:18 EXU.scala 108:16]
  assign io_next_bits_ex2wb_result_data = io_prev_bits_id2ex_is_iem ? 64'h0 : _GEN_0; // @[EXU.scala 132:19 EXU.scala 133:18]
  assign io_csr2ctrl_out_mepc = csru_io_ctrl_out_mepc; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_mtvec = csru_io_ctrl_out_mtvec; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_mie = csru_io_ctrl_out_mie; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_mtie = csru_io_ctrl_out_mtie; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_msie = csru_io_ctrl_out_msie; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_meie = csru_io_ctrl_out_meie; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_mtip = csru_io_ctrl_out_mtip; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_msip = csru_io_ctrl_out_msip; // @[EXU.scala 118:16]
  assign io_csr2ctrl_out_meip = csru_io_ctrl_out_meip; // @[EXU.scala 118:16]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_mdu_op_mul_signed = io_prev_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 61:17]
  assign mdu_io_mdu_op_is_mu = io_prev_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 61:17]
  assign mdu_io_mdu_op_mul_32 = io_prev_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 61:17]
  assign mdu_io_mdu_op_div_signed = io_prev_bits_id2ex_mdu_op_div_signed; // @[EXU.scala 61:17]
  assign mdu_io_mdu_op_is_div = io_prev_bits_id2ex_mdu_op_is_div; // @[EXU.scala 61:17]
  assign mdu_io_mdu_op_is_du = io_prev_bits_id2ex_mdu_op_is_du; // @[EXU.scala 61:17]
  assign mdu_io_src1 = io_prev_bits_id2ex_alu_src1; // @[EXU.scala 58:15]
  assign mdu_io_src2 = io_prev_bits_id2ex_alu_src2; // @[EXU.scala 59:15]
  assign csru_clock = clock;
  assign csru_reset = reset;
  assign csru_io_exu_csr_we = io_prev_bits_id2ex_csr_we; // @[EXU.scala 120:22]
  assign csru_io_exu_csr_hit_is_mepc = io_prev_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mtvec = io_prev_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mstatus = io_prev_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mie = io_prev_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mcause = io_prev_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mip = io_prev_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mtime = io_prev_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mcycle = io_prev_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 119:23]
  assign csru_io_exu_csr_hit_is_mhartid = io_prev_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 119:23]
  assign csru_io_exu_rs1_data = io_prev_bits_id2ex_src1; // @[EXU.scala 122:24]
  assign csru_io_exu_zimm = {{59'd0}, io_prev_bits_id2ex_zimm}; // @[EXU.scala 125:20]
  assign csru_io_exu_operator_csrrw = io_prev_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 121:24]
  assign csru_io_exu_operator_csrrs = io_prev_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 121:24]
  assign csru_io_exu_operator_csrrc = io_prev_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 121:24]
  assign csru_io_exu_operator_csrrwi = io_prev_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 121:24]
  assign csru_io_exu_operator_csrrsi = io_prev_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 121:24]
  assign csru_io_exu_operator_csrrci = io_prev_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 121:24]
  assign csru_io_exu_intr = io_prev_bits_id2ex_intr; // @[EXU.scala 126:20]
  assign csru_io_exu_exec = io_prev_bits_id2ex_exec; // @[EXU.scala 127:20]
  assign csru_io_exu_mret = io_prev_bits_id2ex_mret; // @[EXU.scala 128:20]
  assign csru_io_exu_exce_code = io_prev_bits_id2ex_exce_code; // @[EXU.scala 129:25]
  assign csru_io_exu_pc = io_prev_bits_id2ex_pc; // @[EXU.scala 130:18]
  assign csru_io_sb_clint_msip = io_sb_clint_msip; // @[EXU.scala 117:16]
  assign csru_io_sb_clint_mtip = io_sb_clint_mtip; // @[EXU.scala 117:16]
  assign csru_io_sb_clint_mtime = io_sb_clint_mtime; // @[EXU.scala 117:16]
  assign csru_io_sb_meip = io_sb_meip; // @[EXU.scala 117:16]
endmodule
module ysyx_040978_MEMReg(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input         io_prev_bits_id2mem_fencei,
  input         io_prev_bits_id2mem_size_byte,
  input         io_prev_bits_id2mem_size_hword,
  input         io_prev_bits_id2mem_size_word,
  input         io_prev_bits_id2mem_size_dword,
  input         io_prev_bits_id2mem_sext_flag,
  input         io_prev_bits_id2mem_memory_rd_en,
  input         io_prev_bits_id2mem_memory_we_en,
  input         io_prev_bits_id2wb_intr_exce_ret,
  input         io_prev_bits_id2wb_fencei,
  input         io_prev_bits_id2wb_wb_sel,
  input         io_prev_bits_id2wb_regfile_we_en,
  input  [4:0]  io_prev_bits_id2wb_regfile_we_addr,
  input  [38:0] io_prev_bits_ex2mem_addr,
  input  [63:0] io_prev_bits_ex2mem_we_data,
  input  [7:0]  io_prev_bits_ex2mem_we_mask,
  input  [63:0] io_prev_bits_ex2wb_result_data,
  input         io_next_ready,
  output        io_next_valid,
  output        io_next_bits_id2mem_fencei,
  output        io_next_bits_id2mem_size_byte,
  output        io_next_bits_id2mem_size_hword,
  output        io_next_bits_id2mem_size_word,
  output        io_next_bits_id2mem_size_dword,
  output        io_next_bits_id2mem_sext_flag,
  output        io_next_bits_id2mem_memory_rd_en,
  output        io_next_bits_id2mem_memory_we_en,
  output        io_next_bits_id2wb_intr_exce_ret,
  output        io_next_bits_id2wb_fencei,
  output        io_next_bits_id2wb_wb_sel,
  output        io_next_bits_id2wb_regfile_we_en,
  output [4:0]  io_next_bits_id2wb_regfile_we_addr,
  output [38:0] io_next_bits_ex2mem_addr,
  output [63:0] io_next_bits_ex2mem_we_data,
  output [7:0]  io_next_bits_ex2mem_we_mask,
  output [63:0] io_next_bits_ex2wb_result_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  io_next_valid_r; // @[Reg.scala 27:20]
  wire  data_id2mem_fencei = io_prev_valid & io_prev_bits_id2mem_fencei; // @[MEMU.scala 21:17]
  wire  data_id2mem_size_byte = io_prev_valid & io_prev_bits_id2mem_size_byte; // @[MEMU.scala 21:17]
  wire  data_id2mem_size_hword = io_prev_valid & io_prev_bits_id2mem_size_hword; // @[MEMU.scala 21:17]
  wire  data_id2mem_size_word = io_prev_valid & io_prev_bits_id2mem_size_word; // @[MEMU.scala 21:17]
  wire  data_id2mem_size_dword = io_prev_valid & io_prev_bits_id2mem_size_dword; // @[MEMU.scala 21:17]
  wire  data_id2mem_sext_flag = io_prev_valid & io_prev_bits_id2mem_sext_flag; // @[MEMU.scala 21:17]
  wire  data_id2mem_memory_rd_en = io_prev_valid & io_prev_bits_id2mem_memory_rd_en; // @[MEMU.scala 21:17]
  wire  data_id2mem_memory_we_en = io_prev_valid & io_prev_bits_id2mem_memory_we_en; // @[MEMU.scala 21:17]
  wire  data_id2wb_intr_exce_ret = io_prev_valid & io_prev_bits_id2wb_intr_exce_ret; // @[MEMU.scala 21:17]
  wire  data_id2wb_fencei = io_prev_valid & io_prev_bits_id2wb_fencei; // @[MEMU.scala 21:17]
  wire  data_id2wb_wb_sel = io_prev_valid & io_prev_bits_id2wb_wb_sel; // @[MEMU.scala 21:17]
  wire  data_id2wb_regfile_we_en = io_prev_valid & io_prev_bits_id2wb_regfile_we_en; // @[MEMU.scala 21:17]
  reg  reg_id2mem_fencei; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_byte; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_hword; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_word; // @[Reg.scala 27:20]
  reg  reg_id2mem_size_dword; // @[Reg.scala 27:20]
  reg  reg_id2mem_sext_flag; // @[Reg.scala 27:20]
  reg  reg_id2mem_memory_rd_en; // @[Reg.scala 27:20]
  reg  reg_id2mem_memory_we_en; // @[Reg.scala 27:20]
  reg  reg_id2wb_intr_exce_ret; // @[Reg.scala 27:20]
  reg  reg_id2wb_fencei; // @[Reg.scala 27:20]
  reg  reg_id2wb_wb_sel; // @[Reg.scala 27:20]
  reg  reg_id2wb_regfile_we_en; // @[Reg.scala 27:20]
  reg [4:0] reg_id2wb_regfile_we_addr; // @[Reg.scala 27:20]
  reg [38:0] reg_ex2mem_addr; // @[Reg.scala 27:20]
  reg [63:0] reg_ex2mem_we_data; // @[Reg.scala 27:20]
  reg [7:0] reg_ex2mem_we_mask; // @[Reg.scala 27:20]
  reg [63:0] reg_ex2wb_result_data; // @[Reg.scala 27:20]
  assign io_prev_ready = io_next_ready; // @[MEMU.scala 17:11]
  assign io_next_valid = io_next_valid_r; // @[MEMU.scala 19:11]
  assign io_next_bits_id2mem_fencei = reg_id2mem_fencei; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_size_byte = reg_id2mem_size_byte; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_size_hword = reg_id2mem_size_hword; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_size_word = reg_id2mem_size_word; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_size_dword = reg_id2mem_size_dword; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_sext_flag = reg_id2mem_sext_flag; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_memory_rd_en = reg_id2mem_memory_rd_en; // @[MEMU.scala 23:12]
  assign io_next_bits_id2mem_memory_we_en = reg_id2mem_memory_we_en; // @[MEMU.scala 23:12]
  assign io_next_bits_id2wb_intr_exce_ret = reg_id2wb_intr_exce_ret; // @[MEMU.scala 23:12]
  assign io_next_bits_id2wb_fencei = reg_id2wb_fencei; // @[MEMU.scala 23:12]
  assign io_next_bits_id2wb_wb_sel = reg_id2wb_wb_sel; // @[MEMU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_en = reg_id2wb_regfile_we_en; // @[MEMU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_addr = reg_id2wb_regfile_we_addr; // @[MEMU.scala 23:12]
  assign io_next_bits_ex2mem_addr = reg_ex2mem_addr; // @[MEMU.scala 23:12]
  assign io_next_bits_ex2mem_we_data = reg_ex2mem_we_data; // @[MEMU.scala 23:12]
  assign io_next_bits_ex2mem_we_mask = reg_ex2mem_we_mask; // @[MEMU.scala 23:12]
  assign io_next_bits_ex2wb_result_data = reg_ex2wb_result_data; // @[MEMU.scala 23:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      io_next_valid_r <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      io_next_valid_r <= io_prev_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_fencei <= data_id2mem_fencei; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_byte <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_byte <= data_id2mem_size_byte; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_hword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_hword <= data_id2mem_size_hword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_word <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_word <= data_id2mem_size_word; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_size_dword <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_size_dword <= data_id2mem_size_dword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_sext_flag <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_sext_flag <= data_id2mem_sext_flag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_memory_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_memory_rd_en <= data_id2mem_memory_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2mem_memory_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2mem_memory_we_en <= data_id2mem_memory_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_intr_exce_ret <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_intr_exce_ret <= data_id2wb_intr_exce_ret; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_fencei <= data_id2wb_fencei; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_wb_sel <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_wb_sel <= data_id2wb_wb_sel; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      reg_id2wb_regfile_we_en <= data_id2wb_regfile_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[MEMU.scala 21:17]
        reg_id2wb_regfile_we_addr <= io_prev_bits_id2wb_regfile_we_addr;
      end else begin
        reg_id2wb_regfile_we_addr <= 5'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_ex2mem_addr <= 39'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[MEMU.scala 21:17]
        reg_ex2mem_addr <= io_prev_bits_ex2mem_addr;
      end else begin
        reg_ex2mem_addr <= 39'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_ex2mem_we_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[MEMU.scala 21:17]
        reg_ex2mem_we_data <= io_prev_bits_ex2mem_we_data;
      end else begin
        reg_ex2mem_we_data <= 64'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_ex2mem_we_mask <= 8'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[MEMU.scala 21:17]
        reg_ex2mem_we_mask <= io_prev_bits_ex2mem_we_mask;
      end else begin
        reg_ex2mem_we_mask <= 8'h0;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_ex2wb_result_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_next_ready) begin // @[Reg.scala 28:19]
      if (io_prev_valid) begin // @[MEMU.scala 21:17]
        reg_ex2wb_result_data <= io_prev_bits_ex2wb_result_data;
      end else begin
        reg_ex2wb_result_data <= 64'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_next_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_id2mem_fencei = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_id2mem_size_byte = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_id2mem_size_hword = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_id2mem_size_word = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_id2mem_size_dword = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  reg_id2mem_sext_flag = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  reg_id2mem_memory_rd_en = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_id2mem_memory_we_en = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  reg_id2wb_intr_exce_ret = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_id2wb_fencei = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_id2wb_wb_sel = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reg_id2wb_regfile_we_en = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  reg_id2wb_regfile_we_addr = _RAND_13[4:0];
  _RAND_14 = {2{`RANDOM}};
  reg_ex2mem_addr = _RAND_14[38:0];
  _RAND_15 = {2{`RANDOM}};
  reg_ex2mem_we_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  reg_ex2mem_we_mask = _RAND_16[7:0];
  _RAND_17 = {2{`RANDOM}};
  reg_ex2wb_result_data = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_DAXIManager(
  input          clock,
  input          reset,
  input          io_in_rd_en,
  input          io_in_we_en,
  input  [31:0]  io_in_addr,
  input  [127:0] io_in_data,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  input          io_maxi_aw_ready,
  output         io_maxi_aw_valid,
  output [31:0]  io_maxi_aw_bits_addr,
  output [7:0]   io_maxi_aw_bits_len,
  output [2:0]   io_maxi_aw_bits_size,
  input          io_maxi_w_ready,
  output         io_maxi_w_valid,
  output [63:0]  io_maxi_w_bits_data,
  output [7:0]   io_maxi_w_bits_strb,
  output         io_maxi_w_bits_last,
  input          io_maxi_b_valid,
  output         io_out_finish,
  output         io_out_ready,
  output [127:0] io_out_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [127:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] curr_state; // @[AXI4Manager.scala 179:35]
  reg  stage_out2_rd_en; // @[Reg.scala 27:20]
  reg  stage_out2_we_en; // @[Reg.scala 27:20]
  reg [31:0] stage_out2_addr; // @[Reg.scala 27:20]
  reg [127:0] stage_out2_data; // @[Reg.scala 27:20]
  reg [15:0] stage_out2_wmask; // @[Reg.scala 27:20]
  wire  stage_en = curr_state == 3'h0; // @[AXI4Manager.scala 204:26]
  wire [15:0] _GEN_0 = stage_en ? 16'hffff : stage_out2_wmask; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [127:0] _GEN_1 = stage_en ? io_in_data : stage_out2_data; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [31:0] _GEN_2 = stage_en ? io_in_addr : stage_out2_addr; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_8 = stage_en ? io_in_we_en : stage_out2_we_en; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_9 = stage_en ? io_in_rd_en : stage_out2_rd_en; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  r_last = io_maxi_r_bits_last & io_maxi_r_valid; // @[AXI4Manager.scala 199:42]
  wire [27:0] a_addr_hi = _GEN_2[31:4]; // @[AXI4Manager.scala 210:39]
  wire [31:0] a_addr = {a_addr_hi,4'h0}; // @[Cat.scala 30:58]
  wire  rdata64_x8 = io_maxi_r_valid & ~io_maxi_r_bits_last; // @[AXI4Manager.scala 213:101]
  reg [63:0] memory_data_lo; // @[Reg.scala 27:20]
  wire [127:0] memory_data = {io_maxi_r_bits_data,memory_data_lo}; // @[Cat.scala 30:58]
  wire  _T = 3'h0 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_11 = io_maxi_ar_ready ? 3'h2 : 3'h1; // @[AXI4Manager.scala 222:29 AXI4Manager.scala 222:42 AXI4Manager.scala 222:79]
  wire [2:0] _GEN_12 = io_maxi_aw_ready ? 3'h5 : 3'h4; // @[AXI4Manager.scala 224:29 AXI4Manager.scala 224:42 AXI4Manager.scala 224:79]
  wire [2:0] _GEN_13 = _GEN_8 ? _GEN_12 : 3'h0; // @[AXI4Manager.scala 223:26 AXI4Manager.scala 225:42]
  wire [2:0] _GEN_14 = _GEN_9 ? _GEN_11 : _GEN_13; // @[AXI4Manager.scala 221:20]
  wire  _T_1 = 3'h1 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h4 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h2 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_15 = io_maxi_r_valid ? 3'h3 : 3'h2; // @[AXI4Manager.scala 236:29 AXI4Manager.scala 236:42 AXI4Manager.scala 237:42]
  wire  _T_4 = 3'h3 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_16 = r_last ? 3'h0 : 3'h3; // @[AXI4Manager.scala 240:29 AXI4Manager.scala 240:42 AXI4Manager.scala 241:42]
  wire  _T_5 = 3'h5 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_17 = io_maxi_w_ready ? 3'h6 : 3'h5; // @[AXI4Manager.scala 244:29 AXI4Manager.scala 244:42 AXI4Manager.scala 245:42]
  wire  _T_6 = 3'h6 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_18 = io_maxi_w_ready ? 3'h7 : 3'h6; // @[AXI4Manager.scala 248:29 AXI4Manager.scala 248:42 AXI4Manager.scala 249:42]
  wire  _T_7 = 3'h7 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_19 = io_maxi_b_valid ? 3'h0 : 3'h7; // @[AXI4Manager.scala 252:29 AXI4Manager.scala 252:42 AXI4Manager.scala 253:42]
  wire [2:0] _GEN_20 = _T_7 ? _GEN_19 : 3'h0; // @[Conditional.scala 39:67 AXI4Manager.scala 218:14]
  wire [2:0] _GEN_21 = _T_6 ? _GEN_18 : _GEN_20; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_22 = _T_5 ? _GEN_17 : _GEN_21; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_23 = _T_4 ? _GEN_16 : _GEN_22; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_24 = _T_3 ? _GEN_15 : _GEN_23; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_25 = _T_2 ? _GEN_12 : _GEN_24; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_26 = _T_1 ? _GEN_11 : _GEN_25; // @[Conditional.scala 39:67]
  wire [2:0] next_state = _T ? _GEN_14 : _GEN_26; // @[Conditional.scala 40:58]
  wire  _T_14 = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1; // @[AXI4Manager.scala 260:80]
  wire [1:0] _GEN_31 = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1 ? 2'h3 : 2'h0; // @[AXI4Manager.scala 260:105 AXI.scala 318:19 AXI.scala 310:19]
  wire  _T_21 = next_state == 3'h4 | stage_en & next_state == 3'h5 | curr_state == 3'h4; // @[AXI4Manager.scala 264:81]
  wire [1:0] _GEN_36 = next_state == 3'h4 | stage_en & next_state == 3'h5 | curr_state == 3'h4 ? 2'h3 : 2'h0; // @[AXI4Manager.scala 264:106 AXI.scala 318:19 AXI.scala 310:19]
  wire  _T_22 = curr_state == 3'h5; // @[AXI4Manager.scala 268:19]
  wire [63:0] _GEN_39 = curr_state == 3'h5 ? _GEN_1[63:0] : 64'h0; // @[AXI4Manager.scala 268:31 AXI.scala 358:19 AXI.scala 364:19]
  wire [7:0] _GEN_40 = curr_state == 3'h5 ? _GEN_0[7:0] : 8'h0; // @[AXI4Manager.scala 268:31 AXI.scala 359:19 AXI.scala 365:19]
  reg [127:0] memory_data_buffer; // @[AXI4Manager.scala 280:43]
  assign io_maxi_ar_valid = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1; // @[AXI4Manager.scala 260:80]
  assign io_maxi_ar_bits_addr = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1 ? a_addr : 32'h0
    ; // @[AXI4Manager.scala 260:105 AXI.scala 317:19 AXI.scala 309:19]
  assign io_maxi_ar_bits_len = {{7'd0}, _T_14}; // @[AXI4Manager.scala 260:80]
  assign io_maxi_ar_bits_size = {{1'd0}, _GEN_31}; // @[AXI4Manager.scala 260:105 AXI.scala 318:19 AXI.scala 310:19]
  assign io_maxi_aw_valid = next_state == 3'h4 | stage_en & next_state == 3'h5 | curr_state == 3'h4; // @[AXI4Manager.scala 264:81]
  assign io_maxi_aw_bits_addr = next_state == 3'h4 | stage_en & next_state == 3'h5 | curr_state == 3'h4 ? a_addr : 32'h0
    ; // @[AXI4Manager.scala 264:106 AXI.scala 317:19 AXI.scala 309:19]
  assign io_maxi_aw_bits_len = {{7'd0}, _T_21}; // @[AXI4Manager.scala 264:81]
  assign io_maxi_aw_bits_size = {{1'd0}, _GEN_36}; // @[AXI4Manager.scala 264:106 AXI.scala 318:19 AXI.scala 310:19]
  assign io_maxi_w_valid = curr_state == 3'h6 | _T_22; // @[AXI4Manager.scala 271:31 AXI.scala 357:15]
  assign io_maxi_w_bits_data = curr_state == 3'h6 ? _GEN_1[127:64] : _GEN_39; // @[AXI4Manager.scala 271:31 AXI.scala 358:19]
  assign io_maxi_w_bits_strb = curr_state == 3'h6 ? _GEN_0[15:8] : _GEN_40; // @[AXI4Manager.scala 271:31 AXI.scala 359:19]
  assign io_maxi_w_bits_last = curr_state == 3'h6; // @[AXI4Manager.scala 271:19]
  assign io_out_finish = io_maxi_r_bits_last | io_maxi_b_valid; // @[AXI4Manager.scala 279:34]
  assign io_out_ready = next_state == 3'h0 | stage_en; // @[AXI4Manager.scala 278:38]
  assign io_out_data = curr_state == 3'h2 | curr_state == 3'h3 ? memory_data : memory_data_buffer; // @[AXI4Manager.scala 282:18]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4Manager.scala 179:35]
      curr_state <= 3'h0; // @[AXI4Manager.scala 179:35]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_GEN_9) begin // @[AXI4Manager.scala 221:20]
        curr_state <= _GEN_11;
      end else if (_GEN_8) begin // @[AXI4Manager.scala 223:26]
        curr_state <= _GEN_12;
      end else begin
        curr_state <= 3'h0; // @[AXI4Manager.scala 225:42]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_11;
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_12;
    end else begin
      curr_state <= _GEN_24;
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_we_en <= io_in_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_addr <= io_in_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_data <= 128'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_data <= io_in_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_wmask <= 16'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_wmask <= 16'hffff; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      memory_data_lo <= 64'h0; // @[Reg.scala 27:20]
    end else if (rdata64_x8) begin // @[Reg.scala 28:19]
      memory_data_lo <= io_maxi_r_bits_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[AXI4Manager.scala 280:43]
      memory_data_buffer <= 128'h0; // @[AXI4Manager.scala 280:43]
    end else if (io_out_finish) begin // @[AXI4Manager.scala 281:28]
      memory_data_buffer <= memory_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  stage_out2_rd_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stage_out2_we_en = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  stage_out2_addr = _RAND_3[31:0];
  _RAND_4 = {4{`RANDOM}};
  stage_out2_data = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  stage_out2_wmask = _RAND_5[15:0];
  _RAND_6 = {2{`RANDOM}};
  memory_data_lo = _RAND_6[63:0];
  _RAND_7 = {4{`RANDOM}};
  memory_data_buffer = _RAND_7[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_AXI4LiteManager(
  input         clock,
  input         reset,
  input         io_in_rd_en,
  input         io_in_we_en,
  input         io_in_size_byte,
  input         io_in_size_hword,
  input         io_in_size_word,
  input         io_in_size_dword,
  input  [31:0] io_in_addr,
  input  [63:0] io_in_data,
  input  [15:0] io_in_wmask,
  input         io_maxi_ar_ready,
  output        io_maxi_ar_valid,
  output [31:0] io_maxi_ar_bits_addr,
  output [2:0]  io_maxi_ar_bits_size,
  input         io_maxi_r_valid,
  input  [63:0] io_maxi_r_bits_data,
  input         io_maxi_r_bits_last,
  input         io_maxi_aw_ready,
  output        io_maxi_aw_valid,
  output [31:0] io_maxi_aw_bits_addr,
  output [2:0]  io_maxi_aw_bits_size,
  input         io_maxi_w_ready,
  output        io_maxi_w_valid,
  output [63:0] io_maxi_w_bits_data,
  output [7:0]  io_maxi_w_bits_strb,
  output        io_maxi_w_bits_last,
  input         io_maxi_b_valid,
  output        io_out_finish,
  output        io_out_ready,
  output [63:0] io_out_data,
  output        clint_we_0,
  output [31:0] _T_24_0,
  input  [63:0] clint_rdata_0,
  output [63:0] clint_wdata_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] curr_state; // @[AXI4LiteManager.scala 47:35]
  reg  stage_out2_rd_en; // @[Reg.scala 27:20]
  reg  stage_out2_we_en; // @[Reg.scala 27:20]
  reg  stage_out2_size_byte; // @[Reg.scala 27:20]
  reg  stage_out2_size_hword; // @[Reg.scala 27:20]
  reg  stage_out2_size_word; // @[Reg.scala 27:20]
  reg  stage_out2_size_dword; // @[Reg.scala 27:20]
  reg [31:0] stage_out2_addr; // @[Reg.scala 27:20]
  reg [63:0] stage_out2_data; // @[Reg.scala 27:20]
  reg [15:0] stage_out2_wmask; // @[Reg.scala 27:20]
  wire  stage_en = curr_state == 3'h0; // @[AXI4LiteManager.scala 73:26]
  wire [15:0] _GEN_0 = stage_en ? io_in_wmask : stage_out2_wmask; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [63:0] _GEN_1 = stage_en ? io_in_data : stage_out2_data; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [31:0] _GEN_2 = stage_en ? io_in_addr : stage_out2_addr; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_3 = stage_en ? io_in_size_dword : stage_out2_size_dword; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_4 = stage_en ? io_in_size_word : stage_out2_size_word; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_5 = stage_en ? io_in_size_hword : stage_out2_size_hword; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_6 = stage_en ? io_in_size_byte : stage_out2_size_byte; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_7 = stage_en ? io_in_we_en : stage_out2_we_en; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_8 = stage_en ? io_in_rd_en : stage_out2_rd_en; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  in2__size_byte = stage_en ? io_in_size_byte : stage_out2_size_byte; // @[AXI4LiteManager.scala 55:24]
  wire  in2__size_hword = stage_en ? io_in_size_hword : stage_out2_size_hword; // @[AXI4LiteManager.scala 55:24]
  wire  in2__size_word = stage_en ? io_in_size_word : stage_out2_size_word; // @[AXI4LiteManager.scala 55:24]
  wire  in2__size_dword = stage_en ? io_in_size_dword : stage_out2_size_dword; // @[AXI4LiteManager.scala 55:24]
  wire  is_uart = _GEN_2 > 32'hfffffff & _GEN_2 < 32'h10000fff; // @[AXI4LiteManager.scala 56:51]
  wire  r_last = io_maxi_r_bits_last & io_maxi_r_valid; // @[AXI4LiteManager.scala 66:42]
  wire  is_clint = _GEN_2[31:16] == 16'h200 & _GEN_2[16:15] != 2'h3; // @[AXI4LiteManager.scala 68:59]
  wire [29:0] a_addr_hi = _GEN_2[31:2]; // @[AXI4LiteManager.scala 77:69]
  wire [31:0] _a_addr_T_1 = {a_addr_hi,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] a_addr = is_uart ? _GEN_2 : _a_addr_T_1; // @[AXI4LiteManager.scala 77:30]
  wire [1:0] _a_size_T = _GEN_3 ? 2'h3 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _a_size_T_1 = _GEN_4 ? 2'h2 : _a_size_T; // @[Mux.scala 98:16]
  wire [1:0] _a_size_T_2 = _GEN_5 ? 2'h1 : _a_size_T_1; // @[Mux.scala 98:16]
  wire [1:0] a_size = _GEN_6 ? 2'h0 : _a_size_T_2; // @[Mux.scala 98:16]
  wire [2:0] start_byte = _GEN_2[2:0]; // @[AXI4LiteManager.scala 84:36]
  wire [5:0] start_bit = {start_byte, 3'h0}; // @[AXI4LiteManager.scala 85:45]
  wire [63:0] rdata_out_1 = io_maxi_r_bits_data >> start_bit; // @[AXI4LiteManager.scala 87:46]
  wire  _rdata_out_T = curr_state == 3'h6; // @[AXI4LiteManager.scala 90:17]
  wire  _rdata_out_T_1 = curr_state == 3'h2; // @[AXI4LiteManager.scala 91:17]
  wire [63:0] _rdata_out_T_2 = _rdata_out_T_1 ? rdata_out_1 : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] rdata_out = _rdata_out_T ? clint_rdata_0 : _rdata_out_T_2; // @[Mux.scala 98:16]
  wire [63:0] _memory_data_T_4 = _GEN_3 ? rdata_out : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _memory_data_T_5 = _GEN_4 ? {{32'd0}, rdata_out[31:0]} : _memory_data_T_4; // @[Mux.scala 98:16]
  wire [63:0] _memory_data_T_6 = _GEN_5 ? {{48'd0}, rdata_out[15:0]} : _memory_data_T_5; // @[Mux.scala 98:16]
  wire [63:0] memory_data = _GEN_6 ? {{56'd0}, rdata_out[7:0]} : _memory_data_T_6; // @[Mux.scala 98:16]
  wire [126:0] _GEN_41 = {{63'd0}, _GEN_1}; // @[AXI4LiteManager.scala 102:33]
  wire [126:0] _wdata_T = _GEN_41 << start_bit; // @[AXI4LiteManager.scala 102:33]
  wire [22:0] _GEN_42 = {{7'd0}, _GEN_0}; // @[AXI4LiteManager.scala 104:31]
  wire [22:0] _wmask_T = _GEN_42 << start_byte; // @[AXI4LiteManager.scala 104:31]
  wire [22:0] _wmask_T_4 = _GEN_3 ? _wmask_T : 23'h0; // @[Mux.scala 98:16]
  wire [22:0] _wmask_T_5 = _GEN_4 ? _wmask_T : _wmask_T_4; // @[Mux.scala 98:16]
  wire [22:0] _wmask_T_6 = _GEN_5 ? _wmask_T : _wmask_T_5; // @[Mux.scala 98:16]
  wire [22:0] wmask = _GEN_6 ? _wmask_T : _wmask_T_6; // @[Mux.scala 98:16]
  wire  _T = 3'h0 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_9 = io_maxi_ar_ready ? 3'h2 : 3'h1; // @[AXI4LiteManager.scala 118:37 AXI4LiteManager.scala 118:50 AXI4LiteManager.scala 119:50]
  wire [2:0] _GEN_10 = is_clint ? 3'h6 : _GEN_9; // @[AXI4LiteManager.scala 117:37 AXI4LiteManager.scala 117:50]
  wire [2:0] _GEN_11 = io_maxi_aw_ready ? 3'h4 : 3'h3; // @[AXI4LiteManager.scala 122:37 AXI4LiteManager.scala 122:50 AXI4LiteManager.scala 123:50]
  wire [2:0] _GEN_12 = is_clint ? 3'h7 : _GEN_11; // @[AXI4LiteManager.scala 121:37 AXI4LiteManager.scala 121:50]
  wire [2:0] _GEN_13 = _GEN_7 ? _GEN_12 : 3'h0; // @[AXI4LiteManager.scala 120:26 AXI4LiteManager.scala 124:50]
  wire [2:0] _GEN_14 = _GEN_8 ? _GEN_10 : _GEN_13; // @[AXI4LiteManager.scala 116:20]
  wire  _T_1 = 3'h1 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h3 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_3 = 3'h2 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_15 = r_last ? 3'h0 : 3'h2; // @[AXI4LiteManager.scala 135:29 AXI4LiteManager.scala 135:42 AXI4LiteManager.scala 136:42]
  wire  _T_4 = 3'h4 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_16 = io_maxi_w_ready ? 3'h5 : 3'h4; // @[AXI4LiteManager.scala 139:29 AXI4LiteManager.scala 139:42 AXI4LiteManager.scala 140:42]
  wire  _T_5 = 3'h5 == curr_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_17 = io_maxi_b_valid ? 3'h0 : 3'h5; // @[AXI4LiteManager.scala 143:29 AXI4LiteManager.scala 143:42 AXI4LiteManager.scala 144:42]
  wire [2:0] _GEN_20 = _T_5 ? _GEN_17 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_21 = _T_4 ? _GEN_16 : _GEN_20; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_22 = _T_3 ? _GEN_15 : _GEN_21; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_23 = _T_2 ? _GEN_11 : _GEN_22; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_24 = _T_1 ? _GEN_9 : _GEN_23; // @[Conditional.scala 39:67]
  wire [2:0] next_state = _T ? _GEN_14 : _GEN_24; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_29 = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1 ? a_size : 2'h0; // @[AXI4LiteManager.scala 151:104 AXI.scala 318:19 AXI.scala 310:19]
  wire [1:0] _GEN_35 = next_state == 3'h3 | stage_en & next_state == 3'h4 | curr_state == 3'h3 ? a_size : 2'h0; // @[AXI4LiteManager.scala 155:106 AXI.scala 318:19 AXI.scala 310:19]
  wire [127:0] wdata = {{1'd0}, _wdata_T}; // @[AXI4LiteManager.scala 102:55 AXI4LiteManager.scala 102:55]
  wire [22:0] _GEN_40 = curr_state == 3'h4 ? wmask : 23'h0; // @[AXI4LiteManager.scala 159:31 AXI.scala 359:19 AXI.scala 365:19]
  wire [31:0] _clint_addr_T = a_addr; // @[AXI4LiteManager.scala 77:30]
  wire [31:0] _T_24 = a_addr; // @[AXI4LiteManager.scala 77:30]
  reg [63:0] memory_data_buffer; // @[AXI4LiteManager.scala 179:43]
  wire [63:0] clint_wdata = wdata[63:0]; // @[AXI4LiteManager.scala 170:23]
  wire  clint_we = next_state == 3'h7; // @[AXI4LiteManager.scala 168:29]
  assign io_maxi_ar_valid = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1; // @[AXI4LiteManager.scala 151:79]
  assign io_maxi_ar_bits_addr = next_state == 3'h1 | stage_en & next_state == 3'h2 | curr_state == 3'h1 ? a_addr : 32'h0
    ; // @[AXI4LiteManager.scala 151:104 AXI.scala 317:19 AXI.scala 309:19]
  assign io_maxi_ar_bits_size = {{1'd0}, _GEN_29}; // @[AXI4LiteManager.scala 151:104 AXI.scala 318:19 AXI.scala 310:19]
  assign io_maxi_aw_valid = next_state == 3'h3 | stage_en & next_state == 3'h4 | curr_state == 3'h3; // @[AXI4LiteManager.scala 155:81]
  assign io_maxi_aw_bits_addr = next_state == 3'h3 | stage_en & next_state == 3'h4 | curr_state == 3'h3 ? a_addr : 32'h0
    ; // @[AXI4LiteManager.scala 155:106 AXI.scala 317:19 AXI.scala 309:19]
  assign io_maxi_aw_bits_size = {{1'd0}, _GEN_35}; // @[AXI4LiteManager.scala 155:106 AXI.scala 318:19 AXI.scala 310:19]
  assign io_maxi_w_valid = curr_state == 3'h4; // @[AXI4LiteManager.scala 159:19]
  assign io_maxi_w_bits_data = curr_state == 3'h4 ? wdata[63:0] : 64'h0; // @[AXI4LiteManager.scala 159:31 AXI.scala 358:19 AXI.scala 364:19]
  assign io_maxi_w_bits_strb = _GEN_40[7:0];
  assign io_maxi_w_bits_last = curr_state == 3'h4; // @[AXI4LiteManager.scala 159:19]
  assign io_out_finish = io_maxi_r_bits_last | io_maxi_b_valid | curr_state == 3'h7 | _rdata_out_T; // @[AXI4LiteManager.scala 178:74]
  assign io_out_ready = next_state == 3'h0 | stage_en; // @[AXI4LiteManager.scala 177:38]
  assign io_out_data = _rdata_out_T_1 | _rdata_out_T ? memory_data : memory_data_buffer; // @[AXI4LiteManager.scala 181:18]
  assign clint_we_0 = clint_we;
  assign _T_24_0 = _clint_addr_T;
  assign clint_wdata_0 = clint_wdata;
  always @(posedge clock) begin
    if (reset) begin // @[AXI4LiteManager.scala 47:35]
      curr_state <= 3'h0; // @[AXI4LiteManager.scala 47:35]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_GEN_8) begin // @[AXI4LiteManager.scala 116:20]
        if (is_clint) begin // @[AXI4LiteManager.scala 117:37]
          curr_state <= 3'h6; // @[AXI4LiteManager.scala 117:50]
        end else begin
          curr_state <= _GEN_9;
        end
      end else if (_GEN_7) begin // @[AXI4LiteManager.scala 120:26]
        curr_state <= _GEN_12;
      end else begin
        curr_state <= 3'h0; // @[AXI4LiteManager.scala 124:50]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_9;
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_11;
    end else begin
      curr_state <= _GEN_22;
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_rd_en <= io_in_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_we_en <= io_in_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_size_byte <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_size_byte <= io_in_size_byte; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_size_hword <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_size_hword <= io_in_size_hword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_size_word <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_size_word <= io_in_size_word; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_size_dword <= 1'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_size_dword <= io_in_size_dword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_addr <= io_in_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_data <= io_in_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage_out2_wmask <= 16'h0; // @[Reg.scala 27:20]
    end else if (stage_en) begin // @[Reg.scala 28:19]
      stage_out2_wmask <= io_in_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[AXI4LiteManager.scala 179:43]
      memory_data_buffer <= 64'h0; // @[AXI4LiteManager.scala 179:43]
    end else if (io_out_finish) begin // @[AXI4LiteManager.scala 180:28]
      if (_GEN_6) begin // @[Mux.scala 98:16]
        memory_data_buffer <= {{56'd0}, rdata_out[7:0]};
      end else if (_GEN_5) begin // @[Mux.scala 98:16]
        memory_data_buffer <= {{48'd0}, rdata_out[15:0]};
      end else begin
        memory_data_buffer <= _memory_data_T_5;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  stage_out2_rd_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stage_out2_we_en = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  stage_out2_size_byte = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  stage_out2_size_hword = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  stage_out2_size_word = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stage_out2_size_dword = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  stage_out2_addr = _RAND_7[31:0];
  _RAND_8 = {2{`RANDOM}};
  stage_out2_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  stage_out2_wmask = _RAND_9[15:0];
  _RAND_10 = {2{`RANDOM}};
  memory_data_buffer = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_DCacheUnit(
  input          clock,
  input          reset,
  output         io_next_valid,
  output         io_next_bits_data_id2wb_intr_exce_ret,
  output         io_next_bits_data_id2wb_fencei,
  output         io_next_bits_data_id2wb_wb_sel,
  output         io_next_bits_data_id2wb_regfile_we_en,
  output [4:0]   io_next_bits_data_id2wb_regfile_we_addr,
  output [63:0]  io_next_bits_data_ex2wb_result_data,
  output [63:0]  io_next_bits_data_mem2wb_memory_data,
  output         io_prev_ready,
  input          io_prev_valid,
  input          io_prev_bits_data_id2mem_sext_flag,
  input          io_prev_bits_data_id2mem_memory_rd_en,
  input          io_prev_bits_data_id2mem_memory_we_en,
  input          io_prev_bits_data_id2wb_intr_exce_ret,
  input          io_prev_bits_data_id2wb_fencei,
  input          io_prev_bits_data_id2wb_wb_sel,
  input          io_prev_bits_data_id2wb_regfile_we_en,
  input  [4:0]   io_prev_bits_data_id2wb_regfile_we_addr,
  input  [63:0]  io_prev_bits_data_ex2mem_we_data,
  input  [63:0]  io_prev_bits_data_ex2wb_result_data,
  input          io_prev_bits_flush,
  input  [63:0]  io_prev_bits_wdata,
  input  [7:0]   io_prev_bits_wmask,
  input          io_prev_bits_size_byte,
  input          io_prev_bits_size_hword,
  input          io_prev_bits_size_word,
  input          io_prev_bits_size_dword,
  input  [38:0]  io_prev_bits_addr,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  input          io_maxi_aw_ready,
  output         io_maxi_aw_valid,
  output [31:0]  io_maxi_aw_bits_addr,
  output [7:0]   io_maxi_aw_bits_len,
  output [2:0]   io_maxi_aw_bits_size,
  input          io_maxi_w_ready,
  output         io_maxi_w_valid,
  output [63:0]  io_maxi_w_bits_data,
  output [7:0]   io_maxi_w_bits_strb,
  output         io_maxi_w_bits_last,
  input          io_maxi_b_valid,
  input          io_mmio_ar_ready,
  output         io_mmio_ar_valid,
  output [31:0]  io_mmio_ar_bits_addr,
  output [2:0]   io_mmio_ar_bits_size,
  input          io_mmio_r_valid,
  input  [63:0]  io_mmio_r_bits_data,
  input          io_mmio_r_bits_last,
  input          io_mmio_aw_ready,
  output         io_mmio_aw_valid,
  output [31:0]  io_mmio_aw_bits_addr,
  output [2:0]   io_mmio_aw_bits_size,
  input          io_mmio_w_ready,
  output         io_mmio_w_valid,
  output [63:0]  io_mmio_w_bits_data,
  output [7:0]   io_mmio_w_bits_strb,
  output         io_mmio_w_bits_last,
  input          io_mmio_b_valid,
  output [5:0]   io_sram4_addr,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,
  output         clint_we,
  output [31:0]  _T_24_0,
  input  [63:0]  clint_rdata,
  output [63:0]  clint_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [63:0] _RAND_335;
  reg [63:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
`endif // RANDOMIZE_REG_INIT
  wire  maxi4_manager_clock; // @[DCache.scala 70:29]
  wire  maxi4_manager_reset; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_in_rd_en; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_in_we_en; // @[DCache.scala 70:29]
  wire [31:0] maxi4_manager_io_in_addr; // @[DCache.scala 70:29]
  wire [127:0] maxi4_manager_io_in_data; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_ar_ready; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_ar_valid; // @[DCache.scala 70:29]
  wire [31:0] maxi4_manager_io_maxi_ar_bits_addr; // @[DCache.scala 70:29]
  wire [7:0] maxi4_manager_io_maxi_ar_bits_len; // @[DCache.scala 70:29]
  wire [2:0] maxi4_manager_io_maxi_ar_bits_size; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_r_valid; // @[DCache.scala 70:29]
  wire [63:0] maxi4_manager_io_maxi_r_bits_data; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_r_bits_last; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_aw_ready; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_aw_valid; // @[DCache.scala 70:29]
  wire [31:0] maxi4_manager_io_maxi_aw_bits_addr; // @[DCache.scala 70:29]
  wire [7:0] maxi4_manager_io_maxi_aw_bits_len; // @[DCache.scala 70:29]
  wire [2:0] maxi4_manager_io_maxi_aw_bits_size; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_w_ready; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_w_valid; // @[DCache.scala 70:29]
  wire [63:0] maxi4_manager_io_maxi_w_bits_data; // @[DCache.scala 70:29]
  wire [7:0] maxi4_manager_io_maxi_w_bits_strb; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_w_bits_last; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_maxi_b_valid; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_out_finish; // @[DCache.scala 70:29]
  wire  maxi4_manager_io_out_ready; // @[DCache.scala 70:29]
  wire [127:0] maxi4_manager_io_out_data; // @[DCache.scala 70:29]
  wire  mmio_manager_clock; // @[DCache.scala 83:28]
  wire  mmio_manager_reset; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_rd_en; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_we_en; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_size_byte; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_size_hword; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_size_word; // @[DCache.scala 83:28]
  wire  mmio_manager_io_in_size_dword; // @[DCache.scala 83:28]
  wire [31:0] mmio_manager_io_in_addr; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_io_in_data; // @[DCache.scala 83:28]
  wire [15:0] mmio_manager_io_in_wmask; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_ar_ready; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_ar_valid; // @[DCache.scala 83:28]
  wire [31:0] mmio_manager_io_maxi_ar_bits_addr; // @[DCache.scala 83:28]
  wire [2:0] mmio_manager_io_maxi_ar_bits_size; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_r_valid; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_io_maxi_r_bits_data; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_r_bits_last; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_aw_ready; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_aw_valid; // @[DCache.scala 83:28]
  wire [31:0] mmio_manager_io_maxi_aw_bits_addr; // @[DCache.scala 83:28]
  wire [2:0] mmio_manager_io_maxi_aw_bits_size; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_w_ready; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_w_valid; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_io_maxi_w_bits_data; // @[DCache.scala 83:28]
  wire [7:0] mmio_manager_io_maxi_w_bits_strb; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_w_bits_last; // @[DCache.scala 83:28]
  wire  mmio_manager_io_maxi_b_valid; // @[DCache.scala 83:28]
  wire  mmio_manager_io_out_finish; // @[DCache.scala 83:28]
  wire  mmio_manager_io_out_ready; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_io_out_data; // @[DCache.scala 83:28]
  wire  mmio_manager_clint_we_0; // @[DCache.scala 83:28]
  wire [31:0] mmio_manager__T_24_0; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_clint_rdata_0; // @[DCache.scala 83:28]
  wire [63:0] mmio_manager_clint_wdata_0; // @[DCache.scala 83:28]
  reg [3:0] curr_state; // @[DCache.scala 65:37]
  wire  _T_16 = curr_state == 4'h2; // @[DCache.scala 269:19]
  reg [38:0] stage1_out_bits_addr; // @[Reg.scala 27:20]
  wire [5:0] stage1_index = stage1_out_bits_addr[9:4]; // @[DCache.scala 160:54]
  reg  lru_list_63; // @[DCache.scala 118:35]
  reg  lru_list_62; // @[DCache.scala 118:35]
  reg  lru_list_61; // @[DCache.scala 118:35]
  reg  lru_list_60; // @[DCache.scala 118:35]
  reg  lru_list_59; // @[DCache.scala 118:35]
  reg  lru_list_58; // @[DCache.scala 118:35]
  reg  lru_list_57; // @[DCache.scala 118:35]
  reg  lru_list_56; // @[DCache.scala 118:35]
  reg  lru_list_55; // @[DCache.scala 118:35]
  reg  lru_list_54; // @[DCache.scala 118:35]
  reg  lru_list_53; // @[DCache.scala 118:35]
  reg  lru_list_52; // @[DCache.scala 118:35]
  reg  lru_list_51; // @[DCache.scala 118:35]
  reg  lru_list_50; // @[DCache.scala 118:35]
  reg  lru_list_49; // @[DCache.scala 118:35]
  reg  lru_list_48; // @[DCache.scala 118:35]
  reg  lru_list_47; // @[DCache.scala 118:35]
  reg  lru_list_46; // @[DCache.scala 118:35]
  reg  lru_list_45; // @[DCache.scala 118:35]
  reg  lru_list_44; // @[DCache.scala 118:35]
  reg  lru_list_43; // @[DCache.scala 118:35]
  reg  lru_list_42; // @[DCache.scala 118:35]
  reg  lru_list_41; // @[DCache.scala 118:35]
  reg  lru_list_40; // @[DCache.scala 118:35]
  reg  lru_list_39; // @[DCache.scala 118:35]
  reg  lru_list_38; // @[DCache.scala 118:35]
  reg  lru_list_37; // @[DCache.scala 118:35]
  reg  lru_list_36; // @[DCache.scala 118:35]
  reg  lru_list_35; // @[DCache.scala 118:35]
  reg  lru_list_34; // @[DCache.scala 118:35]
  reg  lru_list_33; // @[DCache.scala 118:35]
  reg  lru_list_32; // @[DCache.scala 118:35]
  reg  lru_list_31; // @[DCache.scala 118:35]
  reg  lru_list_30; // @[DCache.scala 118:35]
  reg  lru_list_29; // @[DCache.scala 118:35]
  reg  lru_list_28; // @[DCache.scala 118:35]
  reg  lru_list_27; // @[DCache.scala 118:35]
  reg  lru_list_26; // @[DCache.scala 118:35]
  reg  lru_list_25; // @[DCache.scala 118:35]
  reg  lru_list_24; // @[DCache.scala 118:35]
  reg  lru_list_23; // @[DCache.scala 118:35]
  reg  lru_list_22; // @[DCache.scala 118:35]
  reg  lru_list_21; // @[DCache.scala 118:35]
  reg  lru_list_20; // @[DCache.scala 118:35]
  reg  lru_list_19; // @[DCache.scala 118:35]
  reg  lru_list_18; // @[DCache.scala 118:35]
  reg  lru_list_17; // @[DCache.scala 118:35]
  reg  lru_list_16; // @[DCache.scala 118:35]
  reg  lru_list_15; // @[DCache.scala 118:35]
  reg  lru_list_14; // @[DCache.scala 118:35]
  reg  lru_list_13; // @[DCache.scala 118:35]
  reg  lru_list_12; // @[DCache.scala 118:35]
  reg  lru_list_11; // @[DCache.scala 118:35]
  reg  lru_list_10; // @[DCache.scala 118:35]
  reg  lru_list_9; // @[DCache.scala 118:35]
  reg  lru_list_8; // @[DCache.scala 118:35]
  reg  lru_list_7; // @[DCache.scala 118:35]
  reg  lru_list_6; // @[DCache.scala 118:35]
  reg  lru_list_5; // @[DCache.scala 118:35]
  reg  lru_list_4; // @[DCache.scala 118:35]
  reg  lru_list_3; // @[DCache.scala 118:35]
  reg  lru_list_2; // @[DCache.scala 118:35]
  reg  lru_list_1; // @[DCache.scala 118:35]
  reg  lru_list_0; // @[DCache.scala 118:35]
  wire  _GEN_166 = 6'h1 == stage1_index ? lru_list_1 : lru_list_0; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_167 = 6'h2 == stage1_index ? lru_list_2 : _GEN_166; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_168 = 6'h3 == stage1_index ? lru_list_3 : _GEN_167; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_169 = 6'h4 == stage1_index ? lru_list_4 : _GEN_168; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_170 = 6'h5 == stage1_index ? lru_list_5 : _GEN_169; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_171 = 6'h6 == stage1_index ? lru_list_6 : _GEN_170; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_172 = 6'h7 == stage1_index ? lru_list_7 : _GEN_171; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_173 = 6'h8 == stage1_index ? lru_list_8 : _GEN_172; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_174 = 6'h9 == stage1_index ? lru_list_9 : _GEN_173; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_175 = 6'ha == stage1_index ? lru_list_10 : _GEN_174; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_176 = 6'hb == stage1_index ? lru_list_11 : _GEN_175; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_177 = 6'hc == stage1_index ? lru_list_12 : _GEN_176; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_178 = 6'hd == stage1_index ? lru_list_13 : _GEN_177; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_179 = 6'he == stage1_index ? lru_list_14 : _GEN_178; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_180 = 6'hf == stage1_index ? lru_list_15 : _GEN_179; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_181 = 6'h10 == stage1_index ? lru_list_16 : _GEN_180; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_182 = 6'h11 == stage1_index ? lru_list_17 : _GEN_181; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_183 = 6'h12 == stage1_index ? lru_list_18 : _GEN_182; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_184 = 6'h13 == stage1_index ? lru_list_19 : _GEN_183; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_185 = 6'h14 == stage1_index ? lru_list_20 : _GEN_184; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_186 = 6'h15 == stage1_index ? lru_list_21 : _GEN_185; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_187 = 6'h16 == stage1_index ? lru_list_22 : _GEN_186; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_188 = 6'h17 == stage1_index ? lru_list_23 : _GEN_187; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_189 = 6'h18 == stage1_index ? lru_list_24 : _GEN_188; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_190 = 6'h19 == stage1_index ? lru_list_25 : _GEN_189; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_191 = 6'h1a == stage1_index ? lru_list_26 : _GEN_190; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_192 = 6'h1b == stage1_index ? lru_list_27 : _GEN_191; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_193 = 6'h1c == stage1_index ? lru_list_28 : _GEN_192; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_194 = 6'h1d == stage1_index ? lru_list_29 : _GEN_193; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_195 = 6'h1e == stage1_index ? lru_list_30 : _GEN_194; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_196 = 6'h1f == stage1_index ? lru_list_31 : _GEN_195; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_197 = 6'h20 == stage1_index ? lru_list_32 : _GEN_196; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_198 = 6'h21 == stage1_index ? lru_list_33 : _GEN_197; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_199 = 6'h22 == stage1_index ? lru_list_34 : _GEN_198; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_200 = 6'h23 == stage1_index ? lru_list_35 : _GEN_199; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_201 = 6'h24 == stage1_index ? lru_list_36 : _GEN_200; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_202 = 6'h25 == stage1_index ? lru_list_37 : _GEN_201; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_203 = 6'h26 == stage1_index ? lru_list_38 : _GEN_202; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_204 = 6'h27 == stage1_index ? lru_list_39 : _GEN_203; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_205 = 6'h28 == stage1_index ? lru_list_40 : _GEN_204; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_206 = 6'h29 == stage1_index ? lru_list_41 : _GEN_205; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_207 = 6'h2a == stage1_index ? lru_list_42 : _GEN_206; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_208 = 6'h2b == stage1_index ? lru_list_43 : _GEN_207; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_209 = 6'h2c == stage1_index ? lru_list_44 : _GEN_208; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_210 = 6'h2d == stage1_index ? lru_list_45 : _GEN_209; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_211 = 6'h2e == stage1_index ? lru_list_46 : _GEN_210; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_212 = 6'h2f == stage1_index ? lru_list_47 : _GEN_211; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_213 = 6'h30 == stage1_index ? lru_list_48 : _GEN_212; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_214 = 6'h31 == stage1_index ? lru_list_49 : _GEN_213; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_215 = 6'h32 == stage1_index ? lru_list_50 : _GEN_214; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_216 = 6'h33 == stage1_index ? lru_list_51 : _GEN_215; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_217 = 6'h34 == stage1_index ? lru_list_52 : _GEN_216; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_218 = 6'h35 == stage1_index ? lru_list_53 : _GEN_217; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_219 = 6'h36 == stage1_index ? lru_list_54 : _GEN_218; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_220 = 6'h37 == stage1_index ? lru_list_55 : _GEN_219; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_221 = 6'h38 == stage1_index ? lru_list_56 : _GEN_220; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_222 = 6'h39 == stage1_index ? lru_list_57 : _GEN_221; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_223 = 6'h3a == stage1_index ? lru_list_58 : _GEN_222; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_224 = 6'h3b == stage1_index ? lru_list_59 : _GEN_223; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_225 = 6'h3c == stage1_index ? lru_list_60 : _GEN_224; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_226 = 6'h3d == stage1_index ? lru_list_61 : _GEN_225; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_227 = 6'h3e == stage1_index ? lru_list_62 : _GEN_226; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  _GEN_228 = 6'h3f == stage1_index ? lru_list_63 : _GEN_227; // @[DCache.scala 172:35 DCache.scala 172:35]
  wire  next_way = ~_GEN_228; // @[DCache.scala 172:35]
  wire  _T_18 = curr_state == 4'hb; // @[DCache.scala 286:26]
  reg [6:0] value; // @[Counter.scala 60:40]
  wire  flush_way = value[6]; // @[DCache.scala 127:45]
  wire  _T_19 = curr_state == 4'h1; // @[DCache.scala 297:26]
  reg  hit_reg; // @[Reg.scala 27:20]
  wire  _T_20 = ~hit_reg; // @[DCache.scala 298:20]
  wire [29:0] tag_array_out_0 = io_sram6_rdata[29:0]; // @[DCache.scala 110:50]
  wire [29:0] tag_array_out_1 = io_sram7_rdata[29:0]; // @[DCache.scala 111:50]
  reg  dirty_array_0_0; // @[DCache.scala 113:44]
  reg  dirty_array_0_1; // @[DCache.scala 113:44]
  reg  dirty_array_0_2; // @[DCache.scala 113:44]
  reg  dirty_array_0_3; // @[DCache.scala 113:44]
  reg  dirty_array_0_4; // @[DCache.scala 113:44]
  reg  dirty_array_0_5; // @[DCache.scala 113:44]
  reg  dirty_array_0_6; // @[DCache.scala 113:44]
  reg  dirty_array_0_7; // @[DCache.scala 113:44]
  reg  dirty_array_0_8; // @[DCache.scala 113:44]
  reg  dirty_array_0_9; // @[DCache.scala 113:44]
  reg  dirty_array_0_10; // @[DCache.scala 113:44]
  reg  dirty_array_0_11; // @[DCache.scala 113:44]
  reg  dirty_array_0_12; // @[DCache.scala 113:44]
  reg  dirty_array_0_13; // @[DCache.scala 113:44]
  reg  dirty_array_0_14; // @[DCache.scala 113:44]
  reg  dirty_array_0_15; // @[DCache.scala 113:44]
  reg  dirty_array_0_16; // @[DCache.scala 113:44]
  reg  dirty_array_0_17; // @[DCache.scala 113:44]
  reg  dirty_array_0_18; // @[DCache.scala 113:44]
  reg  dirty_array_0_19; // @[DCache.scala 113:44]
  reg  dirty_array_0_20; // @[DCache.scala 113:44]
  reg  dirty_array_0_21; // @[DCache.scala 113:44]
  reg  dirty_array_0_22; // @[DCache.scala 113:44]
  reg  dirty_array_0_23; // @[DCache.scala 113:44]
  reg  dirty_array_0_24; // @[DCache.scala 113:44]
  reg  dirty_array_0_25; // @[DCache.scala 113:44]
  reg  dirty_array_0_26; // @[DCache.scala 113:44]
  reg  dirty_array_0_27; // @[DCache.scala 113:44]
  reg  dirty_array_0_28; // @[DCache.scala 113:44]
  reg  dirty_array_0_29; // @[DCache.scala 113:44]
  reg  dirty_array_0_30; // @[DCache.scala 113:44]
  reg  dirty_array_0_31; // @[DCache.scala 113:44]
  reg  dirty_array_0_32; // @[DCache.scala 113:44]
  reg  dirty_array_0_33; // @[DCache.scala 113:44]
  reg  dirty_array_0_34; // @[DCache.scala 113:44]
  reg  dirty_array_0_35; // @[DCache.scala 113:44]
  reg  dirty_array_0_36; // @[DCache.scala 113:44]
  reg  dirty_array_0_37; // @[DCache.scala 113:44]
  reg  dirty_array_0_38; // @[DCache.scala 113:44]
  reg  dirty_array_0_39; // @[DCache.scala 113:44]
  reg  dirty_array_0_40; // @[DCache.scala 113:44]
  reg  dirty_array_0_41; // @[DCache.scala 113:44]
  reg  dirty_array_0_42; // @[DCache.scala 113:44]
  reg  dirty_array_0_43; // @[DCache.scala 113:44]
  reg  dirty_array_0_44; // @[DCache.scala 113:44]
  reg  dirty_array_0_45; // @[DCache.scala 113:44]
  reg  dirty_array_0_46; // @[DCache.scala 113:44]
  reg  dirty_array_0_47; // @[DCache.scala 113:44]
  reg  dirty_array_0_48; // @[DCache.scala 113:44]
  reg  dirty_array_0_49; // @[DCache.scala 113:44]
  reg  dirty_array_0_50; // @[DCache.scala 113:44]
  reg  dirty_array_0_51; // @[DCache.scala 113:44]
  reg  dirty_array_0_52; // @[DCache.scala 113:44]
  reg  dirty_array_0_53; // @[DCache.scala 113:44]
  reg  dirty_array_0_54; // @[DCache.scala 113:44]
  reg  dirty_array_0_55; // @[DCache.scala 113:44]
  reg  dirty_array_0_56; // @[DCache.scala 113:44]
  reg  dirty_array_0_57; // @[DCache.scala 113:44]
  reg  dirty_array_0_58; // @[DCache.scala 113:44]
  reg  dirty_array_0_59; // @[DCache.scala 113:44]
  reg  dirty_array_0_60; // @[DCache.scala 113:44]
  reg  dirty_array_0_61; // @[DCache.scala 113:44]
  reg  dirty_array_0_62; // @[DCache.scala 113:44]
  reg  dirty_array_0_63; // @[DCache.scala 113:44]
  reg  dirty_array_1_0; // @[DCache.scala 114:44]
  reg  dirty_array_1_1; // @[DCache.scala 114:44]
  reg  dirty_array_1_2; // @[DCache.scala 114:44]
  reg  dirty_array_1_3; // @[DCache.scala 114:44]
  reg  dirty_array_1_4; // @[DCache.scala 114:44]
  reg  dirty_array_1_5; // @[DCache.scala 114:44]
  reg  dirty_array_1_6; // @[DCache.scala 114:44]
  reg  dirty_array_1_7; // @[DCache.scala 114:44]
  reg  dirty_array_1_8; // @[DCache.scala 114:44]
  reg  dirty_array_1_9; // @[DCache.scala 114:44]
  reg  dirty_array_1_10; // @[DCache.scala 114:44]
  reg  dirty_array_1_11; // @[DCache.scala 114:44]
  reg  dirty_array_1_12; // @[DCache.scala 114:44]
  reg  dirty_array_1_13; // @[DCache.scala 114:44]
  reg  dirty_array_1_14; // @[DCache.scala 114:44]
  reg  dirty_array_1_15; // @[DCache.scala 114:44]
  reg  dirty_array_1_16; // @[DCache.scala 114:44]
  reg  dirty_array_1_17; // @[DCache.scala 114:44]
  reg  dirty_array_1_18; // @[DCache.scala 114:44]
  reg  dirty_array_1_19; // @[DCache.scala 114:44]
  reg  dirty_array_1_20; // @[DCache.scala 114:44]
  reg  dirty_array_1_21; // @[DCache.scala 114:44]
  reg  dirty_array_1_22; // @[DCache.scala 114:44]
  reg  dirty_array_1_23; // @[DCache.scala 114:44]
  reg  dirty_array_1_24; // @[DCache.scala 114:44]
  reg  dirty_array_1_25; // @[DCache.scala 114:44]
  reg  dirty_array_1_26; // @[DCache.scala 114:44]
  reg  dirty_array_1_27; // @[DCache.scala 114:44]
  reg  dirty_array_1_28; // @[DCache.scala 114:44]
  reg  dirty_array_1_29; // @[DCache.scala 114:44]
  reg  dirty_array_1_30; // @[DCache.scala 114:44]
  reg  dirty_array_1_31; // @[DCache.scala 114:44]
  reg  dirty_array_1_32; // @[DCache.scala 114:44]
  reg  dirty_array_1_33; // @[DCache.scala 114:44]
  reg  dirty_array_1_34; // @[DCache.scala 114:44]
  reg  dirty_array_1_35; // @[DCache.scala 114:44]
  reg  dirty_array_1_36; // @[DCache.scala 114:44]
  reg  dirty_array_1_37; // @[DCache.scala 114:44]
  reg  dirty_array_1_38; // @[DCache.scala 114:44]
  reg  dirty_array_1_39; // @[DCache.scala 114:44]
  reg  dirty_array_1_40; // @[DCache.scala 114:44]
  reg  dirty_array_1_41; // @[DCache.scala 114:44]
  reg  dirty_array_1_42; // @[DCache.scala 114:44]
  reg  dirty_array_1_43; // @[DCache.scala 114:44]
  reg  dirty_array_1_44; // @[DCache.scala 114:44]
  reg  dirty_array_1_45; // @[DCache.scala 114:44]
  reg  dirty_array_1_46; // @[DCache.scala 114:44]
  reg  dirty_array_1_47; // @[DCache.scala 114:44]
  reg  dirty_array_1_48; // @[DCache.scala 114:44]
  reg  dirty_array_1_49; // @[DCache.scala 114:44]
  reg  dirty_array_1_50; // @[DCache.scala 114:44]
  reg  dirty_array_1_51; // @[DCache.scala 114:44]
  reg  dirty_array_1_52; // @[DCache.scala 114:44]
  reg  dirty_array_1_53; // @[DCache.scala 114:44]
  reg  dirty_array_1_54; // @[DCache.scala 114:44]
  reg  dirty_array_1_55; // @[DCache.scala 114:44]
  reg  dirty_array_1_56; // @[DCache.scala 114:44]
  reg  dirty_array_1_57; // @[DCache.scala 114:44]
  reg  dirty_array_1_58; // @[DCache.scala 114:44]
  reg  dirty_array_1_59; // @[DCache.scala 114:44]
  reg  dirty_array_1_60; // @[DCache.scala 114:44]
  reg  dirty_array_1_61; // @[DCache.scala 114:44]
  reg  dirty_array_1_62; // @[DCache.scala 114:44]
  reg  dirty_array_1_63; // @[DCache.scala 114:44]
  reg  valid_array_0_0; // @[DCache.scala 115:44]
  reg  valid_array_0_1; // @[DCache.scala 115:44]
  reg  valid_array_0_2; // @[DCache.scala 115:44]
  reg  valid_array_0_3; // @[DCache.scala 115:44]
  reg  valid_array_0_4; // @[DCache.scala 115:44]
  reg  valid_array_0_5; // @[DCache.scala 115:44]
  reg  valid_array_0_6; // @[DCache.scala 115:44]
  reg  valid_array_0_7; // @[DCache.scala 115:44]
  reg  valid_array_0_8; // @[DCache.scala 115:44]
  reg  valid_array_0_9; // @[DCache.scala 115:44]
  reg  valid_array_0_10; // @[DCache.scala 115:44]
  reg  valid_array_0_11; // @[DCache.scala 115:44]
  reg  valid_array_0_12; // @[DCache.scala 115:44]
  reg  valid_array_0_13; // @[DCache.scala 115:44]
  reg  valid_array_0_14; // @[DCache.scala 115:44]
  reg  valid_array_0_15; // @[DCache.scala 115:44]
  reg  valid_array_0_16; // @[DCache.scala 115:44]
  reg  valid_array_0_17; // @[DCache.scala 115:44]
  reg  valid_array_0_18; // @[DCache.scala 115:44]
  reg  valid_array_0_19; // @[DCache.scala 115:44]
  reg  valid_array_0_20; // @[DCache.scala 115:44]
  reg  valid_array_0_21; // @[DCache.scala 115:44]
  reg  valid_array_0_22; // @[DCache.scala 115:44]
  reg  valid_array_0_23; // @[DCache.scala 115:44]
  reg  valid_array_0_24; // @[DCache.scala 115:44]
  reg  valid_array_0_25; // @[DCache.scala 115:44]
  reg  valid_array_0_26; // @[DCache.scala 115:44]
  reg  valid_array_0_27; // @[DCache.scala 115:44]
  reg  valid_array_0_28; // @[DCache.scala 115:44]
  reg  valid_array_0_29; // @[DCache.scala 115:44]
  reg  valid_array_0_30; // @[DCache.scala 115:44]
  reg  valid_array_0_31; // @[DCache.scala 115:44]
  reg  valid_array_0_32; // @[DCache.scala 115:44]
  reg  valid_array_0_33; // @[DCache.scala 115:44]
  reg  valid_array_0_34; // @[DCache.scala 115:44]
  reg  valid_array_0_35; // @[DCache.scala 115:44]
  reg  valid_array_0_36; // @[DCache.scala 115:44]
  reg  valid_array_0_37; // @[DCache.scala 115:44]
  reg  valid_array_0_38; // @[DCache.scala 115:44]
  reg  valid_array_0_39; // @[DCache.scala 115:44]
  reg  valid_array_0_40; // @[DCache.scala 115:44]
  reg  valid_array_0_41; // @[DCache.scala 115:44]
  reg  valid_array_0_42; // @[DCache.scala 115:44]
  reg  valid_array_0_43; // @[DCache.scala 115:44]
  reg  valid_array_0_44; // @[DCache.scala 115:44]
  reg  valid_array_0_45; // @[DCache.scala 115:44]
  reg  valid_array_0_46; // @[DCache.scala 115:44]
  reg  valid_array_0_47; // @[DCache.scala 115:44]
  reg  valid_array_0_48; // @[DCache.scala 115:44]
  reg  valid_array_0_49; // @[DCache.scala 115:44]
  reg  valid_array_0_50; // @[DCache.scala 115:44]
  reg  valid_array_0_51; // @[DCache.scala 115:44]
  reg  valid_array_0_52; // @[DCache.scala 115:44]
  reg  valid_array_0_53; // @[DCache.scala 115:44]
  reg  valid_array_0_54; // @[DCache.scala 115:44]
  reg  valid_array_0_55; // @[DCache.scala 115:44]
  reg  valid_array_0_56; // @[DCache.scala 115:44]
  reg  valid_array_0_57; // @[DCache.scala 115:44]
  reg  valid_array_0_58; // @[DCache.scala 115:44]
  reg  valid_array_0_59; // @[DCache.scala 115:44]
  reg  valid_array_0_60; // @[DCache.scala 115:44]
  reg  valid_array_0_61; // @[DCache.scala 115:44]
  reg  valid_array_0_62; // @[DCache.scala 115:44]
  reg  valid_array_0_63; // @[DCache.scala 115:44]
  reg  valid_array_1_0; // @[DCache.scala 116:44]
  reg  valid_array_1_1; // @[DCache.scala 116:44]
  reg  valid_array_1_2; // @[DCache.scala 116:44]
  reg  valid_array_1_3; // @[DCache.scala 116:44]
  reg  valid_array_1_4; // @[DCache.scala 116:44]
  reg  valid_array_1_5; // @[DCache.scala 116:44]
  reg  valid_array_1_6; // @[DCache.scala 116:44]
  reg  valid_array_1_7; // @[DCache.scala 116:44]
  reg  valid_array_1_8; // @[DCache.scala 116:44]
  reg  valid_array_1_9; // @[DCache.scala 116:44]
  reg  valid_array_1_10; // @[DCache.scala 116:44]
  reg  valid_array_1_11; // @[DCache.scala 116:44]
  reg  valid_array_1_12; // @[DCache.scala 116:44]
  reg  valid_array_1_13; // @[DCache.scala 116:44]
  reg  valid_array_1_14; // @[DCache.scala 116:44]
  reg  valid_array_1_15; // @[DCache.scala 116:44]
  reg  valid_array_1_16; // @[DCache.scala 116:44]
  reg  valid_array_1_17; // @[DCache.scala 116:44]
  reg  valid_array_1_18; // @[DCache.scala 116:44]
  reg  valid_array_1_19; // @[DCache.scala 116:44]
  reg  valid_array_1_20; // @[DCache.scala 116:44]
  reg  valid_array_1_21; // @[DCache.scala 116:44]
  reg  valid_array_1_22; // @[DCache.scala 116:44]
  reg  valid_array_1_23; // @[DCache.scala 116:44]
  reg  valid_array_1_24; // @[DCache.scala 116:44]
  reg  valid_array_1_25; // @[DCache.scala 116:44]
  reg  valid_array_1_26; // @[DCache.scala 116:44]
  reg  valid_array_1_27; // @[DCache.scala 116:44]
  reg  valid_array_1_28; // @[DCache.scala 116:44]
  reg  valid_array_1_29; // @[DCache.scala 116:44]
  reg  valid_array_1_30; // @[DCache.scala 116:44]
  reg  valid_array_1_31; // @[DCache.scala 116:44]
  reg  valid_array_1_32; // @[DCache.scala 116:44]
  reg  valid_array_1_33; // @[DCache.scala 116:44]
  reg  valid_array_1_34; // @[DCache.scala 116:44]
  reg  valid_array_1_35; // @[DCache.scala 116:44]
  reg  valid_array_1_36; // @[DCache.scala 116:44]
  reg  valid_array_1_37; // @[DCache.scala 116:44]
  reg  valid_array_1_38; // @[DCache.scala 116:44]
  reg  valid_array_1_39; // @[DCache.scala 116:44]
  reg  valid_array_1_40; // @[DCache.scala 116:44]
  reg  valid_array_1_41; // @[DCache.scala 116:44]
  reg  valid_array_1_42; // @[DCache.scala 116:44]
  reg  valid_array_1_43; // @[DCache.scala 116:44]
  reg  valid_array_1_44; // @[DCache.scala 116:44]
  reg  valid_array_1_45; // @[DCache.scala 116:44]
  reg  valid_array_1_46; // @[DCache.scala 116:44]
  reg  valid_array_1_47; // @[DCache.scala 116:44]
  reg  valid_array_1_48; // @[DCache.scala 116:44]
  reg  valid_array_1_49; // @[DCache.scala 116:44]
  reg  valid_array_1_50; // @[DCache.scala 116:44]
  reg  valid_array_1_51; // @[DCache.scala 116:44]
  reg  valid_array_1_52; // @[DCache.scala 116:44]
  reg  valid_array_1_53; // @[DCache.scala 116:44]
  reg  valid_array_1_54; // @[DCache.scala 116:44]
  reg  valid_array_1_55; // @[DCache.scala 116:44]
  reg  valid_array_1_56; // @[DCache.scala 116:44]
  reg  valid_array_1_57; // @[DCache.scala 116:44]
  reg  valid_array_1_58; // @[DCache.scala 116:44]
  reg  valid_array_1_59; // @[DCache.scala 116:44]
  reg  valid_array_1_60; // @[DCache.scala 116:44]
  reg  valid_array_1_61; // @[DCache.scala 116:44]
  reg  valid_array_1_62; // @[DCache.scala 116:44]
  reg  valid_array_1_63; // @[DCache.scala 116:44]
  reg  flush_skip; // @[DCache.scala 122:40]
  reg  flush_cnt_end_latch_en; // @[DCache.scala 125:49]
  wire [5:0] flush_index = value[5:0]; // @[DCache.scala 128:46]
  wire  _GEN_1 = 6'h1 == flush_index ? valid_array_0_1 : valid_array_0_0; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_2 = 6'h2 == flush_index ? valid_array_0_2 : _GEN_1; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_3 = 6'h3 == flush_index ? valid_array_0_3 : _GEN_2; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_4 = 6'h4 == flush_index ? valid_array_0_4 : _GEN_3; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_5 = 6'h5 == flush_index ? valid_array_0_5 : _GEN_4; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_6 = 6'h6 == flush_index ? valid_array_0_6 : _GEN_5; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_7 = 6'h7 == flush_index ? valid_array_0_7 : _GEN_6; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_8 = 6'h8 == flush_index ? valid_array_0_8 : _GEN_7; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_9 = 6'h9 == flush_index ? valid_array_0_9 : _GEN_8; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_10 = 6'ha == flush_index ? valid_array_0_10 : _GEN_9; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_11 = 6'hb == flush_index ? valid_array_0_11 : _GEN_10; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_12 = 6'hc == flush_index ? valid_array_0_12 : _GEN_11; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_13 = 6'hd == flush_index ? valid_array_0_13 : _GEN_12; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_14 = 6'he == flush_index ? valid_array_0_14 : _GEN_13; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_15 = 6'hf == flush_index ? valid_array_0_15 : _GEN_14; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_16 = 6'h10 == flush_index ? valid_array_0_16 : _GEN_15; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_17 = 6'h11 == flush_index ? valid_array_0_17 : _GEN_16; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_18 = 6'h12 == flush_index ? valid_array_0_18 : _GEN_17; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_19 = 6'h13 == flush_index ? valid_array_0_19 : _GEN_18; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_20 = 6'h14 == flush_index ? valid_array_0_20 : _GEN_19; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_21 = 6'h15 == flush_index ? valid_array_0_21 : _GEN_20; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_22 = 6'h16 == flush_index ? valid_array_0_22 : _GEN_21; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_23 = 6'h17 == flush_index ? valid_array_0_23 : _GEN_22; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_24 = 6'h18 == flush_index ? valid_array_0_24 : _GEN_23; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_25 = 6'h19 == flush_index ? valid_array_0_25 : _GEN_24; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_26 = 6'h1a == flush_index ? valid_array_0_26 : _GEN_25; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_27 = 6'h1b == flush_index ? valid_array_0_27 : _GEN_26; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_28 = 6'h1c == flush_index ? valid_array_0_28 : _GEN_27; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_29 = 6'h1d == flush_index ? valid_array_0_29 : _GEN_28; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_30 = 6'h1e == flush_index ? valid_array_0_30 : _GEN_29; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_31 = 6'h1f == flush_index ? valid_array_0_31 : _GEN_30; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_32 = 6'h20 == flush_index ? valid_array_0_32 : _GEN_31; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_33 = 6'h21 == flush_index ? valid_array_0_33 : _GEN_32; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_34 = 6'h22 == flush_index ? valid_array_0_34 : _GEN_33; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_35 = 6'h23 == flush_index ? valid_array_0_35 : _GEN_34; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_36 = 6'h24 == flush_index ? valid_array_0_36 : _GEN_35; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_37 = 6'h25 == flush_index ? valid_array_0_37 : _GEN_36; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_38 = 6'h26 == flush_index ? valid_array_0_38 : _GEN_37; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_39 = 6'h27 == flush_index ? valid_array_0_39 : _GEN_38; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_40 = 6'h28 == flush_index ? valid_array_0_40 : _GEN_39; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_41 = 6'h29 == flush_index ? valid_array_0_41 : _GEN_40; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_42 = 6'h2a == flush_index ? valid_array_0_42 : _GEN_41; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_43 = 6'h2b == flush_index ? valid_array_0_43 : _GEN_42; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_44 = 6'h2c == flush_index ? valid_array_0_44 : _GEN_43; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_45 = 6'h2d == flush_index ? valid_array_0_45 : _GEN_44; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_46 = 6'h2e == flush_index ? valid_array_0_46 : _GEN_45; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_47 = 6'h2f == flush_index ? valid_array_0_47 : _GEN_46; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_48 = 6'h30 == flush_index ? valid_array_0_48 : _GEN_47; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_49 = 6'h31 == flush_index ? valid_array_0_49 : _GEN_48; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_50 = 6'h32 == flush_index ? valid_array_0_50 : _GEN_49; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_51 = 6'h33 == flush_index ? valid_array_0_51 : _GEN_50; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_52 = 6'h34 == flush_index ? valid_array_0_52 : _GEN_51; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_53 = 6'h35 == flush_index ? valid_array_0_53 : _GEN_52; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_54 = 6'h36 == flush_index ? valid_array_0_54 : _GEN_53; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_55 = 6'h37 == flush_index ? valid_array_0_55 : _GEN_54; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_56 = 6'h38 == flush_index ? valid_array_0_56 : _GEN_55; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_57 = 6'h39 == flush_index ? valid_array_0_57 : _GEN_56; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_58 = 6'h3a == flush_index ? valid_array_0_58 : _GEN_57; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_59 = 6'h3b == flush_index ? valid_array_0_59 : _GEN_58; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_60 = 6'h3c == flush_index ? valid_array_0_60 : _GEN_59; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_61 = 6'h3d == flush_index ? valid_array_0_61 : _GEN_60; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_62 = 6'h3e == flush_index ? valid_array_0_62 : _GEN_61; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_63 = 6'h3f == flush_index ? valid_array_0_63 : _GEN_62; // @[DCache.scala 129:57 DCache.scala 129:57]
  wire  _GEN_65 = 6'h1 == flush_index ? valid_array_1_1 : valid_array_1_0; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_66 = 6'h2 == flush_index ? valid_array_1_2 : _GEN_65; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_67 = 6'h3 == flush_index ? valid_array_1_3 : _GEN_66; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_68 = 6'h4 == flush_index ? valid_array_1_4 : _GEN_67; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_69 = 6'h5 == flush_index ? valid_array_1_5 : _GEN_68; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_70 = 6'h6 == flush_index ? valid_array_1_6 : _GEN_69; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_71 = 6'h7 == flush_index ? valid_array_1_7 : _GEN_70; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_72 = 6'h8 == flush_index ? valid_array_1_8 : _GEN_71; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_73 = 6'h9 == flush_index ? valid_array_1_9 : _GEN_72; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_74 = 6'ha == flush_index ? valid_array_1_10 : _GEN_73; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_75 = 6'hb == flush_index ? valid_array_1_11 : _GEN_74; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_76 = 6'hc == flush_index ? valid_array_1_12 : _GEN_75; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_77 = 6'hd == flush_index ? valid_array_1_13 : _GEN_76; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_78 = 6'he == flush_index ? valid_array_1_14 : _GEN_77; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_79 = 6'hf == flush_index ? valid_array_1_15 : _GEN_78; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_80 = 6'h10 == flush_index ? valid_array_1_16 : _GEN_79; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_81 = 6'h11 == flush_index ? valid_array_1_17 : _GEN_80; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_82 = 6'h12 == flush_index ? valid_array_1_18 : _GEN_81; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_83 = 6'h13 == flush_index ? valid_array_1_19 : _GEN_82; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_84 = 6'h14 == flush_index ? valid_array_1_20 : _GEN_83; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_85 = 6'h15 == flush_index ? valid_array_1_21 : _GEN_84; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_86 = 6'h16 == flush_index ? valid_array_1_22 : _GEN_85; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_87 = 6'h17 == flush_index ? valid_array_1_23 : _GEN_86; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_88 = 6'h18 == flush_index ? valid_array_1_24 : _GEN_87; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_89 = 6'h19 == flush_index ? valid_array_1_25 : _GEN_88; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_90 = 6'h1a == flush_index ? valid_array_1_26 : _GEN_89; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_91 = 6'h1b == flush_index ? valid_array_1_27 : _GEN_90; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_92 = 6'h1c == flush_index ? valid_array_1_28 : _GEN_91; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_93 = 6'h1d == flush_index ? valid_array_1_29 : _GEN_92; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_94 = 6'h1e == flush_index ? valid_array_1_30 : _GEN_93; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_95 = 6'h1f == flush_index ? valid_array_1_31 : _GEN_94; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_96 = 6'h20 == flush_index ? valid_array_1_32 : _GEN_95; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_97 = 6'h21 == flush_index ? valid_array_1_33 : _GEN_96; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_98 = 6'h22 == flush_index ? valid_array_1_34 : _GEN_97; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_99 = 6'h23 == flush_index ? valid_array_1_35 : _GEN_98; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_100 = 6'h24 == flush_index ? valid_array_1_36 : _GEN_99; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_101 = 6'h25 == flush_index ? valid_array_1_37 : _GEN_100; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_102 = 6'h26 == flush_index ? valid_array_1_38 : _GEN_101; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_103 = 6'h27 == flush_index ? valid_array_1_39 : _GEN_102; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_104 = 6'h28 == flush_index ? valid_array_1_40 : _GEN_103; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_105 = 6'h29 == flush_index ? valid_array_1_41 : _GEN_104; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_106 = 6'h2a == flush_index ? valid_array_1_42 : _GEN_105; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_107 = 6'h2b == flush_index ? valid_array_1_43 : _GEN_106; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_108 = 6'h2c == flush_index ? valid_array_1_44 : _GEN_107; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_109 = 6'h2d == flush_index ? valid_array_1_45 : _GEN_108; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_110 = 6'h2e == flush_index ? valid_array_1_46 : _GEN_109; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_111 = 6'h2f == flush_index ? valid_array_1_47 : _GEN_110; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_112 = 6'h30 == flush_index ? valid_array_1_48 : _GEN_111; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_113 = 6'h31 == flush_index ? valid_array_1_49 : _GEN_112; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_114 = 6'h32 == flush_index ? valid_array_1_50 : _GEN_113; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_115 = 6'h33 == flush_index ? valid_array_1_51 : _GEN_114; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_116 = 6'h34 == flush_index ? valid_array_1_52 : _GEN_115; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_117 = 6'h35 == flush_index ? valid_array_1_53 : _GEN_116; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_118 = 6'h36 == flush_index ? valid_array_1_54 : _GEN_117; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_119 = 6'h37 == flush_index ? valid_array_1_55 : _GEN_118; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_120 = 6'h38 == flush_index ? valid_array_1_56 : _GEN_119; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_121 = 6'h39 == flush_index ? valid_array_1_57 : _GEN_120; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_122 = 6'h3a == flush_index ? valid_array_1_58 : _GEN_121; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_123 = 6'h3b == flush_index ? valid_array_1_59 : _GEN_122; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_124 = 6'h3c == flush_index ? valid_array_1_60 : _GEN_123; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_125 = 6'h3d == flush_index ? valid_array_1_61 : _GEN_124; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_126 = 6'h3e == flush_index ? valid_array_1_62 : _GEN_125; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  _GEN_127 = 6'h3f == flush_index ? valid_array_1_63 : _GEN_126; // @[DCache.scala 129:126 DCache.scala 129:126]
  wire  flush_hit = _GEN_63 & ~flush_way | _GEN_127 & flush_way; // @[DCache.scala 129:96]
  wire  flush_cnt_end_latch_en_wrap = value == 7'h7f; // @[Counter.scala 72:24]
  wire [6:0] _flush_cnt_end_latch_en_value_T_1 = value + 7'h1; // @[Counter.scala 76:24]
  wire  flush_cnt_rst = curr_state == 4'h6; // @[DCache.scala 260:31]
  wire  _T_13 = curr_state == 4'hc; // @[DCache.scala 256:19]
  wire  flush_cnt_en = curr_state == 4'hc & (flush_skip | maxi4_manager_io_out_finish); // @[DCache.scala 256:29]
  reg  stage1_out_valid; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2mem_sext_flag; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2mem_memory_rd_en; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2mem_memory_we_en; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2wb_intr_exce_ret; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2wb_fencei; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2wb_wb_sel; // @[Reg.scala 27:20]
  reg  stage1_out_bits_data_id2wb_regfile_we_en; // @[Reg.scala 27:20]
  reg [4:0] stage1_out_bits_data_id2wb_regfile_we_addr; // @[Reg.scala 27:20]
  reg [63:0] stage1_out_bits_data_ex2mem_we_data; // @[Reg.scala 27:20]
  reg [63:0] stage1_out_bits_data_ex2wb_result_data; // @[Reg.scala 27:20]
  reg [63:0] stage1_out_bits_wdata; // @[Reg.scala 27:20]
  reg [7:0] stage1_out_bits_wmask; // @[Reg.scala 27:20]
  reg  stage1_out_bits_size_byte; // @[Reg.scala 27:20]
  reg  stage1_out_bits_size_hword; // @[Reg.scala 27:20]
  reg  stage1_out_bits_size_word; // @[Reg.scala 27:20]
  reg  stage1_out_bits_size_dword; // @[Reg.scala 27:20]
  wire  _T_26 = 4'h0 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_27 = stage1_out_bits_data_id2mem_memory_rd_en | stage1_out_bits_data_id2mem_memory_we_en; // @[DCache.scala 358:31]
  wire  addr_underflow = ~stage1_out_bits_addr[31]; // @[DCache.scala 181:60]
  wire [3:0] _GEN_3542 = mmio_manager_io_out_ready ? 4'h7 : 4'h8; // @[DCache.scala 360:30 DCache.scala 360:43 DCache.scala 360:77]
  wire  _GEN_359 = 6'h1 == stage1_index ? dirty_array_1_1 : dirty_array_1_0; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_360 = 6'h2 == stage1_index ? dirty_array_1_2 : _GEN_359; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_361 = 6'h3 == stage1_index ? dirty_array_1_3 : _GEN_360; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_362 = 6'h4 == stage1_index ? dirty_array_1_4 : _GEN_361; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_363 = 6'h5 == stage1_index ? dirty_array_1_5 : _GEN_362; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_364 = 6'h6 == stage1_index ? dirty_array_1_6 : _GEN_363; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_365 = 6'h7 == stage1_index ? dirty_array_1_7 : _GEN_364; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_366 = 6'h8 == stage1_index ? dirty_array_1_8 : _GEN_365; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_367 = 6'h9 == stage1_index ? dirty_array_1_9 : _GEN_366; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_368 = 6'ha == stage1_index ? dirty_array_1_10 : _GEN_367; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_369 = 6'hb == stage1_index ? dirty_array_1_11 : _GEN_368; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_370 = 6'hc == stage1_index ? dirty_array_1_12 : _GEN_369; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_371 = 6'hd == stage1_index ? dirty_array_1_13 : _GEN_370; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_372 = 6'he == stage1_index ? dirty_array_1_14 : _GEN_371; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_373 = 6'hf == stage1_index ? dirty_array_1_15 : _GEN_372; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_374 = 6'h10 == stage1_index ? dirty_array_1_16 : _GEN_373; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_375 = 6'h11 == stage1_index ? dirty_array_1_17 : _GEN_374; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_376 = 6'h12 == stage1_index ? dirty_array_1_18 : _GEN_375; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_377 = 6'h13 == stage1_index ? dirty_array_1_19 : _GEN_376; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_378 = 6'h14 == stage1_index ? dirty_array_1_20 : _GEN_377; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_379 = 6'h15 == stage1_index ? dirty_array_1_21 : _GEN_378; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_380 = 6'h16 == stage1_index ? dirty_array_1_22 : _GEN_379; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_381 = 6'h17 == stage1_index ? dirty_array_1_23 : _GEN_380; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_382 = 6'h18 == stage1_index ? dirty_array_1_24 : _GEN_381; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_383 = 6'h19 == stage1_index ? dirty_array_1_25 : _GEN_382; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_384 = 6'h1a == stage1_index ? dirty_array_1_26 : _GEN_383; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_385 = 6'h1b == stage1_index ? dirty_array_1_27 : _GEN_384; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_386 = 6'h1c == stage1_index ? dirty_array_1_28 : _GEN_385; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_387 = 6'h1d == stage1_index ? dirty_array_1_29 : _GEN_386; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_388 = 6'h1e == stage1_index ? dirty_array_1_30 : _GEN_387; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_389 = 6'h1f == stage1_index ? dirty_array_1_31 : _GEN_388; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_390 = 6'h20 == stage1_index ? dirty_array_1_32 : _GEN_389; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_391 = 6'h21 == stage1_index ? dirty_array_1_33 : _GEN_390; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_392 = 6'h22 == stage1_index ? dirty_array_1_34 : _GEN_391; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_393 = 6'h23 == stage1_index ? dirty_array_1_35 : _GEN_392; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_394 = 6'h24 == stage1_index ? dirty_array_1_36 : _GEN_393; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_395 = 6'h25 == stage1_index ? dirty_array_1_37 : _GEN_394; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_396 = 6'h26 == stage1_index ? dirty_array_1_38 : _GEN_395; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_397 = 6'h27 == stage1_index ? dirty_array_1_39 : _GEN_396; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_398 = 6'h28 == stage1_index ? dirty_array_1_40 : _GEN_397; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_399 = 6'h29 == stage1_index ? dirty_array_1_41 : _GEN_398; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_400 = 6'h2a == stage1_index ? dirty_array_1_42 : _GEN_399; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_401 = 6'h2b == stage1_index ? dirty_array_1_43 : _GEN_400; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_402 = 6'h2c == stage1_index ? dirty_array_1_44 : _GEN_401; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_403 = 6'h2d == stage1_index ? dirty_array_1_45 : _GEN_402; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_404 = 6'h2e == stage1_index ? dirty_array_1_46 : _GEN_403; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_405 = 6'h2f == stage1_index ? dirty_array_1_47 : _GEN_404; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_406 = 6'h30 == stage1_index ? dirty_array_1_48 : _GEN_405; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_407 = 6'h31 == stage1_index ? dirty_array_1_49 : _GEN_406; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_408 = 6'h32 == stage1_index ? dirty_array_1_50 : _GEN_407; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_409 = 6'h33 == stage1_index ? dirty_array_1_51 : _GEN_408; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_410 = 6'h34 == stage1_index ? dirty_array_1_52 : _GEN_409; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_411 = 6'h35 == stage1_index ? dirty_array_1_53 : _GEN_410; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_412 = 6'h36 == stage1_index ? dirty_array_1_54 : _GEN_411; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_413 = 6'h37 == stage1_index ? dirty_array_1_55 : _GEN_412; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_414 = 6'h38 == stage1_index ? dirty_array_1_56 : _GEN_413; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_415 = 6'h39 == stage1_index ? dirty_array_1_57 : _GEN_414; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_416 = 6'h3a == stage1_index ? dirty_array_1_58 : _GEN_415; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_417 = 6'h3b == stage1_index ? dirty_array_1_59 : _GEN_416; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_418 = 6'h3c == stage1_index ? dirty_array_1_60 : _GEN_417; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_419 = 6'h3d == stage1_index ? dirty_array_1_61 : _GEN_418; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_420 = 6'h3e == stage1_index ? dirty_array_1_62 : _GEN_419; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_421 = 6'h3f == stage1_index ? dirty_array_1_63 : _GEN_420; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_423 = 6'h1 == stage1_index ? dirty_array_0_1 : dirty_array_0_0; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_424 = 6'h2 == stage1_index ? dirty_array_0_2 : _GEN_423; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_425 = 6'h3 == stage1_index ? dirty_array_0_3 : _GEN_424; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_426 = 6'h4 == stage1_index ? dirty_array_0_4 : _GEN_425; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_427 = 6'h5 == stage1_index ? dirty_array_0_5 : _GEN_426; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_428 = 6'h6 == stage1_index ? dirty_array_0_6 : _GEN_427; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_429 = 6'h7 == stage1_index ? dirty_array_0_7 : _GEN_428; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_430 = 6'h8 == stage1_index ? dirty_array_0_8 : _GEN_429; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_431 = 6'h9 == stage1_index ? dirty_array_0_9 : _GEN_430; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_432 = 6'ha == stage1_index ? dirty_array_0_10 : _GEN_431; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_433 = 6'hb == stage1_index ? dirty_array_0_11 : _GEN_432; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_434 = 6'hc == stage1_index ? dirty_array_0_12 : _GEN_433; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_435 = 6'hd == stage1_index ? dirty_array_0_13 : _GEN_434; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_436 = 6'he == stage1_index ? dirty_array_0_14 : _GEN_435; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_437 = 6'hf == stage1_index ? dirty_array_0_15 : _GEN_436; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_438 = 6'h10 == stage1_index ? dirty_array_0_16 : _GEN_437; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_439 = 6'h11 == stage1_index ? dirty_array_0_17 : _GEN_438; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_440 = 6'h12 == stage1_index ? dirty_array_0_18 : _GEN_439; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_441 = 6'h13 == stage1_index ? dirty_array_0_19 : _GEN_440; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_442 = 6'h14 == stage1_index ? dirty_array_0_20 : _GEN_441; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_443 = 6'h15 == stage1_index ? dirty_array_0_21 : _GEN_442; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_444 = 6'h16 == stage1_index ? dirty_array_0_22 : _GEN_443; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_445 = 6'h17 == stage1_index ? dirty_array_0_23 : _GEN_444; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_446 = 6'h18 == stage1_index ? dirty_array_0_24 : _GEN_445; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_447 = 6'h19 == stage1_index ? dirty_array_0_25 : _GEN_446; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_448 = 6'h1a == stage1_index ? dirty_array_0_26 : _GEN_447; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_449 = 6'h1b == stage1_index ? dirty_array_0_27 : _GEN_448; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_450 = 6'h1c == stage1_index ? dirty_array_0_28 : _GEN_449; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_451 = 6'h1d == stage1_index ? dirty_array_0_29 : _GEN_450; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_452 = 6'h1e == stage1_index ? dirty_array_0_30 : _GEN_451; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_453 = 6'h1f == stage1_index ? dirty_array_0_31 : _GEN_452; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_454 = 6'h20 == stage1_index ? dirty_array_0_32 : _GEN_453; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_455 = 6'h21 == stage1_index ? dirty_array_0_33 : _GEN_454; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_456 = 6'h22 == stage1_index ? dirty_array_0_34 : _GEN_455; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_457 = 6'h23 == stage1_index ? dirty_array_0_35 : _GEN_456; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_458 = 6'h24 == stage1_index ? dirty_array_0_36 : _GEN_457; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_459 = 6'h25 == stage1_index ? dirty_array_0_37 : _GEN_458; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_460 = 6'h26 == stage1_index ? dirty_array_0_38 : _GEN_459; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_461 = 6'h27 == stage1_index ? dirty_array_0_39 : _GEN_460; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_462 = 6'h28 == stage1_index ? dirty_array_0_40 : _GEN_461; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_463 = 6'h29 == stage1_index ? dirty_array_0_41 : _GEN_462; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_464 = 6'h2a == stage1_index ? dirty_array_0_42 : _GEN_463; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_465 = 6'h2b == stage1_index ? dirty_array_0_43 : _GEN_464; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_466 = 6'h2c == stage1_index ? dirty_array_0_44 : _GEN_465; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_467 = 6'h2d == stage1_index ? dirty_array_0_45 : _GEN_466; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_468 = 6'h2e == stage1_index ? dirty_array_0_46 : _GEN_467; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_469 = 6'h2f == stage1_index ? dirty_array_0_47 : _GEN_468; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_470 = 6'h30 == stage1_index ? dirty_array_0_48 : _GEN_469; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_471 = 6'h31 == stage1_index ? dirty_array_0_49 : _GEN_470; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_472 = 6'h32 == stage1_index ? dirty_array_0_50 : _GEN_471; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_473 = 6'h33 == stage1_index ? dirty_array_0_51 : _GEN_472; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_474 = 6'h34 == stage1_index ? dirty_array_0_52 : _GEN_473; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_475 = 6'h35 == stage1_index ? dirty_array_0_53 : _GEN_474; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_476 = 6'h36 == stage1_index ? dirty_array_0_54 : _GEN_475; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_477 = 6'h37 == stage1_index ? dirty_array_0_55 : _GEN_476; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_478 = 6'h38 == stage1_index ? dirty_array_0_56 : _GEN_477; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_479 = 6'h39 == stage1_index ? dirty_array_0_57 : _GEN_478; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_480 = 6'h3a == stage1_index ? dirty_array_0_58 : _GEN_479; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_481 = 6'h3b == stage1_index ? dirty_array_0_59 : _GEN_480; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_482 = 6'h3c == stage1_index ? dirty_array_0_60 : _GEN_481; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_483 = 6'h3d == stage1_index ? dirty_array_0_61 : _GEN_482; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_484 = 6'h3e == stage1_index ? dirty_array_0_62 : _GEN_483; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  _GEN_485 = 6'h3f == stage1_index ? dirty_array_0_63 : _GEN_484; // @[DCache.scala 182:38 DCache.scala 182:38]
  wire  need_writeback = next_way ? _GEN_421 : _GEN_485; // @[DCache.scala 182:38]
  wire [28:0] stage1_tag = stage1_out_bits_addr[38:10]; // @[DCache.scala 161:54]
  wire [29:0] _GEN_3577 = {{1'd0}, stage1_tag}; // @[DCache.scala 173:52]
  wire  _GEN_230 = 6'h1 == stage1_index ? valid_array_0_1 : valid_array_0_0; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_231 = 6'h2 == stage1_index ? valid_array_0_2 : _GEN_230; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_232 = 6'h3 == stage1_index ? valid_array_0_3 : _GEN_231; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_233 = 6'h4 == stage1_index ? valid_array_0_4 : _GEN_232; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_234 = 6'h5 == stage1_index ? valid_array_0_5 : _GEN_233; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_235 = 6'h6 == stage1_index ? valid_array_0_6 : _GEN_234; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_236 = 6'h7 == stage1_index ? valid_array_0_7 : _GEN_235; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_237 = 6'h8 == stage1_index ? valid_array_0_8 : _GEN_236; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_238 = 6'h9 == stage1_index ? valid_array_0_9 : _GEN_237; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_239 = 6'ha == stage1_index ? valid_array_0_10 : _GEN_238; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_240 = 6'hb == stage1_index ? valid_array_0_11 : _GEN_239; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_241 = 6'hc == stage1_index ? valid_array_0_12 : _GEN_240; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_242 = 6'hd == stage1_index ? valid_array_0_13 : _GEN_241; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_243 = 6'he == stage1_index ? valid_array_0_14 : _GEN_242; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_244 = 6'hf == stage1_index ? valid_array_0_15 : _GEN_243; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_245 = 6'h10 == stage1_index ? valid_array_0_16 : _GEN_244; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_246 = 6'h11 == stage1_index ? valid_array_0_17 : _GEN_245; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_247 = 6'h12 == stage1_index ? valid_array_0_18 : _GEN_246; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_248 = 6'h13 == stage1_index ? valid_array_0_19 : _GEN_247; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_249 = 6'h14 == stage1_index ? valid_array_0_20 : _GEN_248; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_250 = 6'h15 == stage1_index ? valid_array_0_21 : _GEN_249; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_251 = 6'h16 == stage1_index ? valid_array_0_22 : _GEN_250; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_252 = 6'h17 == stage1_index ? valid_array_0_23 : _GEN_251; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_253 = 6'h18 == stage1_index ? valid_array_0_24 : _GEN_252; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_254 = 6'h19 == stage1_index ? valid_array_0_25 : _GEN_253; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_255 = 6'h1a == stage1_index ? valid_array_0_26 : _GEN_254; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_256 = 6'h1b == stage1_index ? valid_array_0_27 : _GEN_255; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_257 = 6'h1c == stage1_index ? valid_array_0_28 : _GEN_256; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_258 = 6'h1d == stage1_index ? valid_array_0_29 : _GEN_257; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_259 = 6'h1e == stage1_index ? valid_array_0_30 : _GEN_258; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_260 = 6'h1f == stage1_index ? valid_array_0_31 : _GEN_259; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_261 = 6'h20 == stage1_index ? valid_array_0_32 : _GEN_260; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_262 = 6'h21 == stage1_index ? valid_array_0_33 : _GEN_261; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_263 = 6'h22 == stage1_index ? valid_array_0_34 : _GEN_262; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_264 = 6'h23 == stage1_index ? valid_array_0_35 : _GEN_263; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_265 = 6'h24 == stage1_index ? valid_array_0_36 : _GEN_264; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_266 = 6'h25 == stage1_index ? valid_array_0_37 : _GEN_265; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_267 = 6'h26 == stage1_index ? valid_array_0_38 : _GEN_266; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_268 = 6'h27 == stage1_index ? valid_array_0_39 : _GEN_267; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_269 = 6'h28 == stage1_index ? valid_array_0_40 : _GEN_268; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_270 = 6'h29 == stage1_index ? valid_array_0_41 : _GEN_269; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_271 = 6'h2a == stage1_index ? valid_array_0_42 : _GEN_270; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_272 = 6'h2b == stage1_index ? valid_array_0_43 : _GEN_271; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_273 = 6'h2c == stage1_index ? valid_array_0_44 : _GEN_272; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_274 = 6'h2d == stage1_index ? valid_array_0_45 : _GEN_273; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_275 = 6'h2e == stage1_index ? valid_array_0_46 : _GEN_274; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_276 = 6'h2f == stage1_index ? valid_array_0_47 : _GEN_275; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_277 = 6'h30 == stage1_index ? valid_array_0_48 : _GEN_276; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_278 = 6'h31 == stage1_index ? valid_array_0_49 : _GEN_277; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_279 = 6'h32 == stage1_index ? valid_array_0_50 : _GEN_278; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_280 = 6'h33 == stage1_index ? valid_array_0_51 : _GEN_279; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_281 = 6'h34 == stage1_index ? valid_array_0_52 : _GEN_280; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_282 = 6'h35 == stage1_index ? valid_array_0_53 : _GEN_281; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_283 = 6'h36 == stage1_index ? valid_array_0_54 : _GEN_282; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_284 = 6'h37 == stage1_index ? valid_array_0_55 : _GEN_283; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_285 = 6'h38 == stage1_index ? valid_array_0_56 : _GEN_284; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_286 = 6'h39 == stage1_index ? valid_array_0_57 : _GEN_285; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_287 = 6'h3a == stage1_index ? valid_array_0_58 : _GEN_286; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_288 = 6'h3b == stage1_index ? valid_array_0_59 : _GEN_287; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_289 = 6'h3c == stage1_index ? valid_array_0_60 : _GEN_288; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_290 = 6'h3d == stage1_index ? valid_array_0_61 : _GEN_289; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_291 = 6'h3e == stage1_index ? valid_array_0_62 : _GEN_290; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  _GEN_292 = 6'h3f == stage1_index ? valid_array_0_63 : _GEN_291; // @[DCache.scala 173:99 DCache.scala 173:99]
  wire  tag0_hit = tag_array_out_0 == _GEN_3577 & _GEN_292; // @[DCache.scala 173:68]
  wire  _GEN_294 = 6'h1 == stage1_index ? valid_array_1_1 : valid_array_1_0; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_295 = 6'h2 == stage1_index ? valid_array_1_2 : _GEN_294; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_296 = 6'h3 == stage1_index ? valid_array_1_3 : _GEN_295; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_297 = 6'h4 == stage1_index ? valid_array_1_4 : _GEN_296; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_298 = 6'h5 == stage1_index ? valid_array_1_5 : _GEN_297; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_299 = 6'h6 == stage1_index ? valid_array_1_6 : _GEN_298; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_300 = 6'h7 == stage1_index ? valid_array_1_7 : _GEN_299; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_301 = 6'h8 == stage1_index ? valid_array_1_8 : _GEN_300; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_302 = 6'h9 == stage1_index ? valid_array_1_9 : _GEN_301; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_303 = 6'ha == stage1_index ? valid_array_1_10 : _GEN_302; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_304 = 6'hb == stage1_index ? valid_array_1_11 : _GEN_303; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_305 = 6'hc == stage1_index ? valid_array_1_12 : _GEN_304; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_306 = 6'hd == stage1_index ? valid_array_1_13 : _GEN_305; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_307 = 6'he == stage1_index ? valid_array_1_14 : _GEN_306; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_308 = 6'hf == stage1_index ? valid_array_1_15 : _GEN_307; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_309 = 6'h10 == stage1_index ? valid_array_1_16 : _GEN_308; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_310 = 6'h11 == stage1_index ? valid_array_1_17 : _GEN_309; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_311 = 6'h12 == stage1_index ? valid_array_1_18 : _GEN_310; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_312 = 6'h13 == stage1_index ? valid_array_1_19 : _GEN_311; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_313 = 6'h14 == stage1_index ? valid_array_1_20 : _GEN_312; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_314 = 6'h15 == stage1_index ? valid_array_1_21 : _GEN_313; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_315 = 6'h16 == stage1_index ? valid_array_1_22 : _GEN_314; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_316 = 6'h17 == stage1_index ? valid_array_1_23 : _GEN_315; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_317 = 6'h18 == stage1_index ? valid_array_1_24 : _GEN_316; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_318 = 6'h19 == stage1_index ? valid_array_1_25 : _GEN_317; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_319 = 6'h1a == stage1_index ? valid_array_1_26 : _GEN_318; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_320 = 6'h1b == stage1_index ? valid_array_1_27 : _GEN_319; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_321 = 6'h1c == stage1_index ? valid_array_1_28 : _GEN_320; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_322 = 6'h1d == stage1_index ? valid_array_1_29 : _GEN_321; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_323 = 6'h1e == stage1_index ? valid_array_1_30 : _GEN_322; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_324 = 6'h1f == stage1_index ? valid_array_1_31 : _GEN_323; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_325 = 6'h20 == stage1_index ? valid_array_1_32 : _GEN_324; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_326 = 6'h21 == stage1_index ? valid_array_1_33 : _GEN_325; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_327 = 6'h22 == stage1_index ? valid_array_1_34 : _GEN_326; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_328 = 6'h23 == stage1_index ? valid_array_1_35 : _GEN_327; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_329 = 6'h24 == stage1_index ? valid_array_1_36 : _GEN_328; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_330 = 6'h25 == stage1_index ? valid_array_1_37 : _GEN_329; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_331 = 6'h26 == stage1_index ? valid_array_1_38 : _GEN_330; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_332 = 6'h27 == stage1_index ? valid_array_1_39 : _GEN_331; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_333 = 6'h28 == stage1_index ? valid_array_1_40 : _GEN_332; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_334 = 6'h29 == stage1_index ? valid_array_1_41 : _GEN_333; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_335 = 6'h2a == stage1_index ? valid_array_1_42 : _GEN_334; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_336 = 6'h2b == stage1_index ? valid_array_1_43 : _GEN_335; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_337 = 6'h2c == stage1_index ? valid_array_1_44 : _GEN_336; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_338 = 6'h2d == stage1_index ? valid_array_1_45 : _GEN_337; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_339 = 6'h2e == stage1_index ? valid_array_1_46 : _GEN_338; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_340 = 6'h2f == stage1_index ? valid_array_1_47 : _GEN_339; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_341 = 6'h30 == stage1_index ? valid_array_1_48 : _GEN_340; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_342 = 6'h31 == stage1_index ? valid_array_1_49 : _GEN_341; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_343 = 6'h32 == stage1_index ? valid_array_1_50 : _GEN_342; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_344 = 6'h33 == stage1_index ? valid_array_1_51 : _GEN_343; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_345 = 6'h34 == stage1_index ? valid_array_1_52 : _GEN_344; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_346 = 6'h35 == stage1_index ? valid_array_1_53 : _GEN_345; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_347 = 6'h36 == stage1_index ? valid_array_1_54 : _GEN_346; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_348 = 6'h37 == stage1_index ? valid_array_1_55 : _GEN_347; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_349 = 6'h38 == stage1_index ? valid_array_1_56 : _GEN_348; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_350 = 6'h39 == stage1_index ? valid_array_1_57 : _GEN_349; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_351 = 6'h3a == stage1_index ? valid_array_1_58 : _GEN_350; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_352 = 6'h3b == stage1_index ? valid_array_1_59 : _GEN_351; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_353 = 6'h3c == stage1_index ? valid_array_1_60 : _GEN_352; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_354 = 6'h3d == stage1_index ? valid_array_1_61 : _GEN_353; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_355 = 6'h3e == stage1_index ? valid_array_1_62 : _GEN_354; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  _GEN_356 = 6'h3f == stage1_index ? valid_array_1_63 : _GEN_355; // @[DCache.scala 174:99 DCache.scala 174:99]
  wire  tag1_hit = tag_array_out_1 == _GEN_3577 & _GEN_356; // @[DCache.scala 174:68]
  wire  miss = ~(tag0_hit | tag1_hit); // @[DCache.scala 180:35]
  wire  _T_28 = need_writeback & miss; // @[DCache.scala 361:37]
  wire [3:0] _GEN_3543 = maxi4_manager_io_out_ready ? 4'h4 : 4'h5; // @[DCache.scala 362:30 DCache.scala 362:43 DCache.scala 362:83]
  wire [3:0] _GEN_3544 = maxi4_manager_io_out_ready ? 4'h2 : 4'h3; // @[DCache.scala 364:30 DCache.scala 364:43 DCache.scala 364:78]
  wire [3:0] _GEN_3545 = stage1_out_bits_data_id2mem_memory_we_en ? 4'h1 : curr_state; // @[DCache.scala 366:34 DCache.scala 366:47 DCache.scala 354:14]
  wire [3:0] _GEN_3546 = stage1_out_bits_data_id2mem_memory_rd_en ? 4'h0 : _GEN_3545; // @[DCache.scala 365:34 DCache.scala 365:47]
  wire [3:0] _GEN_3547 = miss ? _GEN_3544 : _GEN_3546; // @[DCache.scala 363:27]
  wire [3:0] _GEN_3548 = need_writeback & miss ? _GEN_3543 : _GEN_3547; // @[DCache.scala 361:44]
  wire [3:0] _GEN_3549 = addr_underflow ? _GEN_3542 : _GEN_3548; // @[DCache.scala 359:32]
  wire [3:0] _GEN_3550 = stage1_out_bits_data_id2mem_memory_rd_en | stage1_out_bits_data_id2mem_memory_we_en ? _GEN_3549
     : curr_state; // @[DCache.scala 358:45 DCache.scala 354:14]
  wire [3:0] _GEN_3551 = io_prev_bits_flush ? 4'h9 : _GEN_3550; // @[DCache.scala 357:31 DCache.scala 357:44]
  wire  _T_29 = 4'h1 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_30 = 4'h3 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3552 = maxi4_manager_io_out_ready ? 4'h2 : curr_state; // @[DCache.scala 370:34 DCache.scala 370:47 DCache.scala 354:14]
  wire  _T_31 = 4'h5 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3553 = maxi4_manager_io_out_ready ? 4'h4 : curr_state; // @[DCache.scala 371:34 DCache.scala 371:47 DCache.scala 354:14]
  wire  _T_32 = 4'h8 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3554 = mmio_manager_io_out_ready ? 4'h7 : curr_state; // @[DCache.scala 372:34 DCache.scala 372:47 DCache.scala 354:14]
  wire  _T_33 = 4'h2 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3555 = maxi4_manager_io_out_finish ? 4'h6 : curr_state; // @[DCache.scala 374:24 DCache.scala 374:37 DCache.scala 354:14]
  wire  _T_34 = 4'h7 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3556 = mmio_manager_io_out_finish ? 4'h6 : curr_state; // @[DCache.scala 377:24 DCache.scala 377:37 DCache.scala 354:14]
  wire  _T_35 = 4'h4 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3557 = maxi4_manager_io_out_finish ? 4'h3 : curr_state; // @[DCache.scala 380:24 DCache.scala 380:37 DCache.scala 354:14]
  wire  _T_36 = 4'h6 == curr_state; // @[Conditional.scala 37:30]
  wire  _T_37 = 4'h9 == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3559 = flush_hit ? 4'ha : 4'hc; // @[DCache.scala 384:22 DCache.scala 384:35 DCache.scala 385:32]
  wire  _T_38 = 4'ha == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3560 = maxi4_manager_io_out_ready ? 4'hb : curr_state; // @[DCache.scala 388:24 DCache.scala 388:37 DCache.scala 354:14]
  wire  _T_39 = 4'hb == curr_state; // @[Conditional.scala 37:30]
  wire  _T_40 = 4'hc == curr_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_3561 = maxi4_manager_io_out_finish ? 4'h9 : curr_state; // @[DCache.scala 396:31 DCache.scala 396:44 DCache.scala 354:14]
  wire [3:0] _GEN_3562 = flush_skip ? 4'h9 : _GEN_3561; // @[DCache.scala 395:30 DCache.scala 395:43]
  wire [3:0] _GEN_3563 = flush_cnt_end_latch_en ? 4'h6 : _GEN_3562; // @[DCache.scala 394:35 DCache.scala 394:48]
  wire [3:0] _GEN_3564 = _T_40 ? _GEN_3563 : curr_state; // @[Conditional.scala 39:67 DCache.scala 354:14]
  wire [3:0] _GEN_3565 = _T_39 ? 4'hc : _GEN_3564; // @[Conditional.scala 39:67 DCache.scala 391:18]
  wire [3:0] _GEN_3566 = _T_38 ? _GEN_3560 : _GEN_3565; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3567 = _T_37 ? _GEN_3559 : _GEN_3566; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3568 = _T_36 ? 4'h0 : _GEN_3567; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3569 = _T_35 ? _GEN_3557 : _GEN_3568; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3570 = _T_34 ? _GEN_3556 : _GEN_3569; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3571 = _T_33 ? _GEN_3555 : _GEN_3570; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3572 = _T_32 ? _GEN_3554 : _GEN_3571; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3573 = _T_31 ? _GEN_3553 : _GEN_3572; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3574 = _T_30 ? _GEN_3552 : _GEN_3573; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_3575 = _T_29 ? 4'h6 : _GEN_3574; // @[Conditional.scala 39:67 DCache.scala 369:27]
  wire [3:0] next_state = _T_26 ? _GEN_3551 : _GEN_3575; // @[Conditional.scala 40:58]
  wire  go_on = next_state == 4'h0; // @[DCache.scala 185:46]
  wire [5:0] prev_index = io_prev_bits_addr[9:4]; // @[DCache.scala 158:48]
  wire  hit_reg_x8 = curr_state == 4'h0; // @[DCache.scala 175:98]
  wire [127:0] writeback_data = next_way ? io_sram5_rdata : io_sram4_rdata; // @[DCache.scala 176:38]
  wire [3:0] addr_array_0_lo = stage1_out_bits_addr[3:0]; // @[DCache.scala 177:90]
  wire [39:0] _addr_array_0_T = {tag_array_out_0,stage1_index,addr_array_0_lo}; // @[Cat.scala 30:58]
  wire [31:0] addr_array_0 = _addr_array_0_T[31:0]; // @[DCache.scala 177:97]
  wire [39:0] _addr_array_1_T = {tag_array_out_1,stage1_index,addr_array_0_lo}; // @[Cat.scala 30:58]
  wire [31:0] addr_array_1 = _addr_array_1_T[31:0]; // @[DCache.scala 178:97]
  wire [31:0] writeback_addr = next_way ? addr_array_1 : addr_array_0; // @[DCache.scala 179:38]
  wire [39:0] _flush_wb_addr_T = {tag_array_out_1,flush_index,4'h0}; // @[Cat.scala 30:58]
  wire [39:0] _flush_wb_addr_T_1 = {tag_array_out_0,flush_index,4'h0}; // @[Cat.scala 30:58]
  wire [39:0] flush_wb_addr = flush_way ? _flush_wb_addr_T : _flush_wb_addr_T_1; // @[DCache.scala 183:38]
  wire [127:0] flush_wb_data = flush_way ? io_sram5_rdata : io_sram4_rdata; // @[DCache.scala 184:38]
  wire [127:0] _cache_line_data_out_T = tag1_hit ? io_sram5_rdata : 128'h0; // @[Mux.scala 98:16]
  wire [127:0] cache_line_data_out = tag0_hit ? io_sram4_rdata : _cache_line_data_out_T; // @[Mux.scala 98:16]
  wire  _T = curr_state == 4'ha; // @[DCache.scala 205:19]
  wire  _GEN_488 = _T_28 ? 1'h0 : miss; // @[DCache.scala 211:36 DCache.scala 203:14]
  wire  _GEN_489 = _T_27 & _T_28; // @[DCache.scala 210:44 DCache.scala 204:14]
  wire  _GEN_490 = _T_27 & _GEN_488; // @[DCache.scala 210:44 DCache.scala 203:14]
  wire  _GEN_491 = addr_underflow ? 1'h0 : _GEN_489; // @[DCache.scala 207:28 DCache.scala 208:20]
  wire  _GEN_492 = addr_underflow ? 1'h0 : _GEN_490; // @[DCache.scala 207:28 DCache.scala 209:20]
  wire  _T_4 = curr_state == 4'h3; // @[DCache.scala 215:26]
  wire  _GEN_494 = curr_state == 4'h5 | _T; // @[DCache.scala 216:37 DCache.scala 216:50]
  wire  _GEN_496 = curr_state == 4'h3 ? 1'h0 : _GEN_494; // @[DCache.scala 215:37 DCache.scala 204:14]
  wire  _GEN_497 = hit_reg_x8 ? _GEN_491 : _GEN_496; // @[DCache.scala 206:38]
  wire  _GEN_498 = hit_reg_x8 ? _GEN_492 : _T_4; // @[DCache.scala 206:38]
  wire  _maxi4_manager_io_in_addr_T_2 = hit_reg_x8 & need_writeback; // @[DCache.scala 221:29]
  wire [38:0] _maxi4_manager_io_in_addr_T_3 = _maxi4_manager_io_in_addr_T_2 ? {{7'd0}, writeback_addr} :
    stage1_out_bits_addr; // @[Mux.scala 98:16]
  wire [39:0] _maxi4_manager_io_in_addr_T_4 = _T ? flush_wb_addr : {{1'd0}, _maxi4_manager_io_in_addr_T_3}; // @[Mux.scala 98:16]
  wire [34:0] maxi4_manager_io_in_addr_hi = _maxi4_manager_io_in_addr_T_4[38:4]; // @[DCache.scala 222:5]
  wire [38:0] _maxi4_manager_io_in_addr_T_5 = {maxi4_manager_io_in_addr_hi,4'h0}; // @[Cat.scala 30:58]
  wire [127:0] _maxi4_manager_io_in_data_T_3 = _maxi4_manager_io_in_addr_T_2 ? writeback_data : {{64'd0},
    stage1_out_bits_wdata}; // @[Mux.scala 98:16]
  wire  _GEN_503 = stage1_out_bits_data_id2mem_memory_we_en ? 1'h0 : stage1_out_bits_data_id2mem_memory_rd_en; // @[DCache.scala 232:29 DCache.scala 229:14]
  wire  _GEN_504 = curr_state == 4'h8 & stage1_out_bits_data_id2mem_memory_we_en; // @[DCache.scala 235:37 DCache.scala 230:14]
  wire  _GEN_505 = curr_state == 4'h8 & _GEN_503; // @[DCache.scala 235:37 DCache.scala 229:14]
  wire  _T_10 = curr_state == 4'h9; // @[DCache.scala 247:19]
  wire  _GEN_508 = next_state == 4'ha ? 1'h0 : flush_skip; // @[DCache.scala 250:38 DCache.scala 251:18 DCache.scala 122:40]
  wire  _GEN_509 = next_state == 4'hc | _GEN_508; // @[DCache.scala 248:31 DCache.scala 249:18]
  wire  _GEN_3579 = 6'h0 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_512 = 6'h0 == stage1_index | lru_list_0; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3580 = 6'h1 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_513 = 6'h1 == stage1_index | lru_list_1; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3581 = 6'h2 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_514 = 6'h2 == stage1_index | lru_list_2; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3582 = 6'h3 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_515 = 6'h3 == stage1_index | lru_list_3; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3583 = 6'h4 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_516 = 6'h4 == stage1_index | lru_list_4; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3584 = 6'h5 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_517 = 6'h5 == stage1_index | lru_list_5; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3585 = 6'h6 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_518 = 6'h6 == stage1_index | lru_list_6; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3586 = 6'h7 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_519 = 6'h7 == stage1_index | lru_list_7; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3587 = 6'h8 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_520 = 6'h8 == stage1_index | lru_list_8; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3588 = 6'h9 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_521 = 6'h9 == stage1_index | lru_list_9; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3589 = 6'ha == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_522 = 6'ha == stage1_index | lru_list_10; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3590 = 6'hb == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_523 = 6'hb == stage1_index | lru_list_11; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3591 = 6'hc == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_524 = 6'hc == stage1_index | lru_list_12; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3592 = 6'hd == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_525 = 6'hd == stage1_index | lru_list_13; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3593 = 6'he == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_526 = 6'he == stage1_index | lru_list_14; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3594 = 6'hf == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_527 = 6'hf == stage1_index | lru_list_15; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3595 = 6'h10 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_528 = 6'h10 == stage1_index | lru_list_16; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3596 = 6'h11 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_529 = 6'h11 == stage1_index | lru_list_17; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3597 = 6'h12 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_530 = 6'h12 == stage1_index | lru_list_18; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3598 = 6'h13 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_531 = 6'h13 == stage1_index | lru_list_19; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3599 = 6'h14 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_532 = 6'h14 == stage1_index | lru_list_20; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3600 = 6'h15 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_533 = 6'h15 == stage1_index | lru_list_21; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3601 = 6'h16 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_534 = 6'h16 == stage1_index | lru_list_22; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3602 = 6'h17 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_535 = 6'h17 == stage1_index | lru_list_23; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3603 = 6'h18 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_536 = 6'h18 == stage1_index | lru_list_24; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3604 = 6'h19 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_537 = 6'h19 == stage1_index | lru_list_25; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3605 = 6'h1a == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_538 = 6'h1a == stage1_index | lru_list_26; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3606 = 6'h1b == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_539 = 6'h1b == stage1_index | lru_list_27; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3607 = 6'h1c == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_540 = 6'h1c == stage1_index | lru_list_28; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3608 = 6'h1d == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_541 = 6'h1d == stage1_index | lru_list_29; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3609 = 6'h1e == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_542 = 6'h1e == stage1_index | lru_list_30; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3610 = 6'h1f == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_543 = 6'h1f == stage1_index | lru_list_31; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3611 = 6'h20 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_544 = 6'h20 == stage1_index | lru_list_32; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3612 = 6'h21 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_545 = 6'h21 == stage1_index | lru_list_33; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3613 = 6'h22 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_546 = 6'h22 == stage1_index | lru_list_34; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3614 = 6'h23 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_547 = 6'h23 == stage1_index | lru_list_35; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3615 = 6'h24 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_548 = 6'h24 == stage1_index | lru_list_36; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3616 = 6'h25 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_549 = 6'h25 == stage1_index | lru_list_37; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3617 = 6'h26 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_550 = 6'h26 == stage1_index | lru_list_38; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3618 = 6'h27 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_551 = 6'h27 == stage1_index | lru_list_39; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3619 = 6'h28 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_552 = 6'h28 == stage1_index | lru_list_40; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3620 = 6'h29 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_553 = 6'h29 == stage1_index | lru_list_41; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3621 = 6'h2a == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_554 = 6'h2a == stage1_index | lru_list_42; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3622 = 6'h2b == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_555 = 6'h2b == stage1_index | lru_list_43; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3623 = 6'h2c == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_556 = 6'h2c == stage1_index | lru_list_44; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3624 = 6'h2d == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_557 = 6'h2d == stage1_index | lru_list_45; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3625 = 6'h2e == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_558 = 6'h2e == stage1_index | lru_list_46; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3626 = 6'h2f == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_559 = 6'h2f == stage1_index | lru_list_47; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3627 = 6'h30 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_560 = 6'h30 == stage1_index | lru_list_48; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3628 = 6'h31 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_561 = 6'h31 == stage1_index | lru_list_49; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3629 = 6'h32 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_562 = 6'h32 == stage1_index | lru_list_50; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3630 = 6'h33 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_563 = 6'h33 == stage1_index | lru_list_51; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3631 = 6'h34 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_564 = 6'h34 == stage1_index | lru_list_52; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3632 = 6'h35 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_565 = 6'h35 == stage1_index | lru_list_53; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3633 = 6'h36 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_566 = 6'h36 == stage1_index | lru_list_54; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3634 = 6'h37 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_567 = 6'h37 == stage1_index | lru_list_55; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3635 = 6'h38 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_568 = 6'h38 == stage1_index | lru_list_56; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3636 = 6'h39 == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_569 = 6'h39 == stage1_index | lru_list_57; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3637 = 6'h3a == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_570 = 6'h3a == stage1_index | lru_list_58; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3638 = 6'h3b == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_571 = 6'h3b == stage1_index | lru_list_59; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3639 = 6'h3c == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_572 = 6'h3c == stage1_index | lru_list_60; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3640 = 6'h3d == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_573 = 6'h3d == stage1_index | lru_list_61; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3641 = 6'h3e == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_574 = 6'h3e == stage1_index | lru_list_62; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_3642 = 6'h3f == stage1_index; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire  _GEN_575 = 6'h3f == stage1_index | lru_list_63; // @[DCache.scala 271:32 DCache.scala 271:32 DCache.scala 118:35]
  wire [125:0] tag_array_in = {{97'd0}, stage1_tag}; // @[DCache.scala 197:38 DCache.scala 462:16]
  wire [127:0] x12 = {2'h0,tag_array_in}; // @[Cat.scala 30:58]
  wire  _GEN_576 = _GEN_3579 | valid_array_1_0; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_577 = _GEN_3580 | valid_array_1_1; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_578 = _GEN_3581 | valid_array_1_2; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_579 = _GEN_3582 | valid_array_1_3; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_580 = _GEN_3583 | valid_array_1_4; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_581 = _GEN_3584 | valid_array_1_5; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_582 = _GEN_3585 | valid_array_1_6; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_583 = _GEN_3586 | valid_array_1_7; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_584 = _GEN_3587 | valid_array_1_8; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_585 = _GEN_3588 | valid_array_1_9; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_586 = _GEN_3589 | valid_array_1_10; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_587 = _GEN_3590 | valid_array_1_11; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_588 = _GEN_3591 | valid_array_1_12; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_589 = _GEN_3592 | valid_array_1_13; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_590 = _GEN_3593 | valid_array_1_14; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_591 = _GEN_3594 | valid_array_1_15; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_592 = _GEN_3595 | valid_array_1_16; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_593 = _GEN_3596 | valid_array_1_17; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_594 = _GEN_3597 | valid_array_1_18; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_595 = _GEN_3598 | valid_array_1_19; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_596 = _GEN_3599 | valid_array_1_20; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_597 = _GEN_3600 | valid_array_1_21; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_598 = _GEN_3601 | valid_array_1_22; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_599 = _GEN_3602 | valid_array_1_23; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_600 = _GEN_3603 | valid_array_1_24; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_601 = _GEN_3604 | valid_array_1_25; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_602 = _GEN_3605 | valid_array_1_26; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_603 = _GEN_3606 | valid_array_1_27; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_604 = _GEN_3607 | valid_array_1_28; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_605 = _GEN_3608 | valid_array_1_29; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_606 = _GEN_3609 | valid_array_1_30; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_607 = _GEN_3610 | valid_array_1_31; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_608 = _GEN_3611 | valid_array_1_32; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_609 = _GEN_3612 | valid_array_1_33; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_610 = _GEN_3613 | valid_array_1_34; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_611 = _GEN_3614 | valid_array_1_35; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_612 = _GEN_3615 | valid_array_1_36; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_613 = _GEN_3616 | valid_array_1_37; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_614 = _GEN_3617 | valid_array_1_38; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_615 = _GEN_3618 | valid_array_1_39; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_616 = _GEN_3619 | valid_array_1_40; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_617 = _GEN_3620 | valid_array_1_41; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_618 = _GEN_3621 | valid_array_1_42; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_619 = _GEN_3622 | valid_array_1_43; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_620 = _GEN_3623 | valid_array_1_44; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_621 = _GEN_3624 | valid_array_1_45; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_622 = _GEN_3625 | valid_array_1_46; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_623 = _GEN_3626 | valid_array_1_47; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_624 = _GEN_3627 | valid_array_1_48; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_625 = _GEN_3628 | valid_array_1_49; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_626 = _GEN_3629 | valid_array_1_50; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_627 = _GEN_3630 | valid_array_1_51; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_628 = _GEN_3631 | valid_array_1_52; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_629 = _GEN_3632 | valid_array_1_53; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_630 = _GEN_3633 | valid_array_1_54; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_631 = _GEN_3634 | valid_array_1_55; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_632 = _GEN_3635 | valid_array_1_56; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_633 = _GEN_3636 | valid_array_1_57; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_634 = _GEN_3637 | valid_array_1_58; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_635 = _GEN_3638 | valid_array_1_59; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_636 = _GEN_3639 | valid_array_1_60; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_637 = _GEN_3640 | valid_array_1_61; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_638 = _GEN_3641 | valid_array_1_62; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _GEN_639 = _GEN_3642 | valid_array_1_63; // @[DCache.scala 275:37 DCache.scala 275:37 DCache.scala 116:44]
  wire  _dirty_array_in_T_2 = _T_16 & stage1_out_bits_data_id2mem_memory_we_en; // @[DCache.scala 465:27]
  wire  dirty_array_in = _T_19 | _dirty_array_in_T_2; // @[Mux.scala 98:16]
  wire  _GEN_640 = 6'h0 == stage1_index ? dirty_array_in : dirty_array_1_0; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_641 = 6'h1 == stage1_index ? dirty_array_in : dirty_array_1_1; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_642 = 6'h2 == stage1_index ? dirty_array_in : dirty_array_1_2; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_643 = 6'h3 == stage1_index ? dirty_array_in : dirty_array_1_3; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_644 = 6'h4 == stage1_index ? dirty_array_in : dirty_array_1_4; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_645 = 6'h5 == stage1_index ? dirty_array_in : dirty_array_1_5; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_646 = 6'h6 == stage1_index ? dirty_array_in : dirty_array_1_6; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_647 = 6'h7 == stage1_index ? dirty_array_in : dirty_array_1_7; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_648 = 6'h8 == stage1_index ? dirty_array_in : dirty_array_1_8; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_649 = 6'h9 == stage1_index ? dirty_array_in : dirty_array_1_9; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_650 = 6'ha == stage1_index ? dirty_array_in : dirty_array_1_10; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_651 = 6'hb == stage1_index ? dirty_array_in : dirty_array_1_11; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_652 = 6'hc == stage1_index ? dirty_array_in : dirty_array_1_12; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_653 = 6'hd == stage1_index ? dirty_array_in : dirty_array_1_13; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_654 = 6'he == stage1_index ? dirty_array_in : dirty_array_1_14; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_655 = 6'hf == stage1_index ? dirty_array_in : dirty_array_1_15; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_656 = 6'h10 == stage1_index ? dirty_array_in : dirty_array_1_16; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_657 = 6'h11 == stage1_index ? dirty_array_in : dirty_array_1_17; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_658 = 6'h12 == stage1_index ? dirty_array_in : dirty_array_1_18; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_659 = 6'h13 == stage1_index ? dirty_array_in : dirty_array_1_19; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_660 = 6'h14 == stage1_index ? dirty_array_in : dirty_array_1_20; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_661 = 6'h15 == stage1_index ? dirty_array_in : dirty_array_1_21; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_662 = 6'h16 == stage1_index ? dirty_array_in : dirty_array_1_22; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_663 = 6'h17 == stage1_index ? dirty_array_in : dirty_array_1_23; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_664 = 6'h18 == stage1_index ? dirty_array_in : dirty_array_1_24; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_665 = 6'h19 == stage1_index ? dirty_array_in : dirty_array_1_25; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_666 = 6'h1a == stage1_index ? dirty_array_in : dirty_array_1_26; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_667 = 6'h1b == stage1_index ? dirty_array_in : dirty_array_1_27; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_668 = 6'h1c == stage1_index ? dirty_array_in : dirty_array_1_28; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_669 = 6'h1d == stage1_index ? dirty_array_in : dirty_array_1_29; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_670 = 6'h1e == stage1_index ? dirty_array_in : dirty_array_1_30; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_671 = 6'h1f == stage1_index ? dirty_array_in : dirty_array_1_31; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_672 = 6'h20 == stage1_index ? dirty_array_in : dirty_array_1_32; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_673 = 6'h21 == stage1_index ? dirty_array_in : dirty_array_1_33; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_674 = 6'h22 == stage1_index ? dirty_array_in : dirty_array_1_34; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_675 = 6'h23 == stage1_index ? dirty_array_in : dirty_array_1_35; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_676 = 6'h24 == stage1_index ? dirty_array_in : dirty_array_1_36; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_677 = 6'h25 == stage1_index ? dirty_array_in : dirty_array_1_37; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_678 = 6'h26 == stage1_index ? dirty_array_in : dirty_array_1_38; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_679 = 6'h27 == stage1_index ? dirty_array_in : dirty_array_1_39; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_680 = 6'h28 == stage1_index ? dirty_array_in : dirty_array_1_40; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_681 = 6'h29 == stage1_index ? dirty_array_in : dirty_array_1_41; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_682 = 6'h2a == stage1_index ? dirty_array_in : dirty_array_1_42; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_683 = 6'h2b == stage1_index ? dirty_array_in : dirty_array_1_43; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_684 = 6'h2c == stage1_index ? dirty_array_in : dirty_array_1_44; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_685 = 6'h2d == stage1_index ? dirty_array_in : dirty_array_1_45; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_686 = 6'h2e == stage1_index ? dirty_array_in : dirty_array_1_46; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_687 = 6'h2f == stage1_index ? dirty_array_in : dirty_array_1_47; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_688 = 6'h30 == stage1_index ? dirty_array_in : dirty_array_1_48; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_689 = 6'h31 == stage1_index ? dirty_array_in : dirty_array_1_49; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_690 = 6'h32 == stage1_index ? dirty_array_in : dirty_array_1_50; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_691 = 6'h33 == stage1_index ? dirty_array_in : dirty_array_1_51; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_692 = 6'h34 == stage1_index ? dirty_array_in : dirty_array_1_52; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_693 = 6'h35 == stage1_index ? dirty_array_in : dirty_array_1_53; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_694 = 6'h36 == stage1_index ? dirty_array_in : dirty_array_1_54; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_695 = 6'h37 == stage1_index ? dirty_array_in : dirty_array_1_55; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_696 = 6'h38 == stage1_index ? dirty_array_in : dirty_array_1_56; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_697 = 6'h39 == stage1_index ? dirty_array_in : dirty_array_1_57; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_698 = 6'h3a == stage1_index ? dirty_array_in : dirty_array_1_58; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_699 = 6'h3b == stage1_index ? dirty_array_in : dirty_array_1_59; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_700 = 6'h3c == stage1_index ? dirty_array_in : dirty_array_1_60; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_701 = 6'h3d == stage1_index ? dirty_array_in : dirty_array_1_61; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_702 = 6'h3e == stage1_index ? dirty_array_in : dirty_array_1_62; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_703 = 6'h3f == stage1_index ? dirty_array_in : dirty_array_1_63; // @[DCache.scala 276:37 DCache.scala 276:37 DCache.scala 114:44]
  wire  _GEN_704 = 6'h0 == stage1_index ? 1'h0 : lru_list_0; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_705 = 6'h1 == stage1_index ? 1'h0 : lru_list_1; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_706 = 6'h2 == stage1_index ? 1'h0 : lru_list_2; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_707 = 6'h3 == stage1_index ? 1'h0 : lru_list_3; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_708 = 6'h4 == stage1_index ? 1'h0 : lru_list_4; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_709 = 6'h5 == stage1_index ? 1'h0 : lru_list_5; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_710 = 6'h6 == stage1_index ? 1'h0 : lru_list_6; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_711 = 6'h7 == stage1_index ? 1'h0 : lru_list_7; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_712 = 6'h8 == stage1_index ? 1'h0 : lru_list_8; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_713 = 6'h9 == stage1_index ? 1'h0 : lru_list_9; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_714 = 6'ha == stage1_index ? 1'h0 : lru_list_10; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_715 = 6'hb == stage1_index ? 1'h0 : lru_list_11; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_716 = 6'hc == stage1_index ? 1'h0 : lru_list_12; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_717 = 6'hd == stage1_index ? 1'h0 : lru_list_13; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_718 = 6'he == stage1_index ? 1'h0 : lru_list_14; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_719 = 6'hf == stage1_index ? 1'h0 : lru_list_15; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_720 = 6'h10 == stage1_index ? 1'h0 : lru_list_16; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_721 = 6'h11 == stage1_index ? 1'h0 : lru_list_17; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_722 = 6'h12 == stage1_index ? 1'h0 : lru_list_18; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_723 = 6'h13 == stage1_index ? 1'h0 : lru_list_19; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_724 = 6'h14 == stage1_index ? 1'h0 : lru_list_20; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_725 = 6'h15 == stage1_index ? 1'h0 : lru_list_21; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_726 = 6'h16 == stage1_index ? 1'h0 : lru_list_22; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_727 = 6'h17 == stage1_index ? 1'h0 : lru_list_23; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_728 = 6'h18 == stage1_index ? 1'h0 : lru_list_24; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_729 = 6'h19 == stage1_index ? 1'h0 : lru_list_25; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_730 = 6'h1a == stage1_index ? 1'h0 : lru_list_26; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_731 = 6'h1b == stage1_index ? 1'h0 : lru_list_27; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_732 = 6'h1c == stage1_index ? 1'h0 : lru_list_28; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_733 = 6'h1d == stage1_index ? 1'h0 : lru_list_29; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_734 = 6'h1e == stage1_index ? 1'h0 : lru_list_30; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_735 = 6'h1f == stage1_index ? 1'h0 : lru_list_31; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_736 = 6'h20 == stage1_index ? 1'h0 : lru_list_32; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_737 = 6'h21 == stage1_index ? 1'h0 : lru_list_33; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_738 = 6'h22 == stage1_index ? 1'h0 : lru_list_34; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_739 = 6'h23 == stage1_index ? 1'h0 : lru_list_35; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_740 = 6'h24 == stage1_index ? 1'h0 : lru_list_36; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_741 = 6'h25 == stage1_index ? 1'h0 : lru_list_37; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_742 = 6'h26 == stage1_index ? 1'h0 : lru_list_38; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_743 = 6'h27 == stage1_index ? 1'h0 : lru_list_39; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_744 = 6'h28 == stage1_index ? 1'h0 : lru_list_40; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_745 = 6'h29 == stage1_index ? 1'h0 : lru_list_41; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_746 = 6'h2a == stage1_index ? 1'h0 : lru_list_42; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_747 = 6'h2b == stage1_index ? 1'h0 : lru_list_43; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_748 = 6'h2c == stage1_index ? 1'h0 : lru_list_44; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_749 = 6'h2d == stage1_index ? 1'h0 : lru_list_45; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_750 = 6'h2e == stage1_index ? 1'h0 : lru_list_46; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_751 = 6'h2f == stage1_index ? 1'h0 : lru_list_47; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_752 = 6'h30 == stage1_index ? 1'h0 : lru_list_48; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_753 = 6'h31 == stage1_index ? 1'h0 : lru_list_49; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_754 = 6'h32 == stage1_index ? 1'h0 : lru_list_50; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_755 = 6'h33 == stage1_index ? 1'h0 : lru_list_51; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_756 = 6'h34 == stage1_index ? 1'h0 : lru_list_52; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_757 = 6'h35 == stage1_index ? 1'h0 : lru_list_53; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_758 = 6'h36 == stage1_index ? 1'h0 : lru_list_54; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_759 = 6'h37 == stage1_index ? 1'h0 : lru_list_55; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_760 = 6'h38 == stage1_index ? 1'h0 : lru_list_56; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_761 = 6'h39 == stage1_index ? 1'h0 : lru_list_57; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_762 = 6'h3a == stage1_index ? 1'h0 : lru_list_58; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_763 = 6'h3b == stage1_index ? 1'h0 : lru_list_59; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_764 = 6'h3c == stage1_index ? 1'h0 : lru_list_60; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_765 = 6'h3d == stage1_index ? 1'h0 : lru_list_61; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_766 = 6'h3e == stage1_index ? 1'h0 : lru_list_62; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_767 = 6'h3f == stage1_index ? 1'h0 : lru_list_63; // @[DCache.scala 278:32 DCache.scala 278:32 DCache.scala 118:35]
  wire  _GEN_768 = _GEN_3579 | valid_array_0_0; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_769 = _GEN_3580 | valid_array_0_1; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_770 = _GEN_3581 | valid_array_0_2; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_771 = _GEN_3582 | valid_array_0_3; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_772 = _GEN_3583 | valid_array_0_4; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_773 = _GEN_3584 | valid_array_0_5; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_774 = _GEN_3585 | valid_array_0_6; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_775 = _GEN_3586 | valid_array_0_7; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_776 = _GEN_3587 | valid_array_0_8; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_777 = _GEN_3588 | valid_array_0_9; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_778 = _GEN_3589 | valid_array_0_10; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_779 = _GEN_3590 | valid_array_0_11; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_780 = _GEN_3591 | valid_array_0_12; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_781 = _GEN_3592 | valid_array_0_13; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_782 = _GEN_3593 | valid_array_0_14; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_783 = _GEN_3594 | valid_array_0_15; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_784 = _GEN_3595 | valid_array_0_16; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_785 = _GEN_3596 | valid_array_0_17; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_786 = _GEN_3597 | valid_array_0_18; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_787 = _GEN_3598 | valid_array_0_19; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_788 = _GEN_3599 | valid_array_0_20; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_789 = _GEN_3600 | valid_array_0_21; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_790 = _GEN_3601 | valid_array_0_22; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_791 = _GEN_3602 | valid_array_0_23; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_792 = _GEN_3603 | valid_array_0_24; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_793 = _GEN_3604 | valid_array_0_25; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_794 = _GEN_3605 | valid_array_0_26; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_795 = _GEN_3606 | valid_array_0_27; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_796 = _GEN_3607 | valid_array_0_28; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_797 = _GEN_3608 | valid_array_0_29; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_798 = _GEN_3609 | valid_array_0_30; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_799 = _GEN_3610 | valid_array_0_31; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_800 = _GEN_3611 | valid_array_0_32; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_801 = _GEN_3612 | valid_array_0_33; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_802 = _GEN_3613 | valid_array_0_34; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_803 = _GEN_3614 | valid_array_0_35; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_804 = _GEN_3615 | valid_array_0_36; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_805 = _GEN_3616 | valid_array_0_37; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_806 = _GEN_3617 | valid_array_0_38; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_807 = _GEN_3618 | valid_array_0_39; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_808 = _GEN_3619 | valid_array_0_40; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_809 = _GEN_3620 | valid_array_0_41; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_810 = _GEN_3621 | valid_array_0_42; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_811 = _GEN_3622 | valid_array_0_43; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_812 = _GEN_3623 | valid_array_0_44; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_813 = _GEN_3624 | valid_array_0_45; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_814 = _GEN_3625 | valid_array_0_46; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_815 = _GEN_3626 | valid_array_0_47; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_816 = _GEN_3627 | valid_array_0_48; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_817 = _GEN_3628 | valid_array_0_49; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_818 = _GEN_3629 | valid_array_0_50; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_819 = _GEN_3630 | valid_array_0_51; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_820 = _GEN_3631 | valid_array_0_52; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_821 = _GEN_3632 | valid_array_0_53; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_822 = _GEN_3633 | valid_array_0_54; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_823 = _GEN_3634 | valid_array_0_55; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_824 = _GEN_3635 | valid_array_0_56; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_825 = _GEN_3636 | valid_array_0_57; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_826 = _GEN_3637 | valid_array_0_58; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_827 = _GEN_3638 | valid_array_0_59; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_828 = _GEN_3639 | valid_array_0_60; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_829 = _GEN_3640 | valid_array_0_61; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_830 = _GEN_3641 | valid_array_0_62; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_831 = _GEN_3642 | valid_array_0_63; // @[DCache.scala 282:37 DCache.scala 282:37 DCache.scala 115:44]
  wire  _GEN_832 = 6'h0 == stage1_index ? dirty_array_in : dirty_array_0_0; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_833 = 6'h1 == stage1_index ? dirty_array_in : dirty_array_0_1; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_834 = 6'h2 == stage1_index ? dirty_array_in : dirty_array_0_2; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_835 = 6'h3 == stage1_index ? dirty_array_in : dirty_array_0_3; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_836 = 6'h4 == stage1_index ? dirty_array_in : dirty_array_0_4; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_837 = 6'h5 == stage1_index ? dirty_array_in : dirty_array_0_5; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_838 = 6'h6 == stage1_index ? dirty_array_in : dirty_array_0_6; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_839 = 6'h7 == stage1_index ? dirty_array_in : dirty_array_0_7; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_840 = 6'h8 == stage1_index ? dirty_array_in : dirty_array_0_8; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_841 = 6'h9 == stage1_index ? dirty_array_in : dirty_array_0_9; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_842 = 6'ha == stage1_index ? dirty_array_in : dirty_array_0_10; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_843 = 6'hb == stage1_index ? dirty_array_in : dirty_array_0_11; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_844 = 6'hc == stage1_index ? dirty_array_in : dirty_array_0_12; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_845 = 6'hd == stage1_index ? dirty_array_in : dirty_array_0_13; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_846 = 6'he == stage1_index ? dirty_array_in : dirty_array_0_14; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_847 = 6'hf == stage1_index ? dirty_array_in : dirty_array_0_15; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_848 = 6'h10 == stage1_index ? dirty_array_in : dirty_array_0_16; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_849 = 6'h11 == stage1_index ? dirty_array_in : dirty_array_0_17; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_850 = 6'h12 == stage1_index ? dirty_array_in : dirty_array_0_18; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_851 = 6'h13 == stage1_index ? dirty_array_in : dirty_array_0_19; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_852 = 6'h14 == stage1_index ? dirty_array_in : dirty_array_0_20; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_853 = 6'h15 == stage1_index ? dirty_array_in : dirty_array_0_21; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_854 = 6'h16 == stage1_index ? dirty_array_in : dirty_array_0_22; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_855 = 6'h17 == stage1_index ? dirty_array_in : dirty_array_0_23; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_856 = 6'h18 == stage1_index ? dirty_array_in : dirty_array_0_24; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_857 = 6'h19 == stage1_index ? dirty_array_in : dirty_array_0_25; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_858 = 6'h1a == stage1_index ? dirty_array_in : dirty_array_0_26; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_859 = 6'h1b == stage1_index ? dirty_array_in : dirty_array_0_27; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_860 = 6'h1c == stage1_index ? dirty_array_in : dirty_array_0_28; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_861 = 6'h1d == stage1_index ? dirty_array_in : dirty_array_0_29; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_862 = 6'h1e == stage1_index ? dirty_array_in : dirty_array_0_30; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_863 = 6'h1f == stage1_index ? dirty_array_in : dirty_array_0_31; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_864 = 6'h20 == stage1_index ? dirty_array_in : dirty_array_0_32; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_865 = 6'h21 == stage1_index ? dirty_array_in : dirty_array_0_33; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_866 = 6'h22 == stage1_index ? dirty_array_in : dirty_array_0_34; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_867 = 6'h23 == stage1_index ? dirty_array_in : dirty_array_0_35; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_868 = 6'h24 == stage1_index ? dirty_array_in : dirty_array_0_36; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_869 = 6'h25 == stage1_index ? dirty_array_in : dirty_array_0_37; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_870 = 6'h26 == stage1_index ? dirty_array_in : dirty_array_0_38; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_871 = 6'h27 == stage1_index ? dirty_array_in : dirty_array_0_39; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_872 = 6'h28 == stage1_index ? dirty_array_in : dirty_array_0_40; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_873 = 6'h29 == stage1_index ? dirty_array_in : dirty_array_0_41; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_874 = 6'h2a == stage1_index ? dirty_array_in : dirty_array_0_42; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_875 = 6'h2b == stage1_index ? dirty_array_in : dirty_array_0_43; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_876 = 6'h2c == stage1_index ? dirty_array_in : dirty_array_0_44; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_877 = 6'h2d == stage1_index ? dirty_array_in : dirty_array_0_45; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_878 = 6'h2e == stage1_index ? dirty_array_in : dirty_array_0_46; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_879 = 6'h2f == stage1_index ? dirty_array_in : dirty_array_0_47; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_880 = 6'h30 == stage1_index ? dirty_array_in : dirty_array_0_48; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_881 = 6'h31 == stage1_index ? dirty_array_in : dirty_array_0_49; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_882 = 6'h32 == stage1_index ? dirty_array_in : dirty_array_0_50; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_883 = 6'h33 == stage1_index ? dirty_array_in : dirty_array_0_51; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_884 = 6'h34 == stage1_index ? dirty_array_in : dirty_array_0_52; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_885 = 6'h35 == stage1_index ? dirty_array_in : dirty_array_0_53; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_886 = 6'h36 == stage1_index ? dirty_array_in : dirty_array_0_54; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_887 = 6'h37 == stage1_index ? dirty_array_in : dirty_array_0_55; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_888 = 6'h38 == stage1_index ? dirty_array_in : dirty_array_0_56; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_889 = 6'h39 == stage1_index ? dirty_array_in : dirty_array_0_57; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_890 = 6'h3a == stage1_index ? dirty_array_in : dirty_array_0_58; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_891 = 6'h3b == stage1_index ? dirty_array_in : dirty_array_0_59; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_892 = 6'h3c == stage1_index ? dirty_array_in : dirty_array_0_60; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_893 = 6'h3d == stage1_index ? dirty_array_in : dirty_array_0_61; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_894 = 6'h3e == stage1_index ? dirty_array_in : dirty_array_0_62; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_895 = 6'h3f == stage1_index ? dirty_array_in : dirty_array_0_63; // @[DCache.scala 283:37 DCache.scala 283:37 DCache.scala 113:44]
  wire  _GEN_961 = next_way ? 1'h0 : 1'h1; // @[DCache.scala 270:19 CacheBase.scala 72:13 CacheBase.scala 81:13]
  wire  _array_rd_index_T_1 = hit_reg_x8 & io_prev_bits_flush; // @[DCache.scala 453:29]
  wire [5:0] _array_rd_index_T_6 = flush_index + 6'h1; // @[DCache.scala 454:74]
  wire  _array_rd_index_T_13 = _T_10 | _T | _T_18 | _T_13; // @[DCache.scala 455:77]
  wire [5:0] _array_rd_index_T_17 = flush_cnt_rst ? prev_index : stage1_index; // @[Mux.scala 98:16]
  wire [5:0] _array_rd_index_T_18 = go_on ? prev_index : _array_rd_index_T_17; // @[Mux.scala 98:16]
  wire [5:0] _array_rd_index_T_19 = _T_19 ? stage1_index : _array_rd_index_T_18; // @[Mux.scala 98:16]
  wire [5:0] _array_rd_index_T_20 = _array_rd_index_T_13 ? flush_index : _array_rd_index_T_19; // @[Mux.scala 98:16]
  wire [5:0] _array_rd_index_T_21 = flush_cnt_en ? _array_rd_index_T_6 : _array_rd_index_T_20; // @[Mux.scala 98:16]
  wire [5:0] array_rd_index = _array_rd_index_T_1 ? flush_index : _array_rd_index_T_21; // @[Mux.scala 98:16]
  wire [5:0] _GEN_962 = next_way ? stage1_index : array_rd_index; // @[DCache.scala 270:19 CacheBase.scala 73:14 CacheBase.scala 82:14]
  wire  _is_save = _T_19 | hit_reg_x8; // @[DCache.scala 431:59]
  wire [127:0] save_data_src = _is_save ? cache_line_data_out : maxi4_manager_io_out_data; // @[DCache.scala 432:41]
  wire [4:0] save_data_size_2 = {1'h0,stage1_out_bits_size_dword,stage1_out_bits_size_word,stage1_out_bits_size_hword,
    stage1_out_bits_size_byte}; // @[Cat.scala 30:58]
  wire [4:0] _GEN_3771 = {{1'd0}, addr_array_0_lo}; // @[DCache.scala 444:65]
  wire [4:0] _save_start_bit_rshift_T_1 = _GEN_3771 + save_data_size_2; // @[DCache.scala 444:65]
  wire [7:0] save_start_bit_rshift = {_save_start_bit_rshift_T_1, 3'h0}; // @[DCache.scala 444:84]
  wire [127:0] save_data_inserted_H1 = save_data_src >> save_start_bit_rshift; // @[Util.scala 15:19]
  wire [382:0] _GEN_3772 = {{255'd0}, save_data_inserted_H1}; // @[Util.scala 16:17]
  wire [382:0] _save_data_inserted_H_T = _GEN_3772 << save_start_bit_rshift; // @[Util.scala 16:17]
  wire [127:0] save_data_inserted_H = _save_data_inserted_H_T[127:0]; // @[Util.scala 16:36 Util.scala 16:36]
  wire [63:0] _save_data_token_T_5 = stage1_out_bits_size_word ? {{32'd0}, stage1_out_bits_data_ex2mem_we_data[31:0]} :
    stage1_out_bits_data_ex2mem_we_data; // @[Mux.scala 98:16]
  wire [63:0] _save_data_token_T_6 = stage1_out_bits_size_hword ? {{48'd0}, stage1_out_bits_data_ex2mem_we_data[15:0]}
     : _save_data_token_T_5; // @[Mux.scala 98:16]
  wire [63:0] save_data_token = stage1_out_bits_size_byte ? {{56'd0}, stage1_out_bits_data_ex2mem_we_data[7:0]} :
    _save_data_token_T_6; // @[Mux.scala 98:16]
  wire [6:0] save_start_bit_lshift2 = {addr_array_0_lo, 3'h0}; // @[DCache.scala 446:64]
  wire [190:0] _GEN_3773 = {{127'd0}, save_data_token}; // @[Util.scala 19:20]
  wire [190:0] _save_data_inserted_M_T = _GEN_3773 << save_start_bit_lshift2; // @[Util.scala 19:20]
  wire [127:0] save_data_inserted_M = _save_data_inserted_M_T[127:0]; // @[Util.scala 19:40 Util.scala 19:40]
  wire [127:0] _save_data_inserted_T = save_data_inserted_H | save_data_inserted_M; // @[Util.scala 22:7]
  wire [7:0] _GEN_3774 = {{1'd0}, save_start_bit_lshift2}; // @[DCache.scala 445:45]
  wire [7:0] save_start_bit_lshift = 8'h80 - _GEN_3774; // @[DCache.scala 445:45]
  wire [382:0] _GEN_3775 = {{255'd0}, save_data_src}; // @[Util.scala 17:19]
  wire [382:0] _save_data_inserted_L1_T = _GEN_3775 << save_start_bit_lshift; // @[Util.scala 17:19]
  wire [127:0] save_data_inserted_L1 = _save_data_inserted_L1_T[127:0]; // @[Util.scala 17:38 Util.scala 17:38]
  wire [127:0] save_data_inserted_L = save_data_inserted_L1 >> save_start_bit_lshift; // @[Util.scala 18:17]
  wire [127:0] save_data_inserted = _save_data_inserted_T | save_data_inserted_L; // @[Util.scala 22:11]
  wire [127:0] save_data = stage1_out_bits_data_id2mem_memory_we_en ? save_data_inserted : maxi4_manager_io_out_data; // @[DCache.scala 448:19]
  wire [127:0] _GEN_963 = next_way ? save_data : 128'h0; // @[DCache.scala 270:19 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire [127:0] _GEN_964 = next_way ? 128'h0 : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 270:19 CacheBase.scala 75:15 CacheBase.scala 84:15]
  wire [127:0] _GEN_966 = next_way ? x12 : 128'h0; // @[DCache.scala 270:19 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire [5:0] _GEN_1097 = next_way ? array_rd_index : stage1_index; // @[DCache.scala 270:19 CacheBase.scala 82:14 CacheBase.scala 73:14]
  wire [127:0] _GEN_1098 = next_way ? 128'h0 : save_data; // @[DCache.scala 270:19 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire [127:0] _GEN_1099 = next_way ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[DCache.scala 270:19 CacheBase.scala 84:15 CacheBase.scala 75:15]
  wire [127:0] _GEN_1101 = next_way ? 128'h0 : x12; // @[DCache.scala 270:19 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire  _GEN_1231 = 6'h0 == flush_index | lru_list_0; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1232 = 6'h1 == flush_index | lru_list_1; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1233 = 6'h2 == flush_index | lru_list_2; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1234 = 6'h3 == flush_index | lru_list_3; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1235 = 6'h4 == flush_index | lru_list_4; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1236 = 6'h5 == flush_index | lru_list_5; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1237 = 6'h6 == flush_index | lru_list_6; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1238 = 6'h7 == flush_index | lru_list_7; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1239 = 6'h8 == flush_index | lru_list_8; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1240 = 6'h9 == flush_index | lru_list_9; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1241 = 6'ha == flush_index | lru_list_10; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1242 = 6'hb == flush_index | lru_list_11; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1243 = 6'hc == flush_index | lru_list_12; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1244 = 6'hd == flush_index | lru_list_13; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1245 = 6'he == flush_index | lru_list_14; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1246 = 6'hf == flush_index | lru_list_15; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1247 = 6'h10 == flush_index | lru_list_16; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1248 = 6'h11 == flush_index | lru_list_17; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1249 = 6'h12 == flush_index | lru_list_18; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1250 = 6'h13 == flush_index | lru_list_19; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1251 = 6'h14 == flush_index | lru_list_20; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1252 = 6'h15 == flush_index | lru_list_21; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1253 = 6'h16 == flush_index | lru_list_22; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1254 = 6'h17 == flush_index | lru_list_23; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1255 = 6'h18 == flush_index | lru_list_24; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1256 = 6'h19 == flush_index | lru_list_25; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1257 = 6'h1a == flush_index | lru_list_26; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1258 = 6'h1b == flush_index | lru_list_27; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1259 = 6'h1c == flush_index | lru_list_28; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1260 = 6'h1d == flush_index | lru_list_29; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1261 = 6'h1e == flush_index | lru_list_30; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1262 = 6'h1f == flush_index | lru_list_31; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1263 = 6'h20 == flush_index | lru_list_32; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1264 = 6'h21 == flush_index | lru_list_33; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1265 = 6'h22 == flush_index | lru_list_34; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1266 = 6'h23 == flush_index | lru_list_35; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1267 = 6'h24 == flush_index | lru_list_36; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1268 = 6'h25 == flush_index | lru_list_37; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1269 = 6'h26 == flush_index | lru_list_38; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1270 = 6'h27 == flush_index | lru_list_39; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1271 = 6'h28 == flush_index | lru_list_40; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1272 = 6'h29 == flush_index | lru_list_41; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1273 = 6'h2a == flush_index | lru_list_42; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1274 = 6'h2b == flush_index | lru_list_43; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1275 = 6'h2c == flush_index | lru_list_44; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1276 = 6'h2d == flush_index | lru_list_45; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1277 = 6'h2e == flush_index | lru_list_46; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1278 = 6'h2f == flush_index | lru_list_47; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1279 = 6'h30 == flush_index | lru_list_48; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1280 = 6'h31 == flush_index | lru_list_49; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1281 = 6'h32 == flush_index | lru_list_50; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1282 = 6'h33 == flush_index | lru_list_51; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1283 = 6'h34 == flush_index | lru_list_52; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1284 = 6'h35 == flush_index | lru_list_53; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1285 = 6'h36 == flush_index | lru_list_54; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1286 = 6'h37 == flush_index | lru_list_55; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1287 = 6'h38 == flush_index | lru_list_56; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1288 = 6'h39 == flush_index | lru_list_57; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1289 = 6'h3a == flush_index | lru_list_58; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1290 = 6'h3b == flush_index | lru_list_59; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1291 = 6'h3c == flush_index | lru_list_60; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1292 = 6'h3d == flush_index | lru_list_61; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1293 = 6'h3e == flush_index | lru_list_62; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1294 = 6'h3f == flush_index | lru_list_63; // @[DCache.scala 288:31 DCache.scala 288:31 DCache.scala 118:35]
  wire  _GEN_1424 = flush_way ? 1'h0 : 1'h1; // @[DCache.scala 287:22 CacheBase.scala 72:13 CacheBase.scala 81:13]
  wire [5:0] _GEN_1425 = flush_way ? flush_index : array_rd_index; // @[DCache.scala 287:22 CacheBase.scala 73:14 CacheBase.scala 82:14]
  wire [127:0] _GEN_1426 = flush_way ? 128'h0 : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 287:22 CacheBase.scala 75:15 CacheBase.scala 84:15]
  wire [5:0] _GEN_1430 = flush_way ? array_rd_index : flush_index; // @[DCache.scala 287:22 CacheBase.scala 82:14 CacheBase.scala 73:14]
  wire [127:0] _GEN_1431 = flush_way ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[DCache.scala 287:22 CacheBase.scala 84:15 CacheBase.scala 75:15]
  wire  _GEN_1626 = 6'h0 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_0; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1627 = 6'h1 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_1; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1628 = 6'h2 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_2; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1629 = 6'h3 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_3; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1630 = 6'h4 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_4; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1631 = 6'h5 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_5; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1632 = 6'h6 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_6; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1633 = 6'h7 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_7; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1634 = 6'h8 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_8; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1635 = 6'h9 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_9; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1636 = 6'ha == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_10; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1637 = 6'hb == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_11; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1638 = 6'hc == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_12; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1639 = 6'hd == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_13; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1640 = 6'he == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_14; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1641 = 6'hf == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_15; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1642 = 6'h10 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_16; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1643 = 6'h11 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_17; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1644 = 6'h12 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_18; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1645 = 6'h13 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_19; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1646 = 6'h14 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_20; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1647 = 6'h15 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_21; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1648 = 6'h16 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_22; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1649 = 6'h17 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_23; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1650 = 6'h18 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_24; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1651 = 6'h19 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_25; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1652 = 6'h1a == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_26; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1653 = 6'h1b == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_27; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1654 = 6'h1c == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_28; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1655 = 6'h1d == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_29; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1656 = 6'h1e == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_30; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1657 = 6'h1f == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_31; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1658 = 6'h20 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_32; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1659 = 6'h21 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_33; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1660 = 6'h22 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_34; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1661 = 6'h23 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_35; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1662 = 6'h24 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_36; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1663 = 6'h25 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_37; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1664 = 6'h26 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_38; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1665 = 6'h27 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_39; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1666 = 6'h28 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_40; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1667 = 6'h29 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_41; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1668 = 6'h2a == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_42; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1669 = 6'h2b == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_43; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1670 = 6'h2c == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_44; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1671 = 6'h2d == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_45; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1672 = 6'h2e == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_46; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1673 = 6'h2f == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_47; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1674 = 6'h30 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_48; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1675 = 6'h31 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_49; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1676 = 6'h32 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_50; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1677 = 6'h33 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_51; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1678 = 6'h34 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_52; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1679 = 6'h35 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_53; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1680 = 6'h36 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_54; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1681 = 6'h37 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_55; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1682 = 6'h38 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_56; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1683 = 6'h39 == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_57; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1684 = 6'h3a == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_58; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1685 = 6'h3b == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_59; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1686 = 6'h3c == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_60; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1687 = 6'h3d == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_61; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1688 = 6'h3e == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_62; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1689 = 6'h3f == stage1_index ? dirty_array_in | _GEN_485 : dirty_array_0_63; // @[DCache.scala 304:39 DCache.scala 304:39 DCache.scala 113:44]
  wire  _GEN_1882 = 6'h0 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_0; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1883 = 6'h1 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_1; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1884 = 6'h2 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_2; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1885 = 6'h3 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_3; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1886 = 6'h4 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_4; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1887 = 6'h5 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_5; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1888 = 6'h6 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_6; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1889 = 6'h7 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_7; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1890 = 6'h8 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_8; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1891 = 6'h9 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_9; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1892 = 6'ha == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_10; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1893 = 6'hb == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_11; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1894 = 6'hc == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_12; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1895 = 6'hd == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_13; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1896 = 6'he == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_14; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1897 = 6'hf == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_15; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1898 = 6'h10 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_16; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1899 = 6'h11 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_17; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1900 = 6'h12 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_18; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1901 = 6'h13 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_19; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1902 = 6'h14 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_20; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1903 = 6'h15 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_21; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1904 = 6'h16 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_22; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1905 = 6'h17 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_23; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1906 = 6'h18 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_24; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1907 = 6'h19 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_25; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1908 = 6'h1a == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_26; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1909 = 6'h1b == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_27; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1910 = 6'h1c == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_28; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1911 = 6'h1d == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_29; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1912 = 6'h1e == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_30; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1913 = 6'h1f == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_31; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1914 = 6'h20 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_32; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1915 = 6'h21 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_33; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1916 = 6'h22 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_34; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1917 = 6'h23 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_35; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1918 = 6'h24 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_36; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1919 = 6'h25 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_37; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1920 = 6'h26 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_38; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1921 = 6'h27 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_39; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1922 = 6'h28 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_40; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1923 = 6'h29 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_41; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1924 = 6'h2a == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_42; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1925 = 6'h2b == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_43; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1926 = 6'h2c == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_44; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1927 = 6'h2d == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_45; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1928 = 6'h2e == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_46; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1929 = 6'h2f == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_47; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1930 = 6'h30 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_48; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1931 = 6'h31 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_49; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1932 = 6'h32 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_50; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1933 = 6'h33 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_51; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1934 = 6'h34 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_52; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1935 = 6'h35 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_53; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1936 = 6'h36 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_54; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1937 = 6'h37 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_55; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1938 = 6'h38 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_56; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1939 = 6'h39 == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_57; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1940 = 6'h3a == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_58; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1941 = 6'h3b == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_59; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1942 = 6'h3c == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_60; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1943 = 6'h3d == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_61; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1944 = 6'h3e == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_62; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1945 = 6'h3f == stage1_index ? dirty_array_in | _GEN_421 : dirty_array_1_63; // @[DCache.scala 311:39 DCache.scala 311:39 DCache.scala 114:44]
  wire  _GEN_1946 = ~hit_reg ? _GEN_704 : _GEN_512; // @[DCache.scala 298:28]
  wire  _GEN_1947 = ~hit_reg ? _GEN_705 : _GEN_513; // @[DCache.scala 298:28]
  wire  _GEN_1948 = ~hit_reg ? _GEN_706 : _GEN_514; // @[DCache.scala 298:28]
  wire  _GEN_1949 = ~hit_reg ? _GEN_707 : _GEN_515; // @[DCache.scala 298:28]
  wire  _GEN_1950 = ~hit_reg ? _GEN_708 : _GEN_516; // @[DCache.scala 298:28]
  wire  _GEN_1951 = ~hit_reg ? _GEN_709 : _GEN_517; // @[DCache.scala 298:28]
  wire  _GEN_1952 = ~hit_reg ? _GEN_710 : _GEN_518; // @[DCache.scala 298:28]
  wire  _GEN_1953 = ~hit_reg ? _GEN_711 : _GEN_519; // @[DCache.scala 298:28]
  wire  _GEN_1954 = ~hit_reg ? _GEN_712 : _GEN_520; // @[DCache.scala 298:28]
  wire  _GEN_1955 = ~hit_reg ? _GEN_713 : _GEN_521; // @[DCache.scala 298:28]
  wire  _GEN_1956 = ~hit_reg ? _GEN_714 : _GEN_522; // @[DCache.scala 298:28]
  wire  _GEN_1957 = ~hit_reg ? _GEN_715 : _GEN_523; // @[DCache.scala 298:28]
  wire  _GEN_1958 = ~hit_reg ? _GEN_716 : _GEN_524; // @[DCache.scala 298:28]
  wire  _GEN_1959 = ~hit_reg ? _GEN_717 : _GEN_525; // @[DCache.scala 298:28]
  wire  _GEN_1960 = ~hit_reg ? _GEN_718 : _GEN_526; // @[DCache.scala 298:28]
  wire  _GEN_1961 = ~hit_reg ? _GEN_719 : _GEN_527; // @[DCache.scala 298:28]
  wire  _GEN_1962 = ~hit_reg ? _GEN_720 : _GEN_528; // @[DCache.scala 298:28]
  wire  _GEN_1963 = ~hit_reg ? _GEN_721 : _GEN_529; // @[DCache.scala 298:28]
  wire  _GEN_1964 = ~hit_reg ? _GEN_722 : _GEN_530; // @[DCache.scala 298:28]
  wire  _GEN_1965 = ~hit_reg ? _GEN_723 : _GEN_531; // @[DCache.scala 298:28]
  wire  _GEN_1966 = ~hit_reg ? _GEN_724 : _GEN_532; // @[DCache.scala 298:28]
  wire  _GEN_1967 = ~hit_reg ? _GEN_725 : _GEN_533; // @[DCache.scala 298:28]
  wire  _GEN_1968 = ~hit_reg ? _GEN_726 : _GEN_534; // @[DCache.scala 298:28]
  wire  _GEN_1969 = ~hit_reg ? _GEN_727 : _GEN_535; // @[DCache.scala 298:28]
  wire  _GEN_1970 = ~hit_reg ? _GEN_728 : _GEN_536; // @[DCache.scala 298:28]
  wire  _GEN_1971 = ~hit_reg ? _GEN_729 : _GEN_537; // @[DCache.scala 298:28]
  wire  _GEN_1972 = ~hit_reg ? _GEN_730 : _GEN_538; // @[DCache.scala 298:28]
  wire  _GEN_1973 = ~hit_reg ? _GEN_731 : _GEN_539; // @[DCache.scala 298:28]
  wire  _GEN_1974 = ~hit_reg ? _GEN_732 : _GEN_540; // @[DCache.scala 298:28]
  wire  _GEN_1975 = ~hit_reg ? _GEN_733 : _GEN_541; // @[DCache.scala 298:28]
  wire  _GEN_1976 = ~hit_reg ? _GEN_734 : _GEN_542; // @[DCache.scala 298:28]
  wire  _GEN_1977 = ~hit_reg ? _GEN_735 : _GEN_543; // @[DCache.scala 298:28]
  wire  _GEN_1978 = ~hit_reg ? _GEN_736 : _GEN_544; // @[DCache.scala 298:28]
  wire  _GEN_1979 = ~hit_reg ? _GEN_737 : _GEN_545; // @[DCache.scala 298:28]
  wire  _GEN_1980 = ~hit_reg ? _GEN_738 : _GEN_546; // @[DCache.scala 298:28]
  wire  _GEN_1981 = ~hit_reg ? _GEN_739 : _GEN_547; // @[DCache.scala 298:28]
  wire  _GEN_1982 = ~hit_reg ? _GEN_740 : _GEN_548; // @[DCache.scala 298:28]
  wire  _GEN_1983 = ~hit_reg ? _GEN_741 : _GEN_549; // @[DCache.scala 298:28]
  wire  _GEN_1984 = ~hit_reg ? _GEN_742 : _GEN_550; // @[DCache.scala 298:28]
  wire  _GEN_1985 = ~hit_reg ? _GEN_743 : _GEN_551; // @[DCache.scala 298:28]
  wire  _GEN_1986 = ~hit_reg ? _GEN_744 : _GEN_552; // @[DCache.scala 298:28]
  wire  _GEN_1987 = ~hit_reg ? _GEN_745 : _GEN_553; // @[DCache.scala 298:28]
  wire  _GEN_1988 = ~hit_reg ? _GEN_746 : _GEN_554; // @[DCache.scala 298:28]
  wire  _GEN_1989 = ~hit_reg ? _GEN_747 : _GEN_555; // @[DCache.scala 298:28]
  wire  _GEN_1990 = ~hit_reg ? _GEN_748 : _GEN_556; // @[DCache.scala 298:28]
  wire  _GEN_1991 = ~hit_reg ? _GEN_749 : _GEN_557; // @[DCache.scala 298:28]
  wire  _GEN_1992 = ~hit_reg ? _GEN_750 : _GEN_558; // @[DCache.scala 298:28]
  wire  _GEN_1993 = ~hit_reg ? _GEN_751 : _GEN_559; // @[DCache.scala 298:28]
  wire  _GEN_1994 = ~hit_reg ? _GEN_752 : _GEN_560; // @[DCache.scala 298:28]
  wire  _GEN_1995 = ~hit_reg ? _GEN_753 : _GEN_561; // @[DCache.scala 298:28]
  wire  _GEN_1996 = ~hit_reg ? _GEN_754 : _GEN_562; // @[DCache.scala 298:28]
  wire  _GEN_1997 = ~hit_reg ? _GEN_755 : _GEN_563; // @[DCache.scala 298:28]
  wire  _GEN_1998 = ~hit_reg ? _GEN_756 : _GEN_564; // @[DCache.scala 298:28]
  wire  _GEN_1999 = ~hit_reg ? _GEN_757 : _GEN_565; // @[DCache.scala 298:28]
  wire  _GEN_2000 = ~hit_reg ? _GEN_758 : _GEN_566; // @[DCache.scala 298:28]
  wire  _GEN_2001 = ~hit_reg ? _GEN_759 : _GEN_567; // @[DCache.scala 298:28]
  wire  _GEN_2002 = ~hit_reg ? _GEN_760 : _GEN_568; // @[DCache.scala 298:28]
  wire  _GEN_2003 = ~hit_reg ? _GEN_761 : _GEN_569; // @[DCache.scala 298:28]
  wire  _GEN_2004 = ~hit_reg ? _GEN_762 : _GEN_570; // @[DCache.scala 298:28]
  wire  _GEN_2005 = ~hit_reg ? _GEN_763 : _GEN_571; // @[DCache.scala 298:28]
  wire  _GEN_2006 = ~hit_reg ? _GEN_764 : _GEN_572; // @[DCache.scala 298:28]
  wire  _GEN_2007 = ~hit_reg ? _GEN_765 : _GEN_573; // @[DCache.scala 298:28]
  wire  _GEN_2008 = ~hit_reg ? _GEN_766 : _GEN_574; // @[DCache.scala 298:28]
  wire  _GEN_2009 = ~hit_reg ? _GEN_767 : _GEN_575; // @[DCache.scala 298:28]
  wire  _GEN_2011 = ~hit_reg ? 1'h0 : 1'h1; // @[DCache.scala 298:28 CacheBase.scala 72:13 CacheBase.scala 81:13]
  wire [5:0] _GEN_2012 = ~hit_reg ? stage1_index : array_rd_index; // @[DCache.scala 298:28 CacheBase.scala 73:14 CacheBase.scala 82:14]
  wire [127:0] _GEN_2013 = ~hit_reg ? save_data : 128'h0; // @[DCache.scala 298:28 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire [127:0] _GEN_2014 = ~hit_reg ? 128'h0 : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 298:28 CacheBase.scala 75:15 CacheBase.scala 84:15]
  wire [127:0] _GEN_2016 = ~hit_reg ? x12 : 128'h0; // @[DCache.scala 298:28 CacheBase.scala 74:15 CacheBase.scala 83:15]
  wire  _GEN_2018 = ~hit_reg ? _GEN_768 : valid_array_0_0; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2019 = ~hit_reg ? _GEN_769 : valid_array_0_1; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2020 = ~hit_reg ? _GEN_770 : valid_array_0_2; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2021 = ~hit_reg ? _GEN_771 : valid_array_0_3; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2022 = ~hit_reg ? _GEN_772 : valid_array_0_4; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2023 = ~hit_reg ? _GEN_773 : valid_array_0_5; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2024 = ~hit_reg ? _GEN_774 : valid_array_0_6; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2025 = ~hit_reg ? _GEN_775 : valid_array_0_7; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2026 = ~hit_reg ? _GEN_776 : valid_array_0_8; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2027 = ~hit_reg ? _GEN_777 : valid_array_0_9; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2028 = ~hit_reg ? _GEN_778 : valid_array_0_10; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2029 = ~hit_reg ? _GEN_779 : valid_array_0_11; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2030 = ~hit_reg ? _GEN_780 : valid_array_0_12; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2031 = ~hit_reg ? _GEN_781 : valid_array_0_13; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2032 = ~hit_reg ? _GEN_782 : valid_array_0_14; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2033 = ~hit_reg ? _GEN_783 : valid_array_0_15; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2034 = ~hit_reg ? _GEN_784 : valid_array_0_16; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2035 = ~hit_reg ? _GEN_785 : valid_array_0_17; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2036 = ~hit_reg ? _GEN_786 : valid_array_0_18; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2037 = ~hit_reg ? _GEN_787 : valid_array_0_19; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2038 = ~hit_reg ? _GEN_788 : valid_array_0_20; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2039 = ~hit_reg ? _GEN_789 : valid_array_0_21; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2040 = ~hit_reg ? _GEN_790 : valid_array_0_22; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2041 = ~hit_reg ? _GEN_791 : valid_array_0_23; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2042 = ~hit_reg ? _GEN_792 : valid_array_0_24; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2043 = ~hit_reg ? _GEN_793 : valid_array_0_25; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2044 = ~hit_reg ? _GEN_794 : valid_array_0_26; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2045 = ~hit_reg ? _GEN_795 : valid_array_0_27; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2046 = ~hit_reg ? _GEN_796 : valid_array_0_28; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2047 = ~hit_reg ? _GEN_797 : valid_array_0_29; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2048 = ~hit_reg ? _GEN_798 : valid_array_0_30; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2049 = ~hit_reg ? _GEN_799 : valid_array_0_31; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2050 = ~hit_reg ? _GEN_800 : valid_array_0_32; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2051 = ~hit_reg ? _GEN_801 : valid_array_0_33; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2052 = ~hit_reg ? _GEN_802 : valid_array_0_34; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2053 = ~hit_reg ? _GEN_803 : valid_array_0_35; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2054 = ~hit_reg ? _GEN_804 : valid_array_0_36; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2055 = ~hit_reg ? _GEN_805 : valid_array_0_37; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2056 = ~hit_reg ? _GEN_806 : valid_array_0_38; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2057 = ~hit_reg ? _GEN_807 : valid_array_0_39; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2058 = ~hit_reg ? _GEN_808 : valid_array_0_40; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2059 = ~hit_reg ? _GEN_809 : valid_array_0_41; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2060 = ~hit_reg ? _GEN_810 : valid_array_0_42; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2061 = ~hit_reg ? _GEN_811 : valid_array_0_43; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2062 = ~hit_reg ? _GEN_812 : valid_array_0_44; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2063 = ~hit_reg ? _GEN_813 : valid_array_0_45; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2064 = ~hit_reg ? _GEN_814 : valid_array_0_46; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2065 = ~hit_reg ? _GEN_815 : valid_array_0_47; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2066 = ~hit_reg ? _GEN_816 : valid_array_0_48; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2067 = ~hit_reg ? _GEN_817 : valid_array_0_49; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2068 = ~hit_reg ? _GEN_818 : valid_array_0_50; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2069 = ~hit_reg ? _GEN_819 : valid_array_0_51; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2070 = ~hit_reg ? _GEN_820 : valid_array_0_52; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2071 = ~hit_reg ? _GEN_821 : valid_array_0_53; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2072 = ~hit_reg ? _GEN_822 : valid_array_0_54; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2073 = ~hit_reg ? _GEN_823 : valid_array_0_55; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2074 = ~hit_reg ? _GEN_824 : valid_array_0_56; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2075 = ~hit_reg ? _GEN_825 : valid_array_0_57; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2076 = ~hit_reg ? _GEN_826 : valid_array_0_58; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2077 = ~hit_reg ? _GEN_827 : valid_array_0_59; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2078 = ~hit_reg ? _GEN_828 : valid_array_0_60; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2079 = ~hit_reg ? _GEN_829 : valid_array_0_61; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2080 = ~hit_reg ? _GEN_830 : valid_array_0_62; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2081 = ~hit_reg ? _GEN_831 : valid_array_0_63; // @[DCache.scala 298:28 DCache.scala 115:44]
  wire  _GEN_2082 = ~hit_reg ? _GEN_1626 : dirty_array_0_0; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2083 = ~hit_reg ? _GEN_1627 : dirty_array_0_1; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2084 = ~hit_reg ? _GEN_1628 : dirty_array_0_2; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2085 = ~hit_reg ? _GEN_1629 : dirty_array_0_3; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2086 = ~hit_reg ? _GEN_1630 : dirty_array_0_4; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2087 = ~hit_reg ? _GEN_1631 : dirty_array_0_5; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2088 = ~hit_reg ? _GEN_1632 : dirty_array_0_6; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2089 = ~hit_reg ? _GEN_1633 : dirty_array_0_7; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2090 = ~hit_reg ? _GEN_1634 : dirty_array_0_8; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2091 = ~hit_reg ? _GEN_1635 : dirty_array_0_9; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2092 = ~hit_reg ? _GEN_1636 : dirty_array_0_10; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2093 = ~hit_reg ? _GEN_1637 : dirty_array_0_11; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2094 = ~hit_reg ? _GEN_1638 : dirty_array_0_12; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2095 = ~hit_reg ? _GEN_1639 : dirty_array_0_13; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2096 = ~hit_reg ? _GEN_1640 : dirty_array_0_14; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2097 = ~hit_reg ? _GEN_1641 : dirty_array_0_15; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2098 = ~hit_reg ? _GEN_1642 : dirty_array_0_16; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2099 = ~hit_reg ? _GEN_1643 : dirty_array_0_17; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2100 = ~hit_reg ? _GEN_1644 : dirty_array_0_18; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2101 = ~hit_reg ? _GEN_1645 : dirty_array_0_19; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2102 = ~hit_reg ? _GEN_1646 : dirty_array_0_20; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2103 = ~hit_reg ? _GEN_1647 : dirty_array_0_21; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2104 = ~hit_reg ? _GEN_1648 : dirty_array_0_22; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2105 = ~hit_reg ? _GEN_1649 : dirty_array_0_23; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2106 = ~hit_reg ? _GEN_1650 : dirty_array_0_24; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2107 = ~hit_reg ? _GEN_1651 : dirty_array_0_25; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2108 = ~hit_reg ? _GEN_1652 : dirty_array_0_26; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2109 = ~hit_reg ? _GEN_1653 : dirty_array_0_27; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2110 = ~hit_reg ? _GEN_1654 : dirty_array_0_28; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2111 = ~hit_reg ? _GEN_1655 : dirty_array_0_29; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2112 = ~hit_reg ? _GEN_1656 : dirty_array_0_30; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2113 = ~hit_reg ? _GEN_1657 : dirty_array_0_31; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2114 = ~hit_reg ? _GEN_1658 : dirty_array_0_32; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2115 = ~hit_reg ? _GEN_1659 : dirty_array_0_33; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2116 = ~hit_reg ? _GEN_1660 : dirty_array_0_34; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2117 = ~hit_reg ? _GEN_1661 : dirty_array_0_35; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2118 = ~hit_reg ? _GEN_1662 : dirty_array_0_36; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2119 = ~hit_reg ? _GEN_1663 : dirty_array_0_37; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2120 = ~hit_reg ? _GEN_1664 : dirty_array_0_38; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2121 = ~hit_reg ? _GEN_1665 : dirty_array_0_39; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2122 = ~hit_reg ? _GEN_1666 : dirty_array_0_40; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2123 = ~hit_reg ? _GEN_1667 : dirty_array_0_41; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2124 = ~hit_reg ? _GEN_1668 : dirty_array_0_42; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2125 = ~hit_reg ? _GEN_1669 : dirty_array_0_43; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2126 = ~hit_reg ? _GEN_1670 : dirty_array_0_44; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2127 = ~hit_reg ? _GEN_1671 : dirty_array_0_45; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2128 = ~hit_reg ? _GEN_1672 : dirty_array_0_46; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2129 = ~hit_reg ? _GEN_1673 : dirty_array_0_47; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2130 = ~hit_reg ? _GEN_1674 : dirty_array_0_48; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2131 = ~hit_reg ? _GEN_1675 : dirty_array_0_49; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2132 = ~hit_reg ? _GEN_1676 : dirty_array_0_50; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2133 = ~hit_reg ? _GEN_1677 : dirty_array_0_51; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2134 = ~hit_reg ? _GEN_1678 : dirty_array_0_52; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2135 = ~hit_reg ? _GEN_1679 : dirty_array_0_53; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2136 = ~hit_reg ? _GEN_1680 : dirty_array_0_54; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2137 = ~hit_reg ? _GEN_1681 : dirty_array_0_55; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2138 = ~hit_reg ? _GEN_1682 : dirty_array_0_56; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2139 = ~hit_reg ? _GEN_1683 : dirty_array_0_57; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2140 = ~hit_reg ? _GEN_1684 : dirty_array_0_58; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2141 = ~hit_reg ? _GEN_1685 : dirty_array_0_59; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2142 = ~hit_reg ? _GEN_1686 : dirty_array_0_60; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2143 = ~hit_reg ? _GEN_1687 : dirty_array_0_61; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2144 = ~hit_reg ? _GEN_1688 : dirty_array_0_62; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire  _GEN_2145 = ~hit_reg ? _GEN_1689 : dirty_array_0_63; // @[DCache.scala 298:28 DCache.scala 113:44]
  wire [5:0] _GEN_2147 = ~hit_reg ? array_rd_index : stage1_index; // @[DCache.scala 298:28 CacheBase.scala 82:14 CacheBase.scala 73:14]
  wire [127:0] _GEN_2148 = ~hit_reg ? 128'h0 : save_data; // @[DCache.scala 298:28 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire [127:0] _GEN_2149 = ~hit_reg ? 128'hffffffffffffffffffffffffffffffff : 128'h0; // @[DCache.scala 298:28 CacheBase.scala 84:15 CacheBase.scala 75:15]
  wire [127:0] _GEN_2151 = ~hit_reg ? 128'h0 : x12; // @[DCache.scala 298:28 CacheBase.scala 83:15 CacheBase.scala 74:15]
  wire  _GEN_2153 = ~hit_reg ? valid_array_1_0 : _GEN_576; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2154 = ~hit_reg ? valid_array_1_1 : _GEN_577; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2155 = ~hit_reg ? valid_array_1_2 : _GEN_578; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2156 = ~hit_reg ? valid_array_1_3 : _GEN_579; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2157 = ~hit_reg ? valid_array_1_4 : _GEN_580; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2158 = ~hit_reg ? valid_array_1_5 : _GEN_581; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2159 = ~hit_reg ? valid_array_1_6 : _GEN_582; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2160 = ~hit_reg ? valid_array_1_7 : _GEN_583; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2161 = ~hit_reg ? valid_array_1_8 : _GEN_584; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2162 = ~hit_reg ? valid_array_1_9 : _GEN_585; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2163 = ~hit_reg ? valid_array_1_10 : _GEN_586; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2164 = ~hit_reg ? valid_array_1_11 : _GEN_587; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2165 = ~hit_reg ? valid_array_1_12 : _GEN_588; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2166 = ~hit_reg ? valid_array_1_13 : _GEN_589; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2167 = ~hit_reg ? valid_array_1_14 : _GEN_590; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2168 = ~hit_reg ? valid_array_1_15 : _GEN_591; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2169 = ~hit_reg ? valid_array_1_16 : _GEN_592; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2170 = ~hit_reg ? valid_array_1_17 : _GEN_593; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2171 = ~hit_reg ? valid_array_1_18 : _GEN_594; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2172 = ~hit_reg ? valid_array_1_19 : _GEN_595; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2173 = ~hit_reg ? valid_array_1_20 : _GEN_596; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2174 = ~hit_reg ? valid_array_1_21 : _GEN_597; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2175 = ~hit_reg ? valid_array_1_22 : _GEN_598; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2176 = ~hit_reg ? valid_array_1_23 : _GEN_599; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2177 = ~hit_reg ? valid_array_1_24 : _GEN_600; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2178 = ~hit_reg ? valid_array_1_25 : _GEN_601; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2179 = ~hit_reg ? valid_array_1_26 : _GEN_602; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2180 = ~hit_reg ? valid_array_1_27 : _GEN_603; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2181 = ~hit_reg ? valid_array_1_28 : _GEN_604; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2182 = ~hit_reg ? valid_array_1_29 : _GEN_605; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2183 = ~hit_reg ? valid_array_1_30 : _GEN_606; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2184 = ~hit_reg ? valid_array_1_31 : _GEN_607; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2185 = ~hit_reg ? valid_array_1_32 : _GEN_608; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2186 = ~hit_reg ? valid_array_1_33 : _GEN_609; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2187 = ~hit_reg ? valid_array_1_34 : _GEN_610; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2188 = ~hit_reg ? valid_array_1_35 : _GEN_611; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2189 = ~hit_reg ? valid_array_1_36 : _GEN_612; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2190 = ~hit_reg ? valid_array_1_37 : _GEN_613; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2191 = ~hit_reg ? valid_array_1_38 : _GEN_614; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2192 = ~hit_reg ? valid_array_1_39 : _GEN_615; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2193 = ~hit_reg ? valid_array_1_40 : _GEN_616; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2194 = ~hit_reg ? valid_array_1_41 : _GEN_617; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2195 = ~hit_reg ? valid_array_1_42 : _GEN_618; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2196 = ~hit_reg ? valid_array_1_43 : _GEN_619; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2197 = ~hit_reg ? valid_array_1_44 : _GEN_620; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2198 = ~hit_reg ? valid_array_1_45 : _GEN_621; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2199 = ~hit_reg ? valid_array_1_46 : _GEN_622; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2200 = ~hit_reg ? valid_array_1_47 : _GEN_623; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2201 = ~hit_reg ? valid_array_1_48 : _GEN_624; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2202 = ~hit_reg ? valid_array_1_49 : _GEN_625; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2203 = ~hit_reg ? valid_array_1_50 : _GEN_626; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2204 = ~hit_reg ? valid_array_1_51 : _GEN_627; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2205 = ~hit_reg ? valid_array_1_52 : _GEN_628; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2206 = ~hit_reg ? valid_array_1_53 : _GEN_629; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2207 = ~hit_reg ? valid_array_1_54 : _GEN_630; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2208 = ~hit_reg ? valid_array_1_55 : _GEN_631; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2209 = ~hit_reg ? valid_array_1_56 : _GEN_632; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2210 = ~hit_reg ? valid_array_1_57 : _GEN_633; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2211 = ~hit_reg ? valid_array_1_58 : _GEN_634; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2212 = ~hit_reg ? valid_array_1_59 : _GEN_635; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2213 = ~hit_reg ? valid_array_1_60 : _GEN_636; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2214 = ~hit_reg ? valid_array_1_61 : _GEN_637; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2215 = ~hit_reg ? valid_array_1_62 : _GEN_638; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2216 = ~hit_reg ? valid_array_1_63 : _GEN_639; // @[DCache.scala 298:28 DCache.scala 116:44]
  wire  _GEN_2217 = ~hit_reg ? dirty_array_1_0 : _GEN_1882; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2218 = ~hit_reg ? dirty_array_1_1 : _GEN_1883; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2219 = ~hit_reg ? dirty_array_1_2 : _GEN_1884; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2220 = ~hit_reg ? dirty_array_1_3 : _GEN_1885; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2221 = ~hit_reg ? dirty_array_1_4 : _GEN_1886; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2222 = ~hit_reg ? dirty_array_1_5 : _GEN_1887; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2223 = ~hit_reg ? dirty_array_1_6 : _GEN_1888; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2224 = ~hit_reg ? dirty_array_1_7 : _GEN_1889; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2225 = ~hit_reg ? dirty_array_1_8 : _GEN_1890; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2226 = ~hit_reg ? dirty_array_1_9 : _GEN_1891; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2227 = ~hit_reg ? dirty_array_1_10 : _GEN_1892; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2228 = ~hit_reg ? dirty_array_1_11 : _GEN_1893; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2229 = ~hit_reg ? dirty_array_1_12 : _GEN_1894; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2230 = ~hit_reg ? dirty_array_1_13 : _GEN_1895; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2231 = ~hit_reg ? dirty_array_1_14 : _GEN_1896; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2232 = ~hit_reg ? dirty_array_1_15 : _GEN_1897; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2233 = ~hit_reg ? dirty_array_1_16 : _GEN_1898; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2234 = ~hit_reg ? dirty_array_1_17 : _GEN_1899; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2235 = ~hit_reg ? dirty_array_1_18 : _GEN_1900; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2236 = ~hit_reg ? dirty_array_1_19 : _GEN_1901; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2237 = ~hit_reg ? dirty_array_1_20 : _GEN_1902; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2238 = ~hit_reg ? dirty_array_1_21 : _GEN_1903; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2239 = ~hit_reg ? dirty_array_1_22 : _GEN_1904; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2240 = ~hit_reg ? dirty_array_1_23 : _GEN_1905; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2241 = ~hit_reg ? dirty_array_1_24 : _GEN_1906; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2242 = ~hit_reg ? dirty_array_1_25 : _GEN_1907; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2243 = ~hit_reg ? dirty_array_1_26 : _GEN_1908; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2244 = ~hit_reg ? dirty_array_1_27 : _GEN_1909; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2245 = ~hit_reg ? dirty_array_1_28 : _GEN_1910; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2246 = ~hit_reg ? dirty_array_1_29 : _GEN_1911; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2247 = ~hit_reg ? dirty_array_1_30 : _GEN_1912; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2248 = ~hit_reg ? dirty_array_1_31 : _GEN_1913; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2249 = ~hit_reg ? dirty_array_1_32 : _GEN_1914; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2250 = ~hit_reg ? dirty_array_1_33 : _GEN_1915; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2251 = ~hit_reg ? dirty_array_1_34 : _GEN_1916; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2252 = ~hit_reg ? dirty_array_1_35 : _GEN_1917; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2253 = ~hit_reg ? dirty_array_1_36 : _GEN_1918; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2254 = ~hit_reg ? dirty_array_1_37 : _GEN_1919; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2255 = ~hit_reg ? dirty_array_1_38 : _GEN_1920; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2256 = ~hit_reg ? dirty_array_1_39 : _GEN_1921; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2257 = ~hit_reg ? dirty_array_1_40 : _GEN_1922; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2258 = ~hit_reg ? dirty_array_1_41 : _GEN_1923; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2259 = ~hit_reg ? dirty_array_1_42 : _GEN_1924; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2260 = ~hit_reg ? dirty_array_1_43 : _GEN_1925; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2261 = ~hit_reg ? dirty_array_1_44 : _GEN_1926; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2262 = ~hit_reg ? dirty_array_1_45 : _GEN_1927; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2263 = ~hit_reg ? dirty_array_1_46 : _GEN_1928; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2264 = ~hit_reg ? dirty_array_1_47 : _GEN_1929; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2265 = ~hit_reg ? dirty_array_1_48 : _GEN_1930; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2266 = ~hit_reg ? dirty_array_1_49 : _GEN_1931; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2267 = ~hit_reg ? dirty_array_1_50 : _GEN_1932; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2268 = ~hit_reg ? dirty_array_1_51 : _GEN_1933; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2269 = ~hit_reg ? dirty_array_1_52 : _GEN_1934; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2270 = ~hit_reg ? dirty_array_1_53 : _GEN_1935; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2271 = ~hit_reg ? dirty_array_1_54 : _GEN_1936; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2272 = ~hit_reg ? dirty_array_1_55 : _GEN_1937; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2273 = ~hit_reg ? dirty_array_1_56 : _GEN_1938; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2274 = ~hit_reg ? dirty_array_1_57 : _GEN_1939; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2275 = ~hit_reg ? dirty_array_1_58 : _GEN_1940; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2276 = ~hit_reg ? dirty_array_1_59 : _GEN_1941; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2277 = ~hit_reg ? dirty_array_1_60 : _GEN_1942; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2278 = ~hit_reg ? dirty_array_1_61 : _GEN_1943; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2279 = ~hit_reg ? dirty_array_1_62 : _GEN_1944; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2280 = ~hit_reg ? dirty_array_1_63 : _GEN_1945; // @[DCache.scala 298:28 DCache.scala 114:44]
  wire  _GEN_2346 = curr_state == 4'h1 ? _GEN_2011 : 1'h1; // @[DCache.scala 297:36 CacheBase.scala 81:13]
  wire [5:0] _GEN_2347 = curr_state == 4'h1 ? _GEN_2012 : array_rd_index; // @[DCache.scala 297:36 CacheBase.scala 82:14]
  wire [127:0] _GEN_2348 = curr_state == 4'h1 ? _GEN_2013 : 128'h0; // @[DCache.scala 297:36 CacheBase.scala 83:15]
  wire [127:0] _GEN_2349 = curr_state == 4'h1 ? _GEN_2014 : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 297:36 CacheBase.scala 84:15]
  wire [127:0] _GEN_2351 = curr_state == 4'h1 ? _GEN_2016 : 128'h0; // @[DCache.scala 297:36 CacheBase.scala 83:15]
  wire  _GEN_2353 = curr_state == 4'h1 ? _GEN_2018 : valid_array_0_0; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2354 = curr_state == 4'h1 ? _GEN_2019 : valid_array_0_1; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2355 = curr_state == 4'h1 ? _GEN_2020 : valid_array_0_2; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2356 = curr_state == 4'h1 ? _GEN_2021 : valid_array_0_3; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2357 = curr_state == 4'h1 ? _GEN_2022 : valid_array_0_4; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2358 = curr_state == 4'h1 ? _GEN_2023 : valid_array_0_5; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2359 = curr_state == 4'h1 ? _GEN_2024 : valid_array_0_6; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2360 = curr_state == 4'h1 ? _GEN_2025 : valid_array_0_7; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2361 = curr_state == 4'h1 ? _GEN_2026 : valid_array_0_8; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2362 = curr_state == 4'h1 ? _GEN_2027 : valid_array_0_9; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2363 = curr_state == 4'h1 ? _GEN_2028 : valid_array_0_10; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2364 = curr_state == 4'h1 ? _GEN_2029 : valid_array_0_11; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2365 = curr_state == 4'h1 ? _GEN_2030 : valid_array_0_12; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2366 = curr_state == 4'h1 ? _GEN_2031 : valid_array_0_13; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2367 = curr_state == 4'h1 ? _GEN_2032 : valid_array_0_14; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2368 = curr_state == 4'h1 ? _GEN_2033 : valid_array_0_15; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2369 = curr_state == 4'h1 ? _GEN_2034 : valid_array_0_16; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2370 = curr_state == 4'h1 ? _GEN_2035 : valid_array_0_17; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2371 = curr_state == 4'h1 ? _GEN_2036 : valid_array_0_18; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2372 = curr_state == 4'h1 ? _GEN_2037 : valid_array_0_19; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2373 = curr_state == 4'h1 ? _GEN_2038 : valid_array_0_20; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2374 = curr_state == 4'h1 ? _GEN_2039 : valid_array_0_21; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2375 = curr_state == 4'h1 ? _GEN_2040 : valid_array_0_22; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2376 = curr_state == 4'h1 ? _GEN_2041 : valid_array_0_23; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2377 = curr_state == 4'h1 ? _GEN_2042 : valid_array_0_24; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2378 = curr_state == 4'h1 ? _GEN_2043 : valid_array_0_25; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2379 = curr_state == 4'h1 ? _GEN_2044 : valid_array_0_26; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2380 = curr_state == 4'h1 ? _GEN_2045 : valid_array_0_27; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2381 = curr_state == 4'h1 ? _GEN_2046 : valid_array_0_28; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2382 = curr_state == 4'h1 ? _GEN_2047 : valid_array_0_29; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2383 = curr_state == 4'h1 ? _GEN_2048 : valid_array_0_30; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2384 = curr_state == 4'h1 ? _GEN_2049 : valid_array_0_31; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2385 = curr_state == 4'h1 ? _GEN_2050 : valid_array_0_32; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2386 = curr_state == 4'h1 ? _GEN_2051 : valid_array_0_33; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2387 = curr_state == 4'h1 ? _GEN_2052 : valid_array_0_34; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2388 = curr_state == 4'h1 ? _GEN_2053 : valid_array_0_35; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2389 = curr_state == 4'h1 ? _GEN_2054 : valid_array_0_36; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2390 = curr_state == 4'h1 ? _GEN_2055 : valid_array_0_37; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2391 = curr_state == 4'h1 ? _GEN_2056 : valid_array_0_38; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2392 = curr_state == 4'h1 ? _GEN_2057 : valid_array_0_39; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2393 = curr_state == 4'h1 ? _GEN_2058 : valid_array_0_40; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2394 = curr_state == 4'h1 ? _GEN_2059 : valid_array_0_41; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2395 = curr_state == 4'h1 ? _GEN_2060 : valid_array_0_42; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2396 = curr_state == 4'h1 ? _GEN_2061 : valid_array_0_43; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2397 = curr_state == 4'h1 ? _GEN_2062 : valid_array_0_44; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2398 = curr_state == 4'h1 ? _GEN_2063 : valid_array_0_45; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2399 = curr_state == 4'h1 ? _GEN_2064 : valid_array_0_46; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2400 = curr_state == 4'h1 ? _GEN_2065 : valid_array_0_47; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2401 = curr_state == 4'h1 ? _GEN_2066 : valid_array_0_48; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2402 = curr_state == 4'h1 ? _GEN_2067 : valid_array_0_49; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2403 = curr_state == 4'h1 ? _GEN_2068 : valid_array_0_50; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2404 = curr_state == 4'h1 ? _GEN_2069 : valid_array_0_51; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2405 = curr_state == 4'h1 ? _GEN_2070 : valid_array_0_52; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2406 = curr_state == 4'h1 ? _GEN_2071 : valid_array_0_53; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2407 = curr_state == 4'h1 ? _GEN_2072 : valid_array_0_54; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2408 = curr_state == 4'h1 ? _GEN_2073 : valid_array_0_55; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2409 = curr_state == 4'h1 ? _GEN_2074 : valid_array_0_56; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2410 = curr_state == 4'h1 ? _GEN_2075 : valid_array_0_57; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2411 = curr_state == 4'h1 ? _GEN_2076 : valid_array_0_58; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2412 = curr_state == 4'h1 ? _GEN_2077 : valid_array_0_59; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2413 = curr_state == 4'h1 ? _GEN_2078 : valid_array_0_60; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2414 = curr_state == 4'h1 ? _GEN_2079 : valid_array_0_61; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2415 = curr_state == 4'h1 ? _GEN_2080 : valid_array_0_62; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2416 = curr_state == 4'h1 ? _GEN_2081 : valid_array_0_63; // @[DCache.scala 297:36 DCache.scala 115:44]
  wire  _GEN_2417 = curr_state == 4'h1 ? _GEN_2082 : dirty_array_0_0; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2418 = curr_state == 4'h1 ? _GEN_2083 : dirty_array_0_1; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2419 = curr_state == 4'h1 ? _GEN_2084 : dirty_array_0_2; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2420 = curr_state == 4'h1 ? _GEN_2085 : dirty_array_0_3; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2421 = curr_state == 4'h1 ? _GEN_2086 : dirty_array_0_4; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2422 = curr_state == 4'h1 ? _GEN_2087 : dirty_array_0_5; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2423 = curr_state == 4'h1 ? _GEN_2088 : dirty_array_0_6; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2424 = curr_state == 4'h1 ? _GEN_2089 : dirty_array_0_7; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2425 = curr_state == 4'h1 ? _GEN_2090 : dirty_array_0_8; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2426 = curr_state == 4'h1 ? _GEN_2091 : dirty_array_0_9; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2427 = curr_state == 4'h1 ? _GEN_2092 : dirty_array_0_10; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2428 = curr_state == 4'h1 ? _GEN_2093 : dirty_array_0_11; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2429 = curr_state == 4'h1 ? _GEN_2094 : dirty_array_0_12; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2430 = curr_state == 4'h1 ? _GEN_2095 : dirty_array_0_13; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2431 = curr_state == 4'h1 ? _GEN_2096 : dirty_array_0_14; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2432 = curr_state == 4'h1 ? _GEN_2097 : dirty_array_0_15; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2433 = curr_state == 4'h1 ? _GEN_2098 : dirty_array_0_16; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2434 = curr_state == 4'h1 ? _GEN_2099 : dirty_array_0_17; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2435 = curr_state == 4'h1 ? _GEN_2100 : dirty_array_0_18; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2436 = curr_state == 4'h1 ? _GEN_2101 : dirty_array_0_19; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2437 = curr_state == 4'h1 ? _GEN_2102 : dirty_array_0_20; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2438 = curr_state == 4'h1 ? _GEN_2103 : dirty_array_0_21; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2439 = curr_state == 4'h1 ? _GEN_2104 : dirty_array_0_22; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2440 = curr_state == 4'h1 ? _GEN_2105 : dirty_array_0_23; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2441 = curr_state == 4'h1 ? _GEN_2106 : dirty_array_0_24; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2442 = curr_state == 4'h1 ? _GEN_2107 : dirty_array_0_25; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2443 = curr_state == 4'h1 ? _GEN_2108 : dirty_array_0_26; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2444 = curr_state == 4'h1 ? _GEN_2109 : dirty_array_0_27; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2445 = curr_state == 4'h1 ? _GEN_2110 : dirty_array_0_28; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2446 = curr_state == 4'h1 ? _GEN_2111 : dirty_array_0_29; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2447 = curr_state == 4'h1 ? _GEN_2112 : dirty_array_0_30; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2448 = curr_state == 4'h1 ? _GEN_2113 : dirty_array_0_31; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2449 = curr_state == 4'h1 ? _GEN_2114 : dirty_array_0_32; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2450 = curr_state == 4'h1 ? _GEN_2115 : dirty_array_0_33; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2451 = curr_state == 4'h1 ? _GEN_2116 : dirty_array_0_34; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2452 = curr_state == 4'h1 ? _GEN_2117 : dirty_array_0_35; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2453 = curr_state == 4'h1 ? _GEN_2118 : dirty_array_0_36; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2454 = curr_state == 4'h1 ? _GEN_2119 : dirty_array_0_37; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2455 = curr_state == 4'h1 ? _GEN_2120 : dirty_array_0_38; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2456 = curr_state == 4'h1 ? _GEN_2121 : dirty_array_0_39; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2457 = curr_state == 4'h1 ? _GEN_2122 : dirty_array_0_40; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2458 = curr_state == 4'h1 ? _GEN_2123 : dirty_array_0_41; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2459 = curr_state == 4'h1 ? _GEN_2124 : dirty_array_0_42; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2460 = curr_state == 4'h1 ? _GEN_2125 : dirty_array_0_43; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2461 = curr_state == 4'h1 ? _GEN_2126 : dirty_array_0_44; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2462 = curr_state == 4'h1 ? _GEN_2127 : dirty_array_0_45; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2463 = curr_state == 4'h1 ? _GEN_2128 : dirty_array_0_46; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2464 = curr_state == 4'h1 ? _GEN_2129 : dirty_array_0_47; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2465 = curr_state == 4'h1 ? _GEN_2130 : dirty_array_0_48; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2466 = curr_state == 4'h1 ? _GEN_2131 : dirty_array_0_49; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2467 = curr_state == 4'h1 ? _GEN_2132 : dirty_array_0_50; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2468 = curr_state == 4'h1 ? _GEN_2133 : dirty_array_0_51; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2469 = curr_state == 4'h1 ? _GEN_2134 : dirty_array_0_52; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2470 = curr_state == 4'h1 ? _GEN_2135 : dirty_array_0_53; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2471 = curr_state == 4'h1 ? _GEN_2136 : dirty_array_0_54; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2472 = curr_state == 4'h1 ? _GEN_2137 : dirty_array_0_55; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2473 = curr_state == 4'h1 ? _GEN_2138 : dirty_array_0_56; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2474 = curr_state == 4'h1 ? _GEN_2139 : dirty_array_0_57; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2475 = curr_state == 4'h1 ? _GEN_2140 : dirty_array_0_58; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2476 = curr_state == 4'h1 ? _GEN_2141 : dirty_array_0_59; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2477 = curr_state == 4'h1 ? _GEN_2142 : dirty_array_0_60; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2478 = curr_state == 4'h1 ? _GEN_2143 : dirty_array_0_61; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2479 = curr_state == 4'h1 ? _GEN_2144 : dirty_array_0_62; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2480 = curr_state == 4'h1 ? _GEN_2145 : dirty_array_0_63; // @[DCache.scala 297:36 DCache.scala 113:44]
  wire  _GEN_2481 = curr_state == 4'h1 ? _T_20 : 1'h1; // @[DCache.scala 297:36 CacheBase.scala 81:13]
  wire [5:0] _GEN_2482 = curr_state == 4'h1 ? _GEN_2147 : array_rd_index; // @[DCache.scala 297:36 CacheBase.scala 82:14]
  wire [127:0] _GEN_2483 = curr_state == 4'h1 ? _GEN_2148 : 128'h0; // @[DCache.scala 297:36 CacheBase.scala 83:15]
  wire [127:0] _GEN_2484 = curr_state == 4'h1 ? _GEN_2149 : 128'hffffffffffffffffffffffffffffffff; // @[DCache.scala 297:36 CacheBase.scala 84:15]
  wire [127:0] _GEN_2486 = curr_state == 4'h1 ? _GEN_2151 : 128'h0; // @[DCache.scala 297:36 CacheBase.scala 83:15]
  wire  _GEN_2488 = curr_state == 4'h1 ? _GEN_2153 : valid_array_1_0; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2489 = curr_state == 4'h1 ? _GEN_2154 : valid_array_1_1; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2490 = curr_state == 4'h1 ? _GEN_2155 : valid_array_1_2; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2491 = curr_state == 4'h1 ? _GEN_2156 : valid_array_1_3; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2492 = curr_state == 4'h1 ? _GEN_2157 : valid_array_1_4; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2493 = curr_state == 4'h1 ? _GEN_2158 : valid_array_1_5; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2494 = curr_state == 4'h1 ? _GEN_2159 : valid_array_1_6; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2495 = curr_state == 4'h1 ? _GEN_2160 : valid_array_1_7; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2496 = curr_state == 4'h1 ? _GEN_2161 : valid_array_1_8; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2497 = curr_state == 4'h1 ? _GEN_2162 : valid_array_1_9; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2498 = curr_state == 4'h1 ? _GEN_2163 : valid_array_1_10; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2499 = curr_state == 4'h1 ? _GEN_2164 : valid_array_1_11; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2500 = curr_state == 4'h1 ? _GEN_2165 : valid_array_1_12; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2501 = curr_state == 4'h1 ? _GEN_2166 : valid_array_1_13; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2502 = curr_state == 4'h1 ? _GEN_2167 : valid_array_1_14; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2503 = curr_state == 4'h1 ? _GEN_2168 : valid_array_1_15; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2504 = curr_state == 4'h1 ? _GEN_2169 : valid_array_1_16; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2505 = curr_state == 4'h1 ? _GEN_2170 : valid_array_1_17; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2506 = curr_state == 4'h1 ? _GEN_2171 : valid_array_1_18; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2507 = curr_state == 4'h1 ? _GEN_2172 : valid_array_1_19; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2508 = curr_state == 4'h1 ? _GEN_2173 : valid_array_1_20; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2509 = curr_state == 4'h1 ? _GEN_2174 : valid_array_1_21; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2510 = curr_state == 4'h1 ? _GEN_2175 : valid_array_1_22; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2511 = curr_state == 4'h1 ? _GEN_2176 : valid_array_1_23; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2512 = curr_state == 4'h1 ? _GEN_2177 : valid_array_1_24; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2513 = curr_state == 4'h1 ? _GEN_2178 : valid_array_1_25; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2514 = curr_state == 4'h1 ? _GEN_2179 : valid_array_1_26; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2515 = curr_state == 4'h1 ? _GEN_2180 : valid_array_1_27; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2516 = curr_state == 4'h1 ? _GEN_2181 : valid_array_1_28; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2517 = curr_state == 4'h1 ? _GEN_2182 : valid_array_1_29; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2518 = curr_state == 4'h1 ? _GEN_2183 : valid_array_1_30; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2519 = curr_state == 4'h1 ? _GEN_2184 : valid_array_1_31; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2520 = curr_state == 4'h1 ? _GEN_2185 : valid_array_1_32; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2521 = curr_state == 4'h1 ? _GEN_2186 : valid_array_1_33; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2522 = curr_state == 4'h1 ? _GEN_2187 : valid_array_1_34; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2523 = curr_state == 4'h1 ? _GEN_2188 : valid_array_1_35; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2524 = curr_state == 4'h1 ? _GEN_2189 : valid_array_1_36; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2525 = curr_state == 4'h1 ? _GEN_2190 : valid_array_1_37; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2526 = curr_state == 4'h1 ? _GEN_2191 : valid_array_1_38; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2527 = curr_state == 4'h1 ? _GEN_2192 : valid_array_1_39; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2528 = curr_state == 4'h1 ? _GEN_2193 : valid_array_1_40; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2529 = curr_state == 4'h1 ? _GEN_2194 : valid_array_1_41; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2530 = curr_state == 4'h1 ? _GEN_2195 : valid_array_1_42; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2531 = curr_state == 4'h1 ? _GEN_2196 : valid_array_1_43; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2532 = curr_state == 4'h1 ? _GEN_2197 : valid_array_1_44; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2533 = curr_state == 4'h1 ? _GEN_2198 : valid_array_1_45; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2534 = curr_state == 4'h1 ? _GEN_2199 : valid_array_1_46; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2535 = curr_state == 4'h1 ? _GEN_2200 : valid_array_1_47; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2536 = curr_state == 4'h1 ? _GEN_2201 : valid_array_1_48; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2537 = curr_state == 4'h1 ? _GEN_2202 : valid_array_1_49; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2538 = curr_state == 4'h1 ? _GEN_2203 : valid_array_1_50; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2539 = curr_state == 4'h1 ? _GEN_2204 : valid_array_1_51; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2540 = curr_state == 4'h1 ? _GEN_2205 : valid_array_1_52; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2541 = curr_state == 4'h1 ? _GEN_2206 : valid_array_1_53; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2542 = curr_state == 4'h1 ? _GEN_2207 : valid_array_1_54; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2543 = curr_state == 4'h1 ? _GEN_2208 : valid_array_1_55; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2544 = curr_state == 4'h1 ? _GEN_2209 : valid_array_1_56; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2545 = curr_state == 4'h1 ? _GEN_2210 : valid_array_1_57; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2546 = curr_state == 4'h1 ? _GEN_2211 : valid_array_1_58; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2547 = curr_state == 4'h1 ? _GEN_2212 : valid_array_1_59; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2548 = curr_state == 4'h1 ? _GEN_2213 : valid_array_1_60; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2549 = curr_state == 4'h1 ? _GEN_2214 : valid_array_1_61; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2550 = curr_state == 4'h1 ? _GEN_2215 : valid_array_1_62; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2551 = curr_state == 4'h1 ? _GEN_2216 : valid_array_1_63; // @[DCache.scala 297:36 DCache.scala 116:44]
  wire  _GEN_2552 = curr_state == 4'h1 ? _GEN_2217 : dirty_array_1_0; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2553 = curr_state == 4'h1 ? _GEN_2218 : dirty_array_1_1; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2554 = curr_state == 4'h1 ? _GEN_2219 : dirty_array_1_2; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2555 = curr_state == 4'h1 ? _GEN_2220 : dirty_array_1_3; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2556 = curr_state == 4'h1 ? _GEN_2221 : dirty_array_1_4; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2557 = curr_state == 4'h1 ? _GEN_2222 : dirty_array_1_5; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2558 = curr_state == 4'h1 ? _GEN_2223 : dirty_array_1_6; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2559 = curr_state == 4'h1 ? _GEN_2224 : dirty_array_1_7; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2560 = curr_state == 4'h1 ? _GEN_2225 : dirty_array_1_8; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2561 = curr_state == 4'h1 ? _GEN_2226 : dirty_array_1_9; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2562 = curr_state == 4'h1 ? _GEN_2227 : dirty_array_1_10; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2563 = curr_state == 4'h1 ? _GEN_2228 : dirty_array_1_11; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2564 = curr_state == 4'h1 ? _GEN_2229 : dirty_array_1_12; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2565 = curr_state == 4'h1 ? _GEN_2230 : dirty_array_1_13; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2566 = curr_state == 4'h1 ? _GEN_2231 : dirty_array_1_14; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2567 = curr_state == 4'h1 ? _GEN_2232 : dirty_array_1_15; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2568 = curr_state == 4'h1 ? _GEN_2233 : dirty_array_1_16; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2569 = curr_state == 4'h1 ? _GEN_2234 : dirty_array_1_17; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2570 = curr_state == 4'h1 ? _GEN_2235 : dirty_array_1_18; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2571 = curr_state == 4'h1 ? _GEN_2236 : dirty_array_1_19; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2572 = curr_state == 4'h1 ? _GEN_2237 : dirty_array_1_20; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2573 = curr_state == 4'h1 ? _GEN_2238 : dirty_array_1_21; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2574 = curr_state == 4'h1 ? _GEN_2239 : dirty_array_1_22; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2575 = curr_state == 4'h1 ? _GEN_2240 : dirty_array_1_23; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2576 = curr_state == 4'h1 ? _GEN_2241 : dirty_array_1_24; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2577 = curr_state == 4'h1 ? _GEN_2242 : dirty_array_1_25; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2578 = curr_state == 4'h1 ? _GEN_2243 : dirty_array_1_26; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2579 = curr_state == 4'h1 ? _GEN_2244 : dirty_array_1_27; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2580 = curr_state == 4'h1 ? _GEN_2245 : dirty_array_1_28; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2581 = curr_state == 4'h1 ? _GEN_2246 : dirty_array_1_29; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2582 = curr_state == 4'h1 ? _GEN_2247 : dirty_array_1_30; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2583 = curr_state == 4'h1 ? _GEN_2248 : dirty_array_1_31; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2584 = curr_state == 4'h1 ? _GEN_2249 : dirty_array_1_32; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2585 = curr_state == 4'h1 ? _GEN_2250 : dirty_array_1_33; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2586 = curr_state == 4'h1 ? _GEN_2251 : dirty_array_1_34; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2587 = curr_state == 4'h1 ? _GEN_2252 : dirty_array_1_35; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2588 = curr_state == 4'h1 ? _GEN_2253 : dirty_array_1_36; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2589 = curr_state == 4'h1 ? _GEN_2254 : dirty_array_1_37; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2590 = curr_state == 4'h1 ? _GEN_2255 : dirty_array_1_38; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2591 = curr_state == 4'h1 ? _GEN_2256 : dirty_array_1_39; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2592 = curr_state == 4'h1 ? _GEN_2257 : dirty_array_1_40; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2593 = curr_state == 4'h1 ? _GEN_2258 : dirty_array_1_41; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2594 = curr_state == 4'h1 ? _GEN_2259 : dirty_array_1_42; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2595 = curr_state == 4'h1 ? _GEN_2260 : dirty_array_1_43; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2596 = curr_state == 4'h1 ? _GEN_2261 : dirty_array_1_44; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2597 = curr_state == 4'h1 ? _GEN_2262 : dirty_array_1_45; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2598 = curr_state == 4'h1 ? _GEN_2263 : dirty_array_1_46; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2599 = curr_state == 4'h1 ? _GEN_2264 : dirty_array_1_47; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2600 = curr_state == 4'h1 ? _GEN_2265 : dirty_array_1_48; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2601 = curr_state == 4'h1 ? _GEN_2266 : dirty_array_1_49; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2602 = curr_state == 4'h1 ? _GEN_2267 : dirty_array_1_50; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2603 = curr_state == 4'h1 ? _GEN_2268 : dirty_array_1_51; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2604 = curr_state == 4'h1 ? _GEN_2269 : dirty_array_1_52; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2605 = curr_state == 4'h1 ? _GEN_2270 : dirty_array_1_53; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2606 = curr_state == 4'h1 ? _GEN_2271 : dirty_array_1_54; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2607 = curr_state == 4'h1 ? _GEN_2272 : dirty_array_1_55; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2608 = curr_state == 4'h1 ? _GEN_2273 : dirty_array_1_56; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2609 = curr_state == 4'h1 ? _GEN_2274 : dirty_array_1_57; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2610 = curr_state == 4'h1 ? _GEN_2275 : dirty_array_1_58; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2611 = curr_state == 4'h1 ? _GEN_2276 : dirty_array_1_59; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2612 = curr_state == 4'h1 ? _GEN_2277 : dirty_array_1_60; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2613 = curr_state == 4'h1 ? _GEN_2278 : dirty_array_1_61; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2614 = curr_state == 4'h1 ? _GEN_2279 : dirty_array_1_62; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2615 = curr_state == 4'h1 ? _GEN_2280 : dirty_array_1_63; // @[DCache.scala 297:36 DCache.scala 114:44]
  wire  _GEN_2681 = curr_state == 4'hb ? _GEN_1424 : _GEN_2481; // @[DCache.scala 286:38]
  wire [5:0] _GEN_2682 = curr_state == 4'hb ? _GEN_1425 : _GEN_2482; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2683 = curr_state == 4'hb ? 128'h0 : _GEN_2483; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2684 = curr_state == 4'hb ? _GEN_1426 : _GEN_2484; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2686 = curr_state == 4'hb ? 128'h0 : _GEN_2486; // @[DCache.scala 286:38]
  wire  _GEN_2688 = curr_state == 4'hb ? flush_way : _GEN_2346; // @[DCache.scala 286:38]
  wire [5:0] _GEN_2689 = curr_state == 4'hb ? _GEN_1430 : _GEN_2347; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2690 = curr_state == 4'hb ? 128'h0 : _GEN_2348; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2691 = curr_state == 4'hb ? _GEN_1431 : _GEN_2349; // @[DCache.scala 286:38]
  wire [127:0] _GEN_2693 = curr_state == 4'hb ? 128'h0 : _GEN_2351; // @[DCache.scala 286:38]
  wire [190:0] _GEN_4096 = {{127'd0}, mmio_manager_io_out_data}; // @[DCache.scala 405:37]
  wire [190:0] _read_data_128_T = _GEN_4096 << save_start_bit_lshift2; // @[DCache.scala 405:37]
  wire [190:0] _read_data_128_T_1 = addr_underflow ? _read_data_128_T : {{63'd0}, maxi4_manager_io_out_data}; // @[Mux.scala 98:16]
  wire [190:0] read_data_128 = hit_reg_x8 ? {{63'd0}, cache_line_data_out} : _read_data_128_T_1; // @[Mux.scala 98:16]
  wire [190:0] _read_data_64_T = read_data_128 >> save_start_bit_lshift2; // @[DCache.scala 410:46]
  wire [63:0] read_data_64 = _read_data_64_T[63:0]; // @[DCache.scala 410:59]
  wire [63:0] _raw_read_data_T_3 = stage1_out_bits_size_dword ? read_data_64 : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _raw_read_data_T_4 = stage1_out_bits_size_word ? {{32'd0}, read_data_64[31:0]} : _raw_read_data_T_3; // @[Mux.scala 98:16]
  wire [63:0] _raw_read_data_T_5 = stage1_out_bits_size_hword ? {{48'd0}, read_data_64[15:0]} : _raw_read_data_T_4; // @[Mux.scala 98:16]
  wire [63:0] raw_read_data = stage1_out_bits_size_byte ? {{56'd0}, read_data_64[7:0]} : _raw_read_data_T_5; // @[Mux.scala 98:16]
  wire [63:0] _sext_memory_data_signed_T = stage1_out_bits_size_byte ? {{56'd0}, read_data_64[7:0]} : _raw_read_data_T_5
    ; // @[DCache.scala 420:52]
  wire [7:0] _sext_memory_data_signed_T_2 = raw_read_data[7:0]; // @[DCache.scala 422:52]
  wire [15:0] _sext_memory_data_signed_T_4 = raw_read_data[15:0]; // @[DCache.scala 423:53]
  wire [31:0] _sext_memory_data_signed_T_6 = raw_read_data[31:0]; // @[DCache.scala 424:53]
  wire [63:0] _sext_memory_data_signed_T_9 = stage1_out_bits_size_dword ? $signed(_sext_memory_data_signed_T) : $signed(
    _sext_memory_data_signed_T); // @[Mux.scala 98:16]
  wire [63:0] _sext_memory_data_signed_T_10 = stage1_out_bits_size_word ? $signed({{32{_sext_memory_data_signed_T_6[31
    ]}},_sext_memory_data_signed_T_6}) : $signed(_sext_memory_data_signed_T_9); // @[Mux.scala 98:16]
  wire [63:0] _sext_memory_data_signed_T_11 = stage1_out_bits_size_hword ? $signed({{48{_sext_memory_data_signed_T_4[15
    ]}},_sext_memory_data_signed_T_4}) : $signed(_sext_memory_data_signed_T_10); // @[Mux.scala 98:16]
  wire [63:0] sext_memory_data = stage1_out_bits_size_byte ? $signed({{56{_sext_memory_data_signed_T_2[7]}},
    _sext_memory_data_signed_T_2}) : $signed(_sext_memory_data_signed_T_11); // @[DCache.scala 428:58]
  ysyx_040978_DAXIManager maxi4_manager ( // @[DCache.scala 70:29]
    .clock(maxi4_manager_clock),
    .reset(maxi4_manager_reset),
    .io_in_rd_en(maxi4_manager_io_in_rd_en),
    .io_in_we_en(maxi4_manager_io_in_we_en),
    .io_in_addr(maxi4_manager_io_in_addr),
    .io_in_data(maxi4_manager_io_in_data),
    .io_maxi_ar_ready(maxi4_manager_io_maxi_ar_ready),
    .io_maxi_ar_valid(maxi4_manager_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(maxi4_manager_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(maxi4_manager_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(maxi4_manager_io_maxi_ar_bits_size),
    .io_maxi_r_valid(maxi4_manager_io_maxi_r_valid),
    .io_maxi_r_bits_data(maxi4_manager_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(maxi4_manager_io_maxi_r_bits_last),
    .io_maxi_aw_ready(maxi4_manager_io_maxi_aw_ready),
    .io_maxi_aw_valid(maxi4_manager_io_maxi_aw_valid),
    .io_maxi_aw_bits_addr(maxi4_manager_io_maxi_aw_bits_addr),
    .io_maxi_aw_bits_len(maxi4_manager_io_maxi_aw_bits_len),
    .io_maxi_aw_bits_size(maxi4_manager_io_maxi_aw_bits_size),
    .io_maxi_w_ready(maxi4_manager_io_maxi_w_ready),
    .io_maxi_w_valid(maxi4_manager_io_maxi_w_valid),
    .io_maxi_w_bits_data(maxi4_manager_io_maxi_w_bits_data),
    .io_maxi_w_bits_strb(maxi4_manager_io_maxi_w_bits_strb),
    .io_maxi_w_bits_last(maxi4_manager_io_maxi_w_bits_last),
    .io_maxi_b_valid(maxi4_manager_io_maxi_b_valid),
    .io_out_finish(maxi4_manager_io_out_finish),
    .io_out_ready(maxi4_manager_io_out_ready),
    .io_out_data(maxi4_manager_io_out_data)
  );
  ysyx_040978_AXI4LiteManager mmio_manager ( // @[DCache.scala 83:28]
    .clock(mmio_manager_clock),
    .reset(mmio_manager_reset),
    .io_in_rd_en(mmio_manager_io_in_rd_en),
    .io_in_we_en(mmio_manager_io_in_we_en),
    .io_in_size_byte(mmio_manager_io_in_size_byte),
    .io_in_size_hword(mmio_manager_io_in_size_hword),
    .io_in_size_word(mmio_manager_io_in_size_word),
    .io_in_size_dword(mmio_manager_io_in_size_dword),
    .io_in_addr(mmio_manager_io_in_addr),
    .io_in_data(mmio_manager_io_in_data),
    .io_in_wmask(mmio_manager_io_in_wmask),
    .io_maxi_ar_ready(mmio_manager_io_maxi_ar_ready),
    .io_maxi_ar_valid(mmio_manager_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(mmio_manager_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_size(mmio_manager_io_maxi_ar_bits_size),
    .io_maxi_r_valid(mmio_manager_io_maxi_r_valid),
    .io_maxi_r_bits_data(mmio_manager_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(mmio_manager_io_maxi_r_bits_last),
    .io_maxi_aw_ready(mmio_manager_io_maxi_aw_ready),
    .io_maxi_aw_valid(mmio_manager_io_maxi_aw_valid),
    .io_maxi_aw_bits_addr(mmio_manager_io_maxi_aw_bits_addr),
    .io_maxi_aw_bits_size(mmio_manager_io_maxi_aw_bits_size),
    .io_maxi_w_ready(mmio_manager_io_maxi_w_ready),
    .io_maxi_w_valid(mmio_manager_io_maxi_w_valid),
    .io_maxi_w_bits_data(mmio_manager_io_maxi_w_bits_data),
    .io_maxi_w_bits_strb(mmio_manager_io_maxi_w_bits_strb),
    .io_maxi_w_bits_last(mmio_manager_io_maxi_w_bits_last),
    .io_maxi_b_valid(mmio_manager_io_maxi_b_valid),
    .io_out_finish(mmio_manager_io_out_finish),
    .io_out_ready(mmio_manager_io_out_ready),
    .io_out_data(mmio_manager_io_out_data),
    .clint_we_0(mmio_manager_clint_we_0),
    ._T_24_0(mmio_manager__T_24_0),
    .clint_rdata_0(mmio_manager_clint_rdata_0),
    .clint_wdata_0(mmio_manager_clint_wdata_0)
  );
  assign io_next_valid = go_on & stage1_out_valid; // @[DCache.scala 475:30]
  assign io_next_bits_data_id2wb_intr_exce_ret = stage1_out_bits_data_id2wb_intr_exce_ret; // @[DCache.scala 473:24]
  assign io_next_bits_data_id2wb_fencei = stage1_out_bits_data_id2wb_fencei; // @[DCache.scala 473:24]
  assign io_next_bits_data_id2wb_wb_sel = stage1_out_bits_data_id2wb_wb_sel; // @[DCache.scala 473:24]
  assign io_next_bits_data_id2wb_regfile_we_en = stage1_out_bits_data_id2wb_regfile_we_en; // @[DCache.scala 473:24]
  assign io_next_bits_data_id2wb_regfile_we_addr = stage1_out_bits_data_id2wb_regfile_we_addr; // @[DCache.scala 473:24]
  assign io_next_bits_data_ex2wb_result_data = stage1_out_bits_data_ex2wb_result_data; // @[DCache.scala 474:24]
  assign io_next_bits_data_mem2wb_memory_data = stage1_out_bits_data_id2mem_sext_flag ? sext_memory_data : raw_read_data
    ; // @[DCache.scala 429:30]
  assign io_prev_ready = next_state == 4'h0; // @[DCache.scala 185:46]
  assign io_maxi_ar_valid = maxi4_manager_io_maxi_ar_valid; // @[DCache.scala 71:25]
  assign io_maxi_ar_bits_addr = maxi4_manager_io_maxi_ar_bits_addr; // @[DCache.scala 71:25]
  assign io_maxi_ar_bits_len = maxi4_manager_io_maxi_ar_bits_len; // @[DCache.scala 71:25]
  assign io_maxi_ar_bits_size = maxi4_manager_io_maxi_ar_bits_size; // @[DCache.scala 71:25]
  assign io_maxi_aw_valid = maxi4_manager_io_maxi_aw_valid; // @[DCache.scala 71:25]
  assign io_maxi_aw_bits_addr = maxi4_manager_io_maxi_aw_bits_addr; // @[DCache.scala 71:25]
  assign io_maxi_aw_bits_len = maxi4_manager_io_maxi_aw_bits_len; // @[DCache.scala 71:25]
  assign io_maxi_aw_bits_size = maxi4_manager_io_maxi_aw_bits_size; // @[DCache.scala 71:25]
  assign io_maxi_w_valid = maxi4_manager_io_maxi_w_valid; // @[DCache.scala 71:25]
  assign io_maxi_w_bits_data = maxi4_manager_io_maxi_w_bits_data; // @[DCache.scala 71:25]
  assign io_maxi_w_bits_strb = maxi4_manager_io_maxi_w_bits_strb; // @[DCache.scala 71:25]
  assign io_maxi_w_bits_last = maxi4_manager_io_maxi_w_bits_last; // @[DCache.scala 71:25]
  assign io_mmio_ar_valid = mmio_manager_io_maxi_ar_valid; // @[DCache.scala 84:24]
  assign io_mmio_ar_bits_addr = mmio_manager_io_maxi_ar_bits_addr; // @[DCache.scala 84:24]
  assign io_mmio_ar_bits_size = mmio_manager_io_maxi_ar_bits_size; // @[DCache.scala 84:24]
  assign io_mmio_aw_valid = mmio_manager_io_maxi_aw_valid; // @[DCache.scala 84:24]
  assign io_mmio_aw_bits_addr = mmio_manager_io_maxi_aw_bits_addr; // @[DCache.scala 84:24]
  assign io_mmio_aw_bits_size = mmio_manager_io_maxi_aw_bits_size; // @[DCache.scala 84:24]
  assign io_mmio_w_valid = mmio_manager_io_maxi_w_valid; // @[DCache.scala 84:24]
  assign io_mmio_w_bits_data = mmio_manager_io_maxi_w_bits_data; // @[DCache.scala 84:24]
  assign io_mmio_w_bits_strb = mmio_manager_io_maxi_w_bits_strb; // @[DCache.scala 84:24]
  assign io_mmio_w_bits_last = mmio_manager_io_maxi_w_bits_last; // @[DCache.scala 84:24]
  assign io_sram4_addr = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1097 : _GEN_2689; // @[DCache.scala 269:43]
  assign io_sram4_wen = curr_state == 4'h2 & maxi4_manager_io_out_finish ? next_way : _GEN_2688; // @[DCache.scala 269:43]
  assign io_sram4_wmask = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1099 : _GEN_2691; // @[DCache.scala 269:43]
  assign io_sram4_wdata = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1098 : _GEN_2690; // @[DCache.scala 269:43]
  assign io_sram5_addr = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_962 : _GEN_2682; // @[DCache.scala 269:43]
  assign io_sram5_wen = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_961 : _GEN_2681; // @[DCache.scala 269:43]
  assign io_sram5_wmask = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_964 : _GEN_2684; // @[DCache.scala 269:43]
  assign io_sram5_wdata = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_963 : _GEN_2683; // @[DCache.scala 269:43]
  assign io_sram6_addr = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1097 : _GEN_2689; // @[DCache.scala 269:43]
  assign io_sram6_wen = curr_state == 4'h2 & maxi4_manager_io_out_finish ? next_way : _GEN_2688; // @[DCache.scala 269:43]
  assign io_sram6_wmask = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1099 : _GEN_2691; // @[DCache.scala 269:43]
  assign io_sram6_wdata = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_1101 : _GEN_2693; // @[DCache.scala 269:43]
  assign io_sram7_addr = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_962 : _GEN_2682; // @[DCache.scala 269:43]
  assign io_sram7_wen = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_961 : _GEN_2681; // @[DCache.scala 269:43]
  assign io_sram7_wmask = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_964 : _GEN_2684; // @[DCache.scala 269:43]
  assign io_sram7_wdata = curr_state == 4'h2 & maxi4_manager_io_out_finish ? _GEN_966 : _GEN_2686; // @[DCache.scala 269:43]
  assign clint_we = mmio_manager_clint_we_0;
  assign _T_24_0 = mmio_manager__T_24_0;
  assign clint_wdata = mmio_manager_clint_wdata_0;
  assign maxi4_manager_clock = clock;
  assign maxi4_manager_reset = reset;
  assign maxi4_manager_io_in_rd_en = curr_state == 4'ha ? 1'h0 : _GEN_498; // @[DCache.scala 205:30 DCache.scala 203:14]
  assign maxi4_manager_io_in_we_en = curr_state == 4'ha | _GEN_497; // @[DCache.scala 205:30 DCache.scala 205:43]
  assign maxi4_manager_io_in_addr = _maxi4_manager_io_in_addr_T_5[31:0]; // @[DCache.scala 219:13]
  assign maxi4_manager_io_in_data = _T ? flush_wb_data : _maxi4_manager_io_in_data_T_3; // @[Mux.scala 98:16]
  assign maxi4_manager_io_maxi_ar_ready = io_maxi_ar_ready; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_r_valid = io_maxi_r_valid; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_r_bits_data = io_maxi_r_bits_data; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_r_bits_last = io_maxi_r_bits_last; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_aw_ready = io_maxi_aw_ready; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_w_ready = io_maxi_w_ready; // @[DCache.scala 71:25]
  assign maxi4_manager_io_maxi_b_valid = io_maxi_b_valid; // @[DCache.scala 71:25]
  assign mmio_manager_clock = clock;
  assign mmio_manager_reset = reset;
  assign mmio_manager_io_in_rd_en = hit_reg_x8 & addr_underflow ? _GEN_503 : _GEN_505; // @[DCache.scala 231:48]
  assign mmio_manager_io_in_we_en = hit_reg_x8 & addr_underflow ? stage1_out_bits_data_id2mem_memory_we_en : _GEN_504; // @[DCache.scala 231:48]
  assign mmio_manager_io_in_size_byte = stage1_out_bits_size_byte; // @[DCache.scala 242:13]
  assign mmio_manager_io_in_size_hword = stage1_out_bits_size_hword; // @[DCache.scala 242:13]
  assign mmio_manager_io_in_size_word = stage1_out_bits_size_word; // @[DCache.scala 242:13]
  assign mmio_manager_io_in_size_dword = stage1_out_bits_size_dword; // @[DCache.scala 242:13]
  assign mmio_manager_io_in_addr = stage1_out_bits_addr[31:0]; // @[DCache.scala 239:13]
  assign mmio_manager_io_in_data = stage1_out_bits_wdata; // @[DCache.scala 240:14]
  assign mmio_manager_io_in_wmask = {{8'd0}, stage1_out_bits_wmask}; // @[DCache.scala 241:14]
  assign mmio_manager_io_maxi_ar_ready = io_mmio_ar_ready; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_r_valid = io_mmio_r_valid; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_r_bits_data = io_mmio_r_bits_data; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_r_bits_last = io_mmio_r_bits_last; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_aw_ready = io_mmio_aw_ready; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_w_ready = io_mmio_w_ready; // @[DCache.scala 84:24]
  assign mmio_manager_io_maxi_b_valid = io_mmio_b_valid; // @[DCache.scala 84:24]
  assign mmio_manager_clint_rdata_0 = clint_rdata;
  always @(posedge clock) begin
    if (reset) begin // @[DCache.scala 65:37]
      curr_state <= 4'h0; // @[DCache.scala 65:37]
    end else if (_T_26) begin // @[Conditional.scala 40:58]
      if (io_prev_bits_flush) begin // @[DCache.scala 357:31]
        curr_state <= 4'h9; // @[DCache.scala 357:44]
      end else if (stage1_out_bits_data_id2mem_memory_rd_en | stage1_out_bits_data_id2mem_memory_we_en) begin // @[DCache.scala 358:45]
        curr_state <= _GEN_3549;
      end
    end else if (_T_29) begin // @[Conditional.scala 39:67]
      curr_state <= 4'h6; // @[DCache.scala 369:27]
    end else if (_T_30) begin // @[Conditional.scala 39:67]
      curr_state <= _GEN_3552;
    end else begin
      curr_state <= _GEN_3573;
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_addr <= 39'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_addr <= io_prev_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_63 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_63 <= _GEN_575;
      end else if (6'h3f == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_63 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_63 <= _GEN_1294;
      end else begin
        lru_list_63 <= _GEN_1294;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_63 <= _GEN_2009;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_62 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_62 <= _GEN_574;
      end else if (6'h3e == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_62 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_62 <= _GEN_1293;
      end else begin
        lru_list_62 <= _GEN_1293;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_62 <= _GEN_2008;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_61 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_61 <= _GEN_573;
      end else if (6'h3d == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_61 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_61 <= _GEN_1292;
      end else begin
        lru_list_61 <= _GEN_1292;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_61 <= _GEN_2007;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_60 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_60 <= _GEN_572;
      end else if (6'h3c == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_60 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_60 <= _GEN_1291;
      end else begin
        lru_list_60 <= _GEN_1291;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_60 <= _GEN_2006;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_59 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_59 <= _GEN_571;
      end else if (6'h3b == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_59 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_59 <= _GEN_1290;
      end else begin
        lru_list_59 <= _GEN_1290;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_59 <= _GEN_2005;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_58 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_58 <= _GEN_570;
      end else if (6'h3a == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_58 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_58 <= _GEN_1289;
      end else begin
        lru_list_58 <= _GEN_1289;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_58 <= _GEN_2004;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_57 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_57 <= _GEN_569;
      end else if (6'h39 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_57 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_57 <= _GEN_1288;
      end else begin
        lru_list_57 <= _GEN_1288;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_57 <= _GEN_2003;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_56 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_56 <= _GEN_568;
      end else if (6'h38 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_56 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_56 <= _GEN_1287;
      end else begin
        lru_list_56 <= _GEN_1287;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_56 <= _GEN_2002;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_55 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_55 <= _GEN_567;
      end else if (6'h37 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_55 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_55 <= _GEN_1286;
      end else begin
        lru_list_55 <= _GEN_1286;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_55 <= _GEN_2001;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_54 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_54 <= _GEN_566;
      end else if (6'h36 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_54 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_54 <= _GEN_1285;
      end else begin
        lru_list_54 <= _GEN_1285;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_54 <= _GEN_2000;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_53 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_53 <= _GEN_565;
      end else if (6'h35 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_53 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_53 <= _GEN_1284;
      end else begin
        lru_list_53 <= _GEN_1284;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_53 <= _GEN_1999;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_52 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_52 <= _GEN_564;
      end else if (6'h34 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_52 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_52 <= _GEN_1283;
      end else begin
        lru_list_52 <= _GEN_1283;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_52 <= _GEN_1998;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_51 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_51 <= _GEN_563;
      end else if (6'h33 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_51 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_51 <= _GEN_1282;
      end else begin
        lru_list_51 <= _GEN_1282;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_51 <= _GEN_1997;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_50 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_50 <= _GEN_562;
      end else if (6'h32 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_50 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_50 <= _GEN_1281;
      end else begin
        lru_list_50 <= _GEN_1281;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_50 <= _GEN_1996;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_49 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_49 <= _GEN_561;
      end else if (6'h31 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_49 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_49 <= _GEN_1280;
      end else begin
        lru_list_49 <= _GEN_1280;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_49 <= _GEN_1995;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_48 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_48 <= _GEN_560;
      end else if (6'h30 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_48 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_48 <= _GEN_1279;
      end else begin
        lru_list_48 <= _GEN_1279;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_48 <= _GEN_1994;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_47 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_47 <= _GEN_559;
      end else if (6'h2f == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_47 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_47 <= _GEN_1278;
      end else begin
        lru_list_47 <= _GEN_1278;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_47 <= _GEN_1993;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_46 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_46 <= _GEN_558;
      end else if (6'h2e == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_46 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_46 <= _GEN_1277;
      end else begin
        lru_list_46 <= _GEN_1277;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_46 <= _GEN_1992;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_45 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_45 <= _GEN_557;
      end else if (6'h2d == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_45 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_45 <= _GEN_1276;
      end else begin
        lru_list_45 <= _GEN_1276;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_45 <= _GEN_1991;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_44 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_44 <= _GEN_556;
      end else if (6'h2c == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_44 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_44 <= _GEN_1275;
      end else begin
        lru_list_44 <= _GEN_1275;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_44 <= _GEN_1990;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_43 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_43 <= _GEN_555;
      end else if (6'h2b == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_43 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_43 <= _GEN_1274;
      end else begin
        lru_list_43 <= _GEN_1274;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_43 <= _GEN_1989;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_42 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_42 <= _GEN_554;
      end else if (6'h2a == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_42 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_42 <= _GEN_1273;
      end else begin
        lru_list_42 <= _GEN_1273;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_42 <= _GEN_1988;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_41 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_41 <= _GEN_553;
      end else if (6'h29 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_41 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_41 <= _GEN_1272;
      end else begin
        lru_list_41 <= _GEN_1272;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_41 <= _GEN_1987;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_40 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_40 <= _GEN_552;
      end else if (6'h28 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_40 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_40 <= _GEN_1271;
      end else begin
        lru_list_40 <= _GEN_1271;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_40 <= _GEN_1986;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_39 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_39 <= _GEN_551;
      end else if (6'h27 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_39 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_39 <= _GEN_1270;
      end else begin
        lru_list_39 <= _GEN_1270;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_39 <= _GEN_1985;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_38 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_38 <= _GEN_550;
      end else if (6'h26 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_38 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_38 <= _GEN_1269;
      end else begin
        lru_list_38 <= _GEN_1269;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_38 <= _GEN_1984;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_37 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_37 <= _GEN_549;
      end else if (6'h25 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_37 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_37 <= _GEN_1268;
      end else begin
        lru_list_37 <= _GEN_1268;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_37 <= _GEN_1983;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_36 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_36 <= _GEN_548;
      end else if (6'h24 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_36 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_36 <= _GEN_1267;
      end else begin
        lru_list_36 <= _GEN_1267;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_36 <= _GEN_1982;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_35 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_35 <= _GEN_547;
      end else if (6'h23 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_35 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_35 <= _GEN_1266;
      end else begin
        lru_list_35 <= _GEN_1266;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_35 <= _GEN_1981;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_34 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_34 <= _GEN_546;
      end else if (6'h22 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_34 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_34 <= _GEN_1265;
      end else begin
        lru_list_34 <= _GEN_1265;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_34 <= _GEN_1980;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_33 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_33 <= _GEN_545;
      end else if (6'h21 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_33 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_33 <= _GEN_1264;
      end else begin
        lru_list_33 <= _GEN_1264;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_33 <= _GEN_1979;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_32 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_32 <= _GEN_544;
      end else if (6'h20 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_32 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_32 <= _GEN_1263;
      end else begin
        lru_list_32 <= _GEN_1263;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_32 <= _GEN_1978;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_31 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_31 <= _GEN_543;
      end else if (6'h1f == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_31 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_31 <= _GEN_1262;
      end else begin
        lru_list_31 <= _GEN_1262;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_31 <= _GEN_1977;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_30 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_30 <= _GEN_542;
      end else if (6'h1e == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_30 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_30 <= _GEN_1261;
      end else begin
        lru_list_30 <= _GEN_1261;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_30 <= _GEN_1976;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_29 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_29 <= _GEN_541;
      end else if (6'h1d == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_29 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_29 <= _GEN_1260;
      end else begin
        lru_list_29 <= _GEN_1260;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_29 <= _GEN_1975;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_28 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_28 <= _GEN_540;
      end else if (6'h1c == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_28 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_28 <= _GEN_1259;
      end else begin
        lru_list_28 <= _GEN_1259;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_28 <= _GEN_1974;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_27 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_27 <= _GEN_539;
      end else if (6'h1b == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_27 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_27 <= _GEN_1258;
      end else begin
        lru_list_27 <= _GEN_1258;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_27 <= _GEN_1973;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_26 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_26 <= _GEN_538;
      end else if (6'h1a == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_26 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_26 <= _GEN_1257;
      end else begin
        lru_list_26 <= _GEN_1257;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_26 <= _GEN_1972;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_25 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_25 <= _GEN_537;
      end else if (6'h19 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_25 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_25 <= _GEN_1256;
      end else begin
        lru_list_25 <= _GEN_1256;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_25 <= _GEN_1971;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_24 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_24 <= _GEN_536;
      end else if (6'h18 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_24 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_24 <= _GEN_1255;
      end else begin
        lru_list_24 <= _GEN_1255;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_24 <= _GEN_1970;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_23 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_23 <= _GEN_535;
      end else if (6'h17 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_23 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_23 <= _GEN_1254;
      end else begin
        lru_list_23 <= _GEN_1254;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_23 <= _GEN_1969;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_22 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_22 <= _GEN_534;
      end else if (6'h16 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_22 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_22 <= _GEN_1253;
      end else begin
        lru_list_22 <= _GEN_1253;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_22 <= _GEN_1968;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_21 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_21 <= _GEN_533;
      end else if (6'h15 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_21 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_21 <= _GEN_1252;
      end else begin
        lru_list_21 <= _GEN_1252;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_21 <= _GEN_1967;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_20 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_20 <= _GEN_532;
      end else if (6'h14 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_20 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_20 <= _GEN_1251;
      end else begin
        lru_list_20 <= _GEN_1251;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_20 <= _GEN_1966;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_19 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_19 <= _GEN_531;
      end else if (6'h13 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_19 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_19 <= _GEN_1250;
      end else begin
        lru_list_19 <= _GEN_1250;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_19 <= _GEN_1965;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_18 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_18 <= _GEN_530;
      end else if (6'h12 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_18 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_18 <= _GEN_1249;
      end else begin
        lru_list_18 <= _GEN_1249;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_18 <= _GEN_1964;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_17 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_17 <= _GEN_529;
      end else if (6'h11 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_17 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_17 <= _GEN_1248;
      end else begin
        lru_list_17 <= _GEN_1248;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_17 <= _GEN_1963;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_16 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_16 <= _GEN_528;
      end else if (6'h10 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_16 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_16 <= _GEN_1247;
      end else begin
        lru_list_16 <= _GEN_1247;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_16 <= _GEN_1962;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_15 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_15 <= _GEN_527;
      end else if (6'hf == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_15 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_15 <= _GEN_1246;
      end else begin
        lru_list_15 <= _GEN_1246;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_15 <= _GEN_1961;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_14 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_14 <= _GEN_526;
      end else if (6'he == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_14 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_14 <= _GEN_1245;
      end else begin
        lru_list_14 <= _GEN_1245;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_14 <= _GEN_1960;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_13 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_13 <= _GEN_525;
      end else if (6'hd == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_13 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_13 <= _GEN_1244;
      end else begin
        lru_list_13 <= _GEN_1244;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_13 <= _GEN_1959;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_12 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_12 <= _GEN_524;
      end else if (6'hc == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_12 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_12 <= _GEN_1243;
      end else begin
        lru_list_12 <= _GEN_1243;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_12 <= _GEN_1958;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_11 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_11 <= _GEN_523;
      end else if (6'hb == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_11 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_11 <= _GEN_1242;
      end else begin
        lru_list_11 <= _GEN_1242;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_11 <= _GEN_1957;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_10 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_10 <= _GEN_522;
      end else if (6'ha == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_10 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_10 <= _GEN_1241;
      end else begin
        lru_list_10 <= _GEN_1241;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_10 <= _GEN_1956;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_9 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_9 <= _GEN_521;
      end else if (6'h9 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_9 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_9 <= _GEN_1240;
      end else begin
        lru_list_9 <= _GEN_1240;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_9 <= _GEN_1955;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_8 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_8 <= _GEN_520;
      end else if (6'h8 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_8 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_8 <= _GEN_1239;
      end else begin
        lru_list_8 <= _GEN_1239;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_8 <= _GEN_1954;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_7 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_7 <= _GEN_519;
      end else if (6'h7 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_7 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_7 <= _GEN_1238;
      end else begin
        lru_list_7 <= _GEN_1238;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_7 <= _GEN_1953;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_6 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_6 <= _GEN_518;
      end else if (6'h6 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_6 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_6 <= _GEN_1237;
      end else begin
        lru_list_6 <= _GEN_1237;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_6 <= _GEN_1952;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_5 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_5 <= _GEN_517;
      end else if (6'h5 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_5 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_5 <= _GEN_1236;
      end else begin
        lru_list_5 <= _GEN_1236;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_5 <= _GEN_1951;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_4 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_4 <= _GEN_516;
      end else if (6'h4 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_4 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_4 <= _GEN_1235;
      end else begin
        lru_list_4 <= _GEN_1235;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_4 <= _GEN_1950;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_3 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_3 <= _GEN_515;
      end else if (6'h3 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_3 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_3 <= _GEN_1234;
      end else begin
        lru_list_3 <= _GEN_1234;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_3 <= _GEN_1949;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_2 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_2 <= _GEN_514;
      end else if (6'h2 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_2 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_2 <= _GEN_1233;
      end else begin
        lru_list_2 <= _GEN_1233;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_2 <= _GEN_1948;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_1 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_1 <= _GEN_513;
      end else if (6'h1 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_1 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_1 <= _GEN_1232;
      end else begin
        lru_list_1 <= _GEN_1232;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_1 <= _GEN_1947;
    end
    if (reset) begin // @[DCache.scala 118:35]
      lru_list_0 <= 1'h0; // @[DCache.scala 118:35]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        lru_list_0 <= _GEN_512;
      end else if (6'h0 == stage1_index) begin // @[DCache.scala 278:32]
        lru_list_0 <= 1'h0; // @[DCache.scala 278:32]
      end
    end else if (curr_state == 4'hb) begin // @[DCache.scala 286:38]
      if (flush_way) begin // @[DCache.scala 287:22]
        lru_list_0 <= _GEN_1231;
      end else begin
        lru_list_0 <= _GEN_1231;
      end
    end else if (curr_state == 4'h1) begin // @[DCache.scala 297:36]
      lru_list_0 <= _GEN_1946;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 7'h0; // @[Counter.scala 60:40]
    end else if (flush_cnt_rst) begin // @[DCache.scala 144:23]
      value <= 7'h0; // @[Counter.scala 97:11]
    end else if (flush_cnt_en) begin // @[DCache.scala 132:23]
      value <= _flush_cnt_end_latch_en_value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Reg.scala 27:20]
      hit_reg <= 1'h0; // @[Reg.scala 27:20]
    end else if (hit_reg_x8) begin // @[Reg.scala 28:19]
      hit_reg <= tag1_hit; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_0 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_0 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_0 <= _GEN_832;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_0 <= _GEN_2417;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_1 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_1 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_1 <= _GEN_833;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_1 <= _GEN_2418;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_2 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_2 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_2 <= _GEN_834;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_2 <= _GEN_2419;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_3 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_3 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_3 <= _GEN_835;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_3 <= _GEN_2420;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_4 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_4 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_4 <= _GEN_836;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_4 <= _GEN_2421;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_5 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_5 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_5 <= _GEN_837;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_5 <= _GEN_2422;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_6 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_6 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_6 <= _GEN_838;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_6 <= _GEN_2423;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_7 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_7 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_7 <= _GEN_839;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_7 <= _GEN_2424;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_8 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_8 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_8 <= _GEN_840;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_8 <= _GEN_2425;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_9 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_9 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_9 <= _GEN_841;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_9 <= _GEN_2426;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_10 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_10 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_10 <= _GEN_842;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_10 <= _GEN_2427;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_11 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_11 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_11 <= _GEN_843;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_11 <= _GEN_2428;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_12 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_12 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_12 <= _GEN_844;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_12 <= _GEN_2429;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_13 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_13 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_13 <= _GEN_845;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_13 <= _GEN_2430;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_14 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_14 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_14 <= _GEN_846;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_14 <= _GEN_2431;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_15 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_15 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_15 <= _GEN_847;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_15 <= _GEN_2432;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_16 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_16 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_16 <= _GEN_848;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_16 <= _GEN_2433;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_17 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_17 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_17 <= _GEN_849;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_17 <= _GEN_2434;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_18 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_18 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_18 <= _GEN_850;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_18 <= _GEN_2435;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_19 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_19 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_19 <= _GEN_851;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_19 <= _GEN_2436;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_20 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_20 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_20 <= _GEN_852;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_20 <= _GEN_2437;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_21 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_21 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_21 <= _GEN_853;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_21 <= _GEN_2438;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_22 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_22 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_22 <= _GEN_854;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_22 <= _GEN_2439;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_23 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_23 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_23 <= _GEN_855;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_23 <= _GEN_2440;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_24 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_24 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_24 <= _GEN_856;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_24 <= _GEN_2441;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_25 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_25 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_25 <= _GEN_857;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_25 <= _GEN_2442;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_26 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_26 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_26 <= _GEN_858;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_26 <= _GEN_2443;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_27 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_27 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_27 <= _GEN_859;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_27 <= _GEN_2444;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_28 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_28 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_28 <= _GEN_860;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_28 <= _GEN_2445;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_29 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_29 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_29 <= _GEN_861;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_29 <= _GEN_2446;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_30 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_30 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_30 <= _GEN_862;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_30 <= _GEN_2447;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_31 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_31 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_31 <= _GEN_863;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_31 <= _GEN_2448;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_32 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_32 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_32 <= _GEN_864;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_32 <= _GEN_2449;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_33 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_33 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_33 <= _GEN_865;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_33 <= _GEN_2450;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_34 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_34 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_34 <= _GEN_866;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_34 <= _GEN_2451;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_35 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_35 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_35 <= _GEN_867;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_35 <= _GEN_2452;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_36 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_36 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_36 <= _GEN_868;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_36 <= _GEN_2453;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_37 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_37 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_37 <= _GEN_869;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_37 <= _GEN_2454;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_38 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_38 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_38 <= _GEN_870;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_38 <= _GEN_2455;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_39 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_39 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_39 <= _GEN_871;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_39 <= _GEN_2456;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_40 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_40 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_40 <= _GEN_872;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_40 <= _GEN_2457;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_41 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_41 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_41 <= _GEN_873;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_41 <= _GEN_2458;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_42 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_42 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_42 <= _GEN_874;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_42 <= _GEN_2459;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_43 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_43 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_43 <= _GEN_875;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_43 <= _GEN_2460;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_44 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_44 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_44 <= _GEN_876;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_44 <= _GEN_2461;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_45 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_45 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_45 <= _GEN_877;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_45 <= _GEN_2462;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_46 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_46 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_46 <= _GEN_878;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_46 <= _GEN_2463;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_47 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_47 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_47 <= _GEN_879;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_47 <= _GEN_2464;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_48 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_48 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_48 <= _GEN_880;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_48 <= _GEN_2465;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_49 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_49 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_49 <= _GEN_881;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_49 <= _GEN_2466;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_50 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_50 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_50 <= _GEN_882;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_50 <= _GEN_2467;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_51 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_51 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_51 <= _GEN_883;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_51 <= _GEN_2468;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_52 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_52 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_52 <= _GEN_884;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_52 <= _GEN_2469;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_53 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_53 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_53 <= _GEN_885;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_53 <= _GEN_2470;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_54 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_54 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_54 <= _GEN_886;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_54 <= _GEN_2471;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_55 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_55 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_55 <= _GEN_887;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_55 <= _GEN_2472;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_56 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_56 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_56 <= _GEN_888;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_56 <= _GEN_2473;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_57 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_57 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_57 <= _GEN_889;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_57 <= _GEN_2474;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_58 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_58 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_58 <= _GEN_890;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_58 <= _GEN_2475;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_59 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_59 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_59 <= _GEN_891;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_59 <= _GEN_2476;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_60 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_60 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_60 <= _GEN_892;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_60 <= _GEN_2477;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_61 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_61 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_61 <= _GEN_893;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_61 <= _GEN_2478;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_62 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_62 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_62 <= _GEN_894;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_62 <= _GEN_2479;
    end
    if (reset) begin // @[DCache.scala 113:44]
      dirty_array_0_63 <= 1'h0; // @[DCache.scala 113:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_0_63 <= 1'h0; // @[DCache.scala 319:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        dirty_array_0_63 <= _GEN_895;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_0_63 <= _GEN_2480;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_0 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_0 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_0 <= _GEN_640;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_0 <= _GEN_2552;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_1 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_1 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_1 <= _GEN_641;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_1 <= _GEN_2553;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_2 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_2 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_2 <= _GEN_642;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_2 <= _GEN_2554;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_3 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_3 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_3 <= _GEN_643;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_3 <= _GEN_2555;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_4 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_4 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_4 <= _GEN_644;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_4 <= _GEN_2556;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_5 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_5 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_5 <= _GEN_645;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_5 <= _GEN_2557;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_6 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_6 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_6 <= _GEN_646;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_6 <= _GEN_2558;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_7 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_7 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_7 <= _GEN_647;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_7 <= _GEN_2559;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_8 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_8 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_8 <= _GEN_648;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_8 <= _GEN_2560;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_9 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_9 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_9 <= _GEN_649;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_9 <= _GEN_2561;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_10 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_10 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_10 <= _GEN_650;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_10 <= _GEN_2562;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_11 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_11 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_11 <= _GEN_651;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_11 <= _GEN_2563;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_12 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_12 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_12 <= _GEN_652;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_12 <= _GEN_2564;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_13 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_13 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_13 <= _GEN_653;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_13 <= _GEN_2565;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_14 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_14 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_14 <= _GEN_654;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_14 <= _GEN_2566;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_15 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_15 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_15 <= _GEN_655;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_15 <= _GEN_2567;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_16 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_16 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_16 <= _GEN_656;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_16 <= _GEN_2568;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_17 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_17 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_17 <= _GEN_657;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_17 <= _GEN_2569;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_18 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_18 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_18 <= _GEN_658;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_18 <= _GEN_2570;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_19 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_19 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_19 <= _GEN_659;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_19 <= _GEN_2571;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_20 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_20 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_20 <= _GEN_660;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_20 <= _GEN_2572;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_21 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_21 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_21 <= _GEN_661;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_21 <= _GEN_2573;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_22 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_22 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_22 <= _GEN_662;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_22 <= _GEN_2574;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_23 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_23 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_23 <= _GEN_663;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_23 <= _GEN_2575;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_24 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_24 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_24 <= _GEN_664;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_24 <= _GEN_2576;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_25 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_25 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_25 <= _GEN_665;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_25 <= _GEN_2577;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_26 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_26 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_26 <= _GEN_666;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_26 <= _GEN_2578;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_27 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_27 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_27 <= _GEN_667;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_27 <= _GEN_2579;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_28 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_28 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_28 <= _GEN_668;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_28 <= _GEN_2580;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_29 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_29 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_29 <= _GEN_669;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_29 <= _GEN_2581;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_30 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_30 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_30 <= _GEN_670;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_30 <= _GEN_2582;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_31 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_31 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_31 <= _GEN_671;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_31 <= _GEN_2583;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_32 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_32 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_32 <= _GEN_672;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_32 <= _GEN_2584;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_33 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_33 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_33 <= _GEN_673;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_33 <= _GEN_2585;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_34 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_34 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_34 <= _GEN_674;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_34 <= _GEN_2586;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_35 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_35 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_35 <= _GEN_675;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_35 <= _GEN_2587;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_36 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_36 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_36 <= _GEN_676;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_36 <= _GEN_2588;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_37 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_37 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_37 <= _GEN_677;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_37 <= _GEN_2589;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_38 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_38 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_38 <= _GEN_678;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_38 <= _GEN_2590;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_39 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_39 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_39 <= _GEN_679;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_39 <= _GEN_2591;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_40 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_40 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_40 <= _GEN_680;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_40 <= _GEN_2592;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_41 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_41 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_41 <= _GEN_681;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_41 <= _GEN_2593;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_42 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_42 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_42 <= _GEN_682;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_42 <= _GEN_2594;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_43 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_43 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_43 <= _GEN_683;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_43 <= _GEN_2595;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_44 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_44 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_44 <= _GEN_684;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_44 <= _GEN_2596;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_45 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_45 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_45 <= _GEN_685;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_45 <= _GEN_2597;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_46 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_46 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_46 <= _GEN_686;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_46 <= _GEN_2598;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_47 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_47 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_47 <= _GEN_687;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_47 <= _GEN_2599;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_48 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_48 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_48 <= _GEN_688;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_48 <= _GEN_2600;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_49 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_49 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_49 <= _GEN_689;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_49 <= _GEN_2601;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_50 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_50 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_50 <= _GEN_690;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_50 <= _GEN_2602;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_51 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_51 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_51 <= _GEN_691;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_51 <= _GEN_2603;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_52 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_52 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_52 <= _GEN_692;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_52 <= _GEN_2604;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_53 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_53 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_53 <= _GEN_693;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_53 <= _GEN_2605;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_54 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_54 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_54 <= _GEN_694;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_54 <= _GEN_2606;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_55 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_55 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_55 <= _GEN_695;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_55 <= _GEN_2607;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_56 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_56 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_56 <= _GEN_696;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_56 <= _GEN_2608;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_57 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_57 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_57 <= _GEN_697;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_57 <= _GEN_2609;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_58 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_58 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_58 <= _GEN_698;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_58 <= _GEN_2610;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_59 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_59 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_59 <= _GEN_699;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_59 <= _GEN_2611;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_60 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_60 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_60 <= _GEN_700;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_60 <= _GEN_2612;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_61 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_61 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_61 <= _GEN_701;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_61 <= _GEN_2613;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_62 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_62 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_62 <= _GEN_702;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_62 <= _GEN_2614;
    end
    if (reset) begin // @[DCache.scala 114:44]
      dirty_array_1_63 <= 1'h0; // @[DCache.scala 114:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      dirty_array_1_63 <= 1'h0; // @[DCache.scala 317:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        dirty_array_1_63 <= _GEN_703;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      dirty_array_1_63 <= _GEN_2615;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_0 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_0 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_0 <= _GEN_768;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_0 <= _GEN_2353;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_1 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_1 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_1 <= _GEN_769;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_1 <= _GEN_2354;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_2 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_2 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_2 <= _GEN_770;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_2 <= _GEN_2355;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_3 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_3 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_3 <= _GEN_771;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_3 <= _GEN_2356;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_4 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_4 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_4 <= _GEN_772;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_4 <= _GEN_2357;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_5 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_5 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_5 <= _GEN_773;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_5 <= _GEN_2358;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_6 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_6 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_6 <= _GEN_774;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_6 <= _GEN_2359;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_7 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_7 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_7 <= _GEN_775;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_7 <= _GEN_2360;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_8 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_8 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_8 <= _GEN_776;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_8 <= _GEN_2361;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_9 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_9 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_9 <= _GEN_777;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_9 <= _GEN_2362;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_10 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_10 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_10 <= _GEN_778;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_10 <= _GEN_2363;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_11 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_11 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_11 <= _GEN_779;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_11 <= _GEN_2364;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_12 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_12 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_12 <= _GEN_780;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_12 <= _GEN_2365;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_13 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_13 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_13 <= _GEN_781;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_13 <= _GEN_2366;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_14 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_14 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_14 <= _GEN_782;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_14 <= _GEN_2367;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_15 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_15 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_15 <= _GEN_783;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_15 <= _GEN_2368;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_16 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_16 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_16 <= _GEN_784;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_16 <= _GEN_2369;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_17 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_17 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_17 <= _GEN_785;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_17 <= _GEN_2370;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_18 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_18 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_18 <= _GEN_786;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_18 <= _GEN_2371;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_19 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_19 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_19 <= _GEN_787;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_19 <= _GEN_2372;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_20 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_20 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_20 <= _GEN_788;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_20 <= _GEN_2373;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_21 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_21 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_21 <= _GEN_789;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_21 <= _GEN_2374;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_22 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_22 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_22 <= _GEN_790;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_22 <= _GEN_2375;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_23 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_23 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_23 <= _GEN_791;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_23 <= _GEN_2376;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_24 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_24 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_24 <= _GEN_792;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_24 <= _GEN_2377;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_25 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_25 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_25 <= _GEN_793;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_25 <= _GEN_2378;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_26 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_26 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_26 <= _GEN_794;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_26 <= _GEN_2379;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_27 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_27 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_27 <= _GEN_795;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_27 <= _GEN_2380;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_28 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_28 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_28 <= _GEN_796;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_28 <= _GEN_2381;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_29 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_29 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_29 <= _GEN_797;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_29 <= _GEN_2382;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_30 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_30 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_30 <= _GEN_798;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_30 <= _GEN_2383;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_31 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_31 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_31 <= _GEN_799;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_31 <= _GEN_2384;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_32 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_32 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_32 <= _GEN_800;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_32 <= _GEN_2385;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_33 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_33 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_33 <= _GEN_801;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_33 <= _GEN_2386;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_34 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_34 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_34 <= _GEN_802;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_34 <= _GEN_2387;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_35 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_35 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_35 <= _GEN_803;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_35 <= _GEN_2388;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_36 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_36 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_36 <= _GEN_804;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_36 <= _GEN_2389;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_37 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_37 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_37 <= _GEN_805;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_37 <= _GEN_2390;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_38 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_38 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_38 <= _GEN_806;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_38 <= _GEN_2391;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_39 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_39 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_39 <= _GEN_807;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_39 <= _GEN_2392;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_40 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_40 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_40 <= _GEN_808;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_40 <= _GEN_2393;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_41 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_41 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_41 <= _GEN_809;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_41 <= _GEN_2394;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_42 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_42 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_42 <= _GEN_810;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_42 <= _GEN_2395;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_43 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_43 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_43 <= _GEN_811;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_43 <= _GEN_2396;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_44 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_44 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_44 <= _GEN_812;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_44 <= _GEN_2397;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_45 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_45 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_45 <= _GEN_813;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_45 <= _GEN_2398;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_46 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_46 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_46 <= _GEN_814;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_46 <= _GEN_2399;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_47 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_47 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_47 <= _GEN_815;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_47 <= _GEN_2400;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_48 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_48 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_48 <= _GEN_816;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_48 <= _GEN_2401;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_49 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_49 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_49 <= _GEN_817;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_49 <= _GEN_2402;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_50 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_50 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_50 <= _GEN_818;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_50 <= _GEN_2403;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_51 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_51 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_51 <= _GEN_819;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_51 <= _GEN_2404;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_52 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_52 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_52 <= _GEN_820;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_52 <= _GEN_2405;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_53 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_53 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_53 <= _GEN_821;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_53 <= _GEN_2406;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_54 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_54 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_54 <= _GEN_822;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_54 <= _GEN_2407;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_55 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_55 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_55 <= _GEN_823;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_55 <= _GEN_2408;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_56 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_56 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_56 <= _GEN_824;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_56 <= _GEN_2409;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_57 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_57 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_57 <= _GEN_825;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_57 <= _GEN_2410;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_58 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_58 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_58 <= _GEN_826;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_58 <= _GEN_2411;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_59 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_59 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_59 <= _GEN_827;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_59 <= _GEN_2412;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_60 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_60 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_60 <= _GEN_828;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_60 <= _GEN_2413;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_61 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_61 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_61 <= _GEN_829;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_61 <= _GEN_2414;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_62 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_62 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_62 <= _GEN_830;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_62 <= _GEN_2415;
    end
    if (reset) begin // @[DCache.scala 115:44]
      valid_array_0_63 <= 1'h0; // @[DCache.scala 115:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_0_63 <= 1'h0; // @[DCache.scala 318:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (!(next_way)) begin // @[DCache.scala 270:19]
        valid_array_0_63 <= _GEN_831;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_0_63 <= _GEN_2416;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_0 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_0 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_0 <= _GEN_576;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_0 <= _GEN_2488;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_1 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_1 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_1 <= _GEN_577;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_1 <= _GEN_2489;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_2 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_2 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_2 <= _GEN_578;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_2 <= _GEN_2490;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_3 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_3 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_3 <= _GEN_579;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_3 <= _GEN_2491;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_4 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_4 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_4 <= _GEN_580;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_4 <= _GEN_2492;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_5 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_5 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_5 <= _GEN_581;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_5 <= _GEN_2493;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_6 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_6 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_6 <= _GEN_582;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_6 <= _GEN_2494;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_7 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_7 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_7 <= _GEN_583;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_7 <= _GEN_2495;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_8 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_8 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_8 <= _GEN_584;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_8 <= _GEN_2496;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_9 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_9 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_9 <= _GEN_585;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_9 <= _GEN_2497;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_10 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_10 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_10 <= _GEN_586;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_10 <= _GEN_2498;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_11 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_11 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_11 <= _GEN_587;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_11 <= _GEN_2499;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_12 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_12 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_12 <= _GEN_588;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_12 <= _GEN_2500;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_13 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_13 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_13 <= _GEN_589;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_13 <= _GEN_2501;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_14 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_14 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_14 <= _GEN_590;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_14 <= _GEN_2502;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_15 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_15 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_15 <= _GEN_591;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_15 <= _GEN_2503;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_16 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_16 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_16 <= _GEN_592;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_16 <= _GEN_2504;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_17 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_17 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_17 <= _GEN_593;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_17 <= _GEN_2505;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_18 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_18 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_18 <= _GEN_594;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_18 <= _GEN_2506;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_19 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_19 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_19 <= _GEN_595;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_19 <= _GEN_2507;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_20 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_20 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_20 <= _GEN_596;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_20 <= _GEN_2508;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_21 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_21 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_21 <= _GEN_597;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_21 <= _GEN_2509;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_22 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_22 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_22 <= _GEN_598;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_22 <= _GEN_2510;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_23 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_23 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_23 <= _GEN_599;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_23 <= _GEN_2511;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_24 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_24 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_24 <= _GEN_600;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_24 <= _GEN_2512;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_25 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_25 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_25 <= _GEN_601;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_25 <= _GEN_2513;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_26 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_26 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_26 <= _GEN_602;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_26 <= _GEN_2514;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_27 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_27 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_27 <= _GEN_603;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_27 <= _GEN_2515;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_28 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_28 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_28 <= _GEN_604;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_28 <= _GEN_2516;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_29 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_29 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_29 <= _GEN_605;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_29 <= _GEN_2517;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_30 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_30 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_30 <= _GEN_606;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_30 <= _GEN_2518;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_31 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_31 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_31 <= _GEN_607;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_31 <= _GEN_2519;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_32 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_32 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_32 <= _GEN_608;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_32 <= _GEN_2520;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_33 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_33 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_33 <= _GEN_609;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_33 <= _GEN_2521;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_34 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_34 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_34 <= _GEN_610;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_34 <= _GEN_2522;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_35 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_35 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_35 <= _GEN_611;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_35 <= _GEN_2523;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_36 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_36 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_36 <= _GEN_612;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_36 <= _GEN_2524;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_37 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_37 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_37 <= _GEN_613;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_37 <= _GEN_2525;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_38 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_38 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_38 <= _GEN_614;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_38 <= _GEN_2526;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_39 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_39 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_39 <= _GEN_615;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_39 <= _GEN_2527;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_40 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_40 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_40 <= _GEN_616;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_40 <= _GEN_2528;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_41 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_41 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_41 <= _GEN_617;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_41 <= _GEN_2529;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_42 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_42 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_42 <= _GEN_618;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_42 <= _GEN_2530;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_43 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_43 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_43 <= _GEN_619;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_43 <= _GEN_2531;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_44 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_44 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_44 <= _GEN_620;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_44 <= _GEN_2532;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_45 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_45 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_45 <= _GEN_621;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_45 <= _GEN_2533;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_46 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_46 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_46 <= _GEN_622;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_46 <= _GEN_2534;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_47 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_47 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_47 <= _GEN_623;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_47 <= _GEN_2535;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_48 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_48 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_48 <= _GEN_624;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_48 <= _GEN_2536;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_49 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_49 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_49 <= _GEN_625;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_49 <= _GEN_2537;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_50 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_50 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_50 <= _GEN_626;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_50 <= _GEN_2538;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_51 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_51 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_51 <= _GEN_627;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_51 <= _GEN_2539;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_52 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_52 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_52 <= _GEN_628;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_52 <= _GEN_2540;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_53 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_53 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_53 <= _GEN_629;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_53 <= _GEN_2541;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_54 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_54 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_54 <= _GEN_630;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_54 <= _GEN_2542;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_55 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_55 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_55 <= _GEN_631;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_55 <= _GEN_2543;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_56 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_56 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_56 <= _GEN_632;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_56 <= _GEN_2544;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_57 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_57 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_57 <= _GEN_633;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_57 <= _GEN_2545;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_58 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_58 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_58 <= _GEN_634;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_58 <= _GEN_2546;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_59 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_59 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_59 <= _GEN_635;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_59 <= _GEN_2547;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_60 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_60 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_60 <= _GEN_636;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_60 <= _GEN_2548;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_61 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_61 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_61 <= _GEN_637;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_61 <= _GEN_2549;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_62 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_62 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_62 <= _GEN_638;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_62 <= _GEN_2550;
    end
    if (reset) begin // @[DCache.scala 116:44]
      valid_array_1_63 <= 1'h0; // @[DCache.scala 116:44]
    end else if (_T_13 & flush_way & flush_index == 6'h3f) begin // @[DCache.scala 315:84]
      valid_array_1_63 <= 1'h0; // @[DCache.scala 316:19]
    end else if (curr_state == 4'h2 & maxi4_manager_io_out_finish) begin // @[DCache.scala 269:43]
      if (next_way) begin // @[DCache.scala 270:19]
        valid_array_1_63 <= _GEN_639;
      end
    end else if (!(curr_state == 4'hb)) begin // @[DCache.scala 286:38]
      valid_array_1_63 <= _GEN_2551;
    end
    if (reset) begin // @[DCache.scala 122:40]
      flush_skip <= 1'h0; // @[DCache.scala 122:40]
    end else if (curr_state == 4'h9) begin // @[DCache.scala 247:30]
      flush_skip <= _GEN_509;
    end
    if (reset) begin // @[DCache.scala 125:49]
      flush_cnt_end_latch_en <= 1'h0; // @[DCache.scala 125:49]
    end else if (flush_cnt_en) begin // @[DCache.scala 132:23]
      flush_cnt_end_latch_en <= flush_cnt_end_latch_en_wrap; // @[DCache.scala 133:28]
    end else if (flush_cnt_rst) begin // @[DCache.scala 134:28]
      flush_cnt_end_latch_en <= 1'h0; // @[DCache.scala 135:28]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_valid <= io_prev_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2mem_sext_flag <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2mem_sext_flag <= io_prev_bits_data_id2mem_sext_flag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2mem_memory_rd_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2mem_memory_rd_en <= io_prev_bits_data_id2mem_memory_rd_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2mem_memory_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2mem_memory_we_en <= io_prev_bits_data_id2mem_memory_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2wb_intr_exce_ret <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2wb_intr_exce_ret <= io_prev_bits_data_id2wb_intr_exce_ret; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2wb_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2wb_fencei <= io_prev_bits_data_id2wb_fencei; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2wb_wb_sel <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2wb_wb_sel <= io_prev_bits_data_id2wb_wb_sel; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2wb_regfile_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2wb_regfile_we_en <= io_prev_bits_data_id2wb_regfile_we_en; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_id2wb_regfile_we_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_id2wb_regfile_we_addr <= io_prev_bits_data_id2wb_regfile_we_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_ex2mem_we_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_ex2mem_we_data <= io_prev_bits_data_ex2mem_we_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_data_ex2wb_result_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_data_ex2wb_result_data <= io_prev_bits_data_ex2wb_result_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_wdata <= io_prev_bits_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_wmask <= io_prev_bits_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_size_byte <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_size_byte <= io_prev_bits_size_byte; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_size_hword <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_size_hword <= io_prev_bits_size_hword; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_size_word <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_size_word <= io_prev_bits_size_word; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stage1_out_bits_size_dword <= 1'h0; // @[Reg.scala 27:20]
    end else if (go_on) begin // @[Reg.scala 28:19]
      stage1_out_bits_size_dword <= io_prev_bits_size_dword; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[3:0];
  _RAND_1 = {2{`RANDOM}};
  stage1_out_bits_addr = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  lru_list_63 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_list_62 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_list_61 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_list_60 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_list_59 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_list_58 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_list_57 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_list_56 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_list_55 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_list_54 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_list_53 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_list_52 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_list_51 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_list_50 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_list_49 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_list_48 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_list_47 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_list_46 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_list_45 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_list_44 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_list_43 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_list_42 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_list_41 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_list_40 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_list_39 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_list_38 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_list_37 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_list_36 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_list_35 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_list_34 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_list_33 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_list_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_list_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_list_30 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_list_29 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_list_28 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_list_27 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_list_26 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_list_25 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_list_24 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_list_23 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_list_22 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_list_21 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_list_20 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_list_19 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_list_18 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_list_17 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_list_16 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_list_15 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_list_14 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_list_13 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_list_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_list_11 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_list_10 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_list_9 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_list_8 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_list_7 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_list_6 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_list_5 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_list_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_list_3 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_list_2 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_list_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_list_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  value = _RAND_66[6:0];
  _RAND_67 = {1{`RANDOM}};
  hit_reg = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dirty_array_0_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dirty_array_0_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dirty_array_0_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dirty_array_0_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dirty_array_0_4 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dirty_array_0_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dirty_array_0_6 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dirty_array_0_7 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dirty_array_0_8 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dirty_array_0_9 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dirty_array_0_10 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dirty_array_0_11 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dirty_array_0_12 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dirty_array_0_13 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dirty_array_0_14 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dirty_array_0_15 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dirty_array_0_16 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dirty_array_0_17 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dirty_array_0_18 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dirty_array_0_19 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dirty_array_0_20 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dirty_array_0_21 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dirty_array_0_22 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dirty_array_0_23 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dirty_array_0_24 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dirty_array_0_25 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dirty_array_0_26 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dirty_array_0_27 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_array_0_28 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_array_0_29 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_array_0_30 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_array_0_31 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_array_0_32 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_array_0_33 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_array_0_34 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_array_0_35 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_array_0_36 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_array_0_37 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_array_0_38 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_array_0_39 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_array_0_40 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_array_0_41 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_array_0_42 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_array_0_43 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_array_0_44 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_array_0_45 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_array_0_46 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_array_0_47 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_array_0_48 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_array_0_49 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_array_0_50 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_array_0_51 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_array_0_52 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_array_0_53 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_array_0_54 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_array_0_55 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_array_0_56 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_array_0_57 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_array_0_58 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_array_0_59 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_array_0_60 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_array_0_61 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_array_0_62 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  dirty_array_0_63 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  dirty_array_1_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  dirty_array_1_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  dirty_array_1_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  dirty_array_1_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dirty_array_1_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  dirty_array_1_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  dirty_array_1_6 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  dirty_array_1_7 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dirty_array_1_8 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  dirty_array_1_9 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  dirty_array_1_10 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  dirty_array_1_11 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dirty_array_1_12 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  dirty_array_1_13 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  dirty_array_1_14 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  dirty_array_1_15 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dirty_array_1_16 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  dirty_array_1_17 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  dirty_array_1_18 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  dirty_array_1_19 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dirty_array_1_20 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dirty_array_1_21 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dirty_array_1_22 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dirty_array_1_23 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dirty_array_1_24 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dirty_array_1_25 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dirty_array_1_26 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dirty_array_1_27 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dirty_array_1_28 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dirty_array_1_29 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dirty_array_1_30 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dirty_array_1_31 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dirty_array_1_32 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dirty_array_1_33 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dirty_array_1_34 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dirty_array_1_35 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dirty_array_1_36 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dirty_array_1_37 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dirty_array_1_38 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dirty_array_1_39 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dirty_array_1_40 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dirty_array_1_41 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dirty_array_1_42 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dirty_array_1_43 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dirty_array_1_44 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dirty_array_1_45 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dirty_array_1_46 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dirty_array_1_47 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dirty_array_1_48 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dirty_array_1_49 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dirty_array_1_50 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dirty_array_1_51 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dirty_array_1_52 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dirty_array_1_53 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dirty_array_1_54 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dirty_array_1_55 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dirty_array_1_56 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dirty_array_1_57 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dirty_array_1_58 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dirty_array_1_59 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dirty_array_1_60 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dirty_array_1_61 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dirty_array_1_62 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dirty_array_1_63 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_array_0_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_array_0_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_array_0_2 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_array_0_3 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_array_0_4 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_array_0_5 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_array_0_6 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_array_0_7 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_array_0_8 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_array_0_9 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_array_0_10 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_array_0_11 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_array_0_12 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_array_0_13 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_array_0_14 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_array_0_15 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_array_0_16 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_array_0_17 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_array_0_18 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_array_0_19 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_array_0_20 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_array_0_21 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_array_0_22 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_array_0_23 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_array_0_24 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_array_0_25 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_array_0_26 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_array_0_27 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_array_0_28 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_array_0_29 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_array_0_30 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_array_0_31 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_array_0_32 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_array_0_33 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_array_0_34 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_array_0_35 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_array_0_36 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_array_0_37 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_array_0_38 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_array_0_39 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_array_0_40 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_array_0_41 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_array_0_42 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_array_0_43 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_array_0_44 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_array_0_45 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_array_0_46 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_array_0_47 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_array_0_48 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_array_0_49 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_array_0_50 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_array_0_51 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_array_0_52 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_array_0_53 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_array_0_54 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_array_0_55 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_array_0_56 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_array_0_57 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_array_0_58 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_array_0_59 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_array_0_60 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_array_0_61 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_array_0_62 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_array_0_63 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_array_1_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_array_1_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_array_1_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_array_1_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_array_1_4 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_array_1_5 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_array_1_6 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_array_1_7 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_array_1_8 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_array_1_9 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_array_1_10 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_array_1_11 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_array_1_12 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_array_1_13 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_array_1_14 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_array_1_15 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_array_1_16 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_array_1_17 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_array_1_18 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_array_1_19 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_array_1_20 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_array_1_21 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_array_1_22 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_array_1_23 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_array_1_24 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_array_1_25 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_array_1_26 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_array_1_27 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_array_1_28 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_array_1_29 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_array_1_30 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_array_1_31 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_array_1_32 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_array_1_33 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_array_1_34 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_array_1_35 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_array_1_36 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_array_1_37 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_array_1_38 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_array_1_39 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_array_1_40 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_array_1_41 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_array_1_42 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_array_1_43 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_array_1_44 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_array_1_45 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_array_1_46 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_array_1_47 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_array_1_48 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_array_1_49 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_array_1_50 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_array_1_51 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_array_1_52 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_array_1_53 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_array_1_54 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_array_1_55 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_array_1_56 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_array_1_57 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_array_1_58 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_array_1_59 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_array_1_60 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_array_1_61 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_array_1_62 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_array_1_63 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  flush_skip = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  flush_cnt_end_latch_en = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  stage1_out_valid = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  stage1_out_bits_data_id2mem_sext_flag = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  stage1_out_bits_data_id2mem_memory_rd_en = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  stage1_out_bits_data_id2mem_memory_we_en = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  stage1_out_bits_data_id2wb_intr_exce_ret = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  stage1_out_bits_data_id2wb_fencei = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  stage1_out_bits_data_id2wb_wb_sel = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  stage1_out_bits_data_id2wb_regfile_we_en = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  stage1_out_bits_data_id2wb_regfile_we_addr = _RAND_334[4:0];
  _RAND_335 = {2{`RANDOM}};
  stage1_out_bits_data_ex2mem_we_data = _RAND_335[63:0];
  _RAND_336 = {2{`RANDOM}};
  stage1_out_bits_data_ex2wb_result_data = _RAND_336[63:0];
  _RAND_337 = {2{`RANDOM}};
  stage1_out_bits_wdata = _RAND_337[63:0];
  _RAND_338 = {1{`RANDOM}};
  stage1_out_bits_wmask = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  stage1_out_bits_size_byte = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  stage1_out_bits_size_hword = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  stage1_out_bits_size_word = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  stage1_out_bits_size_dword = _RAND_342[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_MEMU(
  input          clock,
  input          reset,
  output         io_prev_ready,
  input          io_prev_valid,
  input          io_prev_bits_id2mem_fencei,
  input          io_prev_bits_id2mem_size_byte,
  input          io_prev_bits_id2mem_size_hword,
  input          io_prev_bits_id2mem_size_word,
  input          io_prev_bits_id2mem_size_dword,
  input          io_prev_bits_id2mem_sext_flag,
  input          io_prev_bits_id2mem_memory_rd_en,
  input          io_prev_bits_id2mem_memory_we_en,
  input          io_prev_bits_id2wb_intr_exce_ret,
  input          io_prev_bits_id2wb_fencei,
  input          io_prev_bits_id2wb_wb_sel,
  input          io_prev_bits_id2wb_regfile_we_en,
  input  [4:0]   io_prev_bits_id2wb_regfile_we_addr,
  input  [38:0]  io_prev_bits_ex2mem_addr,
  input  [63:0]  io_prev_bits_ex2mem_we_data,
  input  [7:0]   io_prev_bits_ex2mem_we_mask,
  input  [63:0]  io_prev_bits_ex2wb_result_data,
  output         io_next_valid,
  output         io_next_bits_id2wb_intr_exce_ret,
  output         io_next_bits_id2wb_fencei,
  output         io_next_bits_id2wb_wb_sel,
  output         io_next_bits_id2wb_regfile_we_en,
  output [4:0]   io_next_bits_id2wb_regfile_we_addr,
  output [63:0]  io_next_bits_ex2wb_result_data,
  output [63:0]  io_next_bits_mem2wb_memory_data,
  input          io_maxi_ar_ready,
  output         io_maxi_ar_valid,
  output [31:0]  io_maxi_ar_bits_addr,
  output [7:0]   io_maxi_ar_bits_len,
  output [2:0]   io_maxi_ar_bits_size,
  input          io_maxi_r_valid,
  input  [63:0]  io_maxi_r_bits_data,
  input          io_maxi_r_bits_last,
  input          io_maxi_aw_ready,
  output         io_maxi_aw_valid,
  output [31:0]  io_maxi_aw_bits_addr,
  output [7:0]   io_maxi_aw_bits_len,
  output [2:0]   io_maxi_aw_bits_size,
  input          io_maxi_w_ready,
  output         io_maxi_w_valid,
  output [63:0]  io_maxi_w_bits_data,
  output [7:0]   io_maxi_w_bits_strb,
  output         io_maxi_w_bits_last,
  input          io_maxi_b_valid,
  input          io_mmio_ar_ready,
  output         io_mmio_ar_valid,
  output [31:0]  io_mmio_ar_bits_addr,
  output [2:0]   io_mmio_ar_bits_size,
  input          io_mmio_r_valid,
  input  [63:0]  io_mmio_r_bits_data,
  input          io_mmio_r_bits_last,
  input          io_mmio_aw_ready,
  output         io_mmio_aw_valid,
  output [31:0]  io_mmio_aw_bits_addr,
  output [2:0]   io_mmio_aw_bits_size,
  input          io_mmio_w_ready,
  output         io_mmio_w_valid,
  output [63:0]  io_mmio_w_bits_data,
  output [7:0]   io_mmio_w_bits_strb,
  output         io_mmio_w_bits_last,
  input          io_mmio_b_valid,
  output [5:0]   io_sram4_addr,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,
  output         clint_we,
  output [31:0]  _T_24,
  input  [63:0]  clint_rdata,
  output [63:0]  clint_wdata
);
  wire  dcache_clock; // @[MEMU.scala 43:30]
  wire  dcache_reset; // @[MEMU.scala 43:30]
  wire  dcache_io_next_valid; // @[MEMU.scala 43:30]
  wire  dcache_io_next_bits_data_id2wb_intr_exce_ret; // @[MEMU.scala 43:30]
  wire  dcache_io_next_bits_data_id2wb_fencei; // @[MEMU.scala 43:30]
  wire  dcache_io_next_bits_data_id2wb_wb_sel; // @[MEMU.scala 43:30]
  wire  dcache_io_next_bits_data_id2wb_regfile_we_en; // @[MEMU.scala 43:30]
  wire [4:0] dcache_io_next_bits_data_id2wb_regfile_we_addr; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_next_bits_data_ex2wb_result_data; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_next_bits_data_mem2wb_memory_data; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_valid; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2mem_sext_flag; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2mem_memory_rd_en; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2mem_memory_we_en; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2wb_intr_exce_ret; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2wb_fencei; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2wb_wb_sel; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_data_id2wb_regfile_we_en; // @[MEMU.scala 43:30]
  wire [4:0] dcache_io_prev_bits_data_id2wb_regfile_we_addr; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_prev_bits_data_ex2mem_we_data; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_prev_bits_data_ex2wb_result_data; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_flush; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_prev_bits_wdata; // @[MEMU.scala 43:30]
  wire [7:0] dcache_io_prev_bits_wmask; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_size_byte; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_size_hword; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_size_word; // @[MEMU.scala 43:30]
  wire  dcache_io_prev_bits_size_dword; // @[MEMU.scala 43:30]
  wire [38:0] dcache_io_prev_bits_addr; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_ar_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_ar_valid; // @[MEMU.scala 43:30]
  wire [31:0] dcache_io_maxi_ar_bits_addr; // @[MEMU.scala 43:30]
  wire [7:0] dcache_io_maxi_ar_bits_len; // @[MEMU.scala 43:30]
  wire [2:0] dcache_io_maxi_ar_bits_size; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_r_valid; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_maxi_r_bits_data; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_r_bits_last; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_aw_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_aw_valid; // @[MEMU.scala 43:30]
  wire [31:0] dcache_io_maxi_aw_bits_addr; // @[MEMU.scala 43:30]
  wire [7:0] dcache_io_maxi_aw_bits_len; // @[MEMU.scala 43:30]
  wire [2:0] dcache_io_maxi_aw_bits_size; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_w_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_w_valid; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_maxi_w_bits_data; // @[MEMU.scala 43:30]
  wire [7:0] dcache_io_maxi_w_bits_strb; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_w_bits_last; // @[MEMU.scala 43:30]
  wire  dcache_io_maxi_b_valid; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_ar_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_ar_valid; // @[MEMU.scala 43:30]
  wire [31:0] dcache_io_mmio_ar_bits_addr; // @[MEMU.scala 43:30]
  wire [2:0] dcache_io_mmio_ar_bits_size; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_r_valid; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_mmio_r_bits_data; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_r_bits_last; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_aw_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_aw_valid; // @[MEMU.scala 43:30]
  wire [31:0] dcache_io_mmio_aw_bits_addr; // @[MEMU.scala 43:30]
  wire [2:0] dcache_io_mmio_aw_bits_size; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_w_ready; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_w_valid; // @[MEMU.scala 43:30]
  wire [63:0] dcache_io_mmio_w_bits_data; // @[MEMU.scala 43:30]
  wire [7:0] dcache_io_mmio_w_bits_strb; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_w_bits_last; // @[MEMU.scala 43:30]
  wire  dcache_io_mmio_b_valid; // @[MEMU.scala 43:30]
  wire [5:0] dcache_io_sram4_addr; // @[MEMU.scala 43:30]
  wire  dcache_io_sram4_wen; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram4_wmask; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram4_wdata; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram4_rdata; // @[MEMU.scala 43:30]
  wire [5:0] dcache_io_sram5_addr; // @[MEMU.scala 43:30]
  wire  dcache_io_sram5_wen; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram5_wmask; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram5_wdata; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram5_rdata; // @[MEMU.scala 43:30]
  wire [5:0] dcache_io_sram6_addr; // @[MEMU.scala 43:30]
  wire  dcache_io_sram6_wen; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram6_wmask; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram6_wdata; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram6_rdata; // @[MEMU.scala 43:30]
  wire [5:0] dcache_io_sram7_addr; // @[MEMU.scala 43:30]
  wire  dcache_io_sram7_wen; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram7_wmask; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram7_wdata; // @[MEMU.scala 43:30]
  wire [127:0] dcache_io_sram7_rdata; // @[MEMU.scala 43:30]
  wire  dcache_clint_we; // @[MEMU.scala 43:30]
  wire [31:0] dcache__T_24_0; // @[MEMU.scala 43:30]
  wire [63:0] dcache_clint_rdata; // @[MEMU.scala 43:30]
  wire [63:0] dcache_clint_wdata; // @[MEMU.scala 43:30]
  ysyx_040978_DCacheUnit dcache ( // @[MEMU.scala 43:30]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_next_valid(dcache_io_next_valid),
    .io_next_bits_data_id2wb_intr_exce_ret(dcache_io_next_bits_data_id2wb_intr_exce_ret),
    .io_next_bits_data_id2wb_fencei(dcache_io_next_bits_data_id2wb_fencei),
    .io_next_bits_data_id2wb_wb_sel(dcache_io_next_bits_data_id2wb_wb_sel),
    .io_next_bits_data_id2wb_regfile_we_en(dcache_io_next_bits_data_id2wb_regfile_we_en),
    .io_next_bits_data_id2wb_regfile_we_addr(dcache_io_next_bits_data_id2wb_regfile_we_addr),
    .io_next_bits_data_ex2wb_result_data(dcache_io_next_bits_data_ex2wb_result_data),
    .io_next_bits_data_mem2wb_memory_data(dcache_io_next_bits_data_mem2wb_memory_data),
    .io_prev_ready(dcache_io_prev_ready),
    .io_prev_valid(dcache_io_prev_valid),
    .io_prev_bits_data_id2mem_sext_flag(dcache_io_prev_bits_data_id2mem_sext_flag),
    .io_prev_bits_data_id2mem_memory_rd_en(dcache_io_prev_bits_data_id2mem_memory_rd_en),
    .io_prev_bits_data_id2mem_memory_we_en(dcache_io_prev_bits_data_id2mem_memory_we_en),
    .io_prev_bits_data_id2wb_intr_exce_ret(dcache_io_prev_bits_data_id2wb_intr_exce_ret),
    .io_prev_bits_data_id2wb_fencei(dcache_io_prev_bits_data_id2wb_fencei),
    .io_prev_bits_data_id2wb_wb_sel(dcache_io_prev_bits_data_id2wb_wb_sel),
    .io_prev_bits_data_id2wb_regfile_we_en(dcache_io_prev_bits_data_id2wb_regfile_we_en),
    .io_prev_bits_data_id2wb_regfile_we_addr(dcache_io_prev_bits_data_id2wb_regfile_we_addr),
    .io_prev_bits_data_ex2mem_we_data(dcache_io_prev_bits_data_ex2mem_we_data),
    .io_prev_bits_data_ex2wb_result_data(dcache_io_prev_bits_data_ex2wb_result_data),
    .io_prev_bits_flush(dcache_io_prev_bits_flush),
    .io_prev_bits_wdata(dcache_io_prev_bits_wdata),
    .io_prev_bits_wmask(dcache_io_prev_bits_wmask),
    .io_prev_bits_size_byte(dcache_io_prev_bits_size_byte),
    .io_prev_bits_size_hword(dcache_io_prev_bits_size_hword),
    .io_prev_bits_size_word(dcache_io_prev_bits_size_word),
    .io_prev_bits_size_dword(dcache_io_prev_bits_size_dword),
    .io_prev_bits_addr(dcache_io_prev_bits_addr),
    .io_maxi_ar_ready(dcache_io_maxi_ar_ready),
    .io_maxi_ar_valid(dcache_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(dcache_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(dcache_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(dcache_io_maxi_ar_bits_size),
    .io_maxi_r_valid(dcache_io_maxi_r_valid),
    .io_maxi_r_bits_data(dcache_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(dcache_io_maxi_r_bits_last),
    .io_maxi_aw_ready(dcache_io_maxi_aw_ready),
    .io_maxi_aw_valid(dcache_io_maxi_aw_valid),
    .io_maxi_aw_bits_addr(dcache_io_maxi_aw_bits_addr),
    .io_maxi_aw_bits_len(dcache_io_maxi_aw_bits_len),
    .io_maxi_aw_bits_size(dcache_io_maxi_aw_bits_size),
    .io_maxi_w_ready(dcache_io_maxi_w_ready),
    .io_maxi_w_valid(dcache_io_maxi_w_valid),
    .io_maxi_w_bits_data(dcache_io_maxi_w_bits_data),
    .io_maxi_w_bits_strb(dcache_io_maxi_w_bits_strb),
    .io_maxi_w_bits_last(dcache_io_maxi_w_bits_last),
    .io_maxi_b_valid(dcache_io_maxi_b_valid),
    .io_mmio_ar_ready(dcache_io_mmio_ar_ready),
    .io_mmio_ar_valid(dcache_io_mmio_ar_valid),
    .io_mmio_ar_bits_addr(dcache_io_mmio_ar_bits_addr),
    .io_mmio_ar_bits_size(dcache_io_mmio_ar_bits_size),
    .io_mmio_r_valid(dcache_io_mmio_r_valid),
    .io_mmio_r_bits_data(dcache_io_mmio_r_bits_data),
    .io_mmio_r_bits_last(dcache_io_mmio_r_bits_last),
    .io_mmio_aw_ready(dcache_io_mmio_aw_ready),
    .io_mmio_aw_valid(dcache_io_mmio_aw_valid),
    .io_mmio_aw_bits_addr(dcache_io_mmio_aw_bits_addr),
    .io_mmio_aw_bits_size(dcache_io_mmio_aw_bits_size),
    .io_mmio_w_ready(dcache_io_mmio_w_ready),
    .io_mmio_w_valid(dcache_io_mmio_w_valid),
    .io_mmio_w_bits_data(dcache_io_mmio_w_bits_data),
    .io_mmio_w_bits_strb(dcache_io_mmio_w_bits_strb),
    .io_mmio_w_bits_last(dcache_io_mmio_w_bits_last),
    .io_mmio_b_valid(dcache_io_mmio_b_valid),
    .io_sram4_addr(dcache_io_sram4_addr),
    .io_sram4_wen(dcache_io_sram4_wen),
    .io_sram4_wmask(dcache_io_sram4_wmask),
    .io_sram4_wdata(dcache_io_sram4_wdata),
    .io_sram4_rdata(dcache_io_sram4_rdata),
    .io_sram5_addr(dcache_io_sram5_addr),
    .io_sram5_wen(dcache_io_sram5_wen),
    .io_sram5_wmask(dcache_io_sram5_wmask),
    .io_sram5_wdata(dcache_io_sram5_wdata),
    .io_sram5_rdata(dcache_io_sram5_rdata),
    .io_sram6_addr(dcache_io_sram6_addr),
    .io_sram6_wen(dcache_io_sram6_wen),
    .io_sram6_wmask(dcache_io_sram6_wmask),
    .io_sram6_wdata(dcache_io_sram6_wdata),
    .io_sram6_rdata(dcache_io_sram6_rdata),
    .io_sram7_addr(dcache_io_sram7_addr),
    .io_sram7_wen(dcache_io_sram7_wen),
    .io_sram7_wmask(dcache_io_sram7_wmask),
    .io_sram7_wdata(dcache_io_sram7_wdata),
    .io_sram7_rdata(dcache_io_sram7_rdata),
    .clint_we(dcache_clint_we),
    ._T_24_0(dcache__T_24_0),
    .clint_rdata(dcache_clint_rdata),
    .clint_wdata(dcache_clint_wdata)
  );
  assign io_prev_ready = dcache_io_prev_ready; // @[MEMU.scala 65:14]
  assign io_next_valid = dcache_io_next_valid; // @[MEMU.scala 64:14]
  assign io_next_bits_id2wb_intr_exce_ret = dcache_io_next_bits_data_id2wb_intr_exce_ret; // @[MEMU.scala 53:13]
  assign io_next_bits_id2wb_fencei = dcache_io_next_bits_data_id2wb_fencei; // @[MEMU.scala 53:13]
  assign io_next_bits_id2wb_wb_sel = dcache_io_next_bits_data_id2wb_wb_sel; // @[MEMU.scala 53:13]
  assign io_next_bits_id2wb_regfile_we_en = dcache_io_next_bits_data_id2wb_regfile_we_en; // @[MEMU.scala 53:13]
  assign io_next_bits_id2wb_regfile_we_addr = dcache_io_next_bits_data_id2wb_regfile_we_addr; // @[MEMU.scala 53:13]
  assign io_next_bits_ex2wb_result_data = dcache_io_next_bits_data_ex2wb_result_data; // @[MEMU.scala 53:13]
  assign io_next_bits_mem2wb_memory_data = dcache_io_next_bits_data_mem2wb_memory_data; // @[MEMU.scala 53:13]
  assign io_maxi_ar_valid = dcache_io_maxi_ar_valid; // @[MEMU.scala 56:18]
  assign io_maxi_ar_bits_addr = dcache_io_maxi_ar_bits_addr; // @[MEMU.scala 56:18]
  assign io_maxi_ar_bits_len = dcache_io_maxi_ar_bits_len; // @[MEMU.scala 56:18]
  assign io_maxi_ar_bits_size = dcache_io_maxi_ar_bits_size; // @[MEMU.scala 56:18]
  assign io_maxi_aw_valid = dcache_io_maxi_aw_valid; // @[MEMU.scala 56:18]
  assign io_maxi_aw_bits_addr = dcache_io_maxi_aw_bits_addr; // @[MEMU.scala 56:18]
  assign io_maxi_aw_bits_len = dcache_io_maxi_aw_bits_len; // @[MEMU.scala 56:18]
  assign io_maxi_aw_bits_size = dcache_io_maxi_aw_bits_size; // @[MEMU.scala 56:18]
  assign io_maxi_w_valid = dcache_io_maxi_w_valid; // @[MEMU.scala 56:18]
  assign io_maxi_w_bits_data = dcache_io_maxi_w_bits_data; // @[MEMU.scala 56:18]
  assign io_maxi_w_bits_strb = dcache_io_maxi_w_bits_strb; // @[MEMU.scala 56:18]
  assign io_maxi_w_bits_last = dcache_io_maxi_w_bits_last; // @[MEMU.scala 56:18]
  assign io_mmio_ar_valid = dcache_io_mmio_ar_valid; // @[MEMU.scala 57:18]
  assign io_mmio_ar_bits_addr = dcache_io_mmio_ar_bits_addr; // @[MEMU.scala 57:18]
  assign io_mmio_ar_bits_size = dcache_io_mmio_ar_bits_size; // @[MEMU.scala 57:18]
  assign io_mmio_aw_valid = dcache_io_mmio_aw_valid; // @[MEMU.scala 57:18]
  assign io_mmio_aw_bits_addr = dcache_io_mmio_aw_bits_addr; // @[MEMU.scala 57:18]
  assign io_mmio_aw_bits_size = dcache_io_mmio_aw_bits_size; // @[MEMU.scala 57:18]
  assign io_mmio_w_valid = dcache_io_mmio_w_valid; // @[MEMU.scala 57:18]
  assign io_mmio_w_bits_data = dcache_io_mmio_w_bits_data; // @[MEMU.scala 57:18]
  assign io_mmio_w_bits_strb = dcache_io_mmio_w_bits_strb; // @[MEMU.scala 57:18]
  assign io_mmio_w_bits_last = dcache_io_mmio_w_bits_last; // @[MEMU.scala 57:18]
  assign io_sram4_addr = dcache_io_sram4_addr; // @[MEMU.scala 59:19]
  assign io_sram4_wen = dcache_io_sram4_wen; // @[MEMU.scala 59:19]
  assign io_sram4_wmask = dcache_io_sram4_wmask; // @[MEMU.scala 59:19]
  assign io_sram4_wdata = dcache_io_sram4_wdata; // @[MEMU.scala 59:19]
  assign io_sram5_addr = dcache_io_sram5_addr; // @[MEMU.scala 60:19]
  assign io_sram5_wen = dcache_io_sram5_wen; // @[MEMU.scala 60:19]
  assign io_sram5_wmask = dcache_io_sram5_wmask; // @[MEMU.scala 60:19]
  assign io_sram5_wdata = dcache_io_sram5_wdata; // @[MEMU.scala 60:19]
  assign io_sram6_addr = dcache_io_sram6_addr; // @[MEMU.scala 61:19]
  assign io_sram6_wen = dcache_io_sram6_wen; // @[MEMU.scala 61:19]
  assign io_sram6_wmask = dcache_io_sram6_wmask; // @[MEMU.scala 61:19]
  assign io_sram6_wdata = dcache_io_sram6_wdata; // @[MEMU.scala 61:19]
  assign io_sram7_addr = dcache_io_sram7_addr; // @[MEMU.scala 62:19]
  assign io_sram7_wen = dcache_io_sram7_wen; // @[MEMU.scala 62:19]
  assign io_sram7_wmask = dcache_io_sram7_wmask; // @[MEMU.scala 62:19]
  assign io_sram7_wdata = dcache_io_sram7_wdata; // @[MEMU.scala 62:19]
  assign clint_we = dcache_clint_we;
  assign _T_24 = dcache__T_24_0;
  assign clint_wdata = dcache_clint_wdata;
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_prev_valid = io_prev_valid; // @[MEMU.scala 46:24]
  assign dcache_io_prev_bits_data_id2mem_sext_flag = io_prev_bits_id2mem_sext_flag; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2mem_memory_rd_en = io_prev_bits_id2mem_memory_rd_en; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2mem_memory_we_en = io_prev_bits_id2mem_memory_we_en; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2wb_intr_exce_ret = io_prev_bits_id2wb_intr_exce_ret; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2wb_fencei = io_prev_bits_id2wb_fencei; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2wb_wb_sel = io_prev_bits_id2wb_wb_sel; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2wb_regfile_we_en = io_prev_bits_id2wb_regfile_we_en; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_id2wb_regfile_we_addr = io_prev_bits_id2wb_regfile_we_addr; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_ex2mem_we_data = io_prev_bits_ex2mem_we_data; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_data_ex2wb_result_data = io_prev_bits_ex2wb_result_data; // @[MEMU.scala 45:28]
  assign dcache_io_prev_bits_flush = io_prev_bits_id2mem_fencei; // @[MEMU.scala 51:29]
  assign dcache_io_prev_bits_wdata = io_prev_bits_ex2mem_we_data; // @[MEMU.scala 48:29]
  assign dcache_io_prev_bits_wmask = io_prev_bits_ex2mem_we_mask; // @[MEMU.scala 49:29]
  assign dcache_io_prev_bits_size_byte = io_prev_bits_id2mem_size_byte; // @[MEMU.scala 50:29]
  assign dcache_io_prev_bits_size_hword = io_prev_bits_id2mem_size_hword; // @[MEMU.scala 50:29]
  assign dcache_io_prev_bits_size_word = io_prev_bits_id2mem_size_word; // @[MEMU.scala 50:29]
  assign dcache_io_prev_bits_size_dword = io_prev_bits_id2mem_size_dword; // @[MEMU.scala 50:29]
  assign dcache_io_prev_bits_addr = io_prev_bits_ex2mem_addr; // @[MEMU.scala 47:29]
  assign dcache_io_maxi_ar_ready = io_maxi_ar_ready; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_r_valid = io_maxi_r_valid; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_r_bits_data = io_maxi_r_bits_data; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_r_bits_last = io_maxi_r_bits_last; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_aw_ready = io_maxi_aw_ready; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_w_ready = io_maxi_w_ready; // @[MEMU.scala 56:18]
  assign dcache_io_maxi_b_valid = io_maxi_b_valid; // @[MEMU.scala 56:18]
  assign dcache_io_mmio_ar_ready = io_mmio_ar_ready; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_r_valid = io_mmio_r_valid; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_r_bits_data = io_mmio_r_bits_data; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_r_bits_last = io_mmio_r_bits_last; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_aw_ready = io_mmio_aw_ready; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_w_ready = io_mmio_w_ready; // @[MEMU.scala 57:18]
  assign dcache_io_mmio_b_valid = io_mmio_b_valid; // @[MEMU.scala 57:18]
  assign dcache_io_sram4_rdata = io_sram4_rdata; // @[MEMU.scala 59:19]
  assign dcache_io_sram5_rdata = io_sram5_rdata; // @[MEMU.scala 60:19]
  assign dcache_io_sram6_rdata = io_sram6_rdata; // @[MEMU.scala 61:19]
  assign dcache_io_sram7_rdata = io_sram7_rdata; // @[MEMU.scala 62:19]
  assign dcache_clint_rdata = clint_rdata;
endmodule
module ysyx_040978_WBReg(
  input         clock,
  input         reset,
  input         io_prev_valid,
  input         io_prev_bits_id2wb_intr_exce_ret,
  input         io_prev_bits_id2wb_fencei,
  input         io_prev_bits_id2wb_wb_sel,
  input         io_prev_bits_id2wb_regfile_we_en,
  input  [4:0]  io_prev_bits_id2wb_regfile_we_addr,
  input  [63:0] io_prev_bits_ex2wb_result_data,
  input  [63:0] io_prev_bits_mem2wb_memory_data,
  output        io_next_valid,
  output        io_next_bits_id2wb_intr_exce_ret,
  output        io_next_bits_id2wb_fencei,
  output        io_next_bits_id2wb_wb_sel,
  output        io_next_bits_id2wb_regfile_we_en,
  output [4:0]  io_next_bits_id2wb_regfile_we_addr,
  output [63:0] io_next_bits_ex2wb_result_data,
  output [63:0] io_next_bits_mem2wb_memory_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  io_next_valid_r; // @[Reg.scala 27:20]
  wire  data_id2wb_intr_exce_ret = io_prev_valid & io_prev_bits_id2wb_intr_exce_ret; // @[WBU.scala 21:17]
  wire  data_id2wb_fencei = io_prev_valid & io_prev_bits_id2wb_fencei; // @[WBU.scala 21:17]
  wire  data_id2wb_wb_sel = io_prev_valid & io_prev_bits_id2wb_wb_sel; // @[WBU.scala 21:17]
  wire  data_id2wb_regfile_we_en = io_prev_valid & io_prev_bits_id2wb_regfile_we_en; // @[WBU.scala 21:17]
  reg  reg_id2wb_intr_exce_ret; // @[Reg.scala 27:20]
  reg  reg_id2wb_fencei; // @[Reg.scala 27:20]
  reg  reg_id2wb_wb_sel; // @[Reg.scala 27:20]
  reg  reg_id2wb_regfile_we_en; // @[Reg.scala 27:20]
  reg [4:0] reg_id2wb_regfile_we_addr; // @[Reg.scala 27:20]
  reg [63:0] reg_ex2wb_result_data; // @[Reg.scala 27:20]
  reg [63:0] reg_mem2wb_memory_data; // @[Reg.scala 27:20]
  assign io_next_valid = io_next_valid_r; // @[WBU.scala 19:11]
  assign io_next_bits_id2wb_intr_exce_ret = reg_id2wb_intr_exce_ret; // @[WBU.scala 23:12]
  assign io_next_bits_id2wb_fencei = reg_id2wb_fencei; // @[WBU.scala 23:12]
  assign io_next_bits_id2wb_wb_sel = reg_id2wb_wb_sel; // @[WBU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_en = reg_id2wb_regfile_we_en; // @[WBU.scala 23:12]
  assign io_next_bits_id2wb_regfile_we_addr = reg_id2wb_regfile_we_addr; // @[WBU.scala 23:12]
  assign io_next_bits_ex2wb_result_data = reg_ex2wb_result_data; // @[WBU.scala 23:12]
  assign io_next_bits_mem2wb_memory_data = reg_mem2wb_memory_data; // @[WBU.scala 23:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      io_next_valid_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      io_next_valid_r <= io_prev_valid;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_intr_exce_ret <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      reg_id2wb_intr_exce_ret <= data_id2wb_intr_exce_ret;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_fencei <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      reg_id2wb_fencei <= data_id2wb_fencei;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_wb_sel <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      reg_id2wb_wb_sel <= data_id2wb_wb_sel;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_en <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      reg_id2wb_regfile_we_en <= data_id2wb_regfile_we_en;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_id2wb_regfile_we_addr <= 5'h0; // @[Reg.scala 27:20]
    end else if (io_prev_valid) begin // @[WBU.scala 21:17]
      reg_id2wb_regfile_we_addr <= io_prev_bits_id2wb_regfile_we_addr;
    end else begin
      reg_id2wb_regfile_we_addr <= 5'h0;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_ex2wb_result_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_prev_valid) begin // @[WBU.scala 21:17]
      reg_ex2wb_result_data <= io_prev_bits_ex2wb_result_data;
    end else begin
      reg_ex2wb_result_data <= 64'h0;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg_mem2wb_memory_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_prev_valid) begin // @[WBU.scala 21:17]
      reg_mem2wb_memory_data <= io_prev_bits_mem2wb_memory_data;
    end else begin
      reg_mem2wb_memory_data <= 64'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_next_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_id2wb_intr_exce_ret = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_id2wb_fencei = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_id2wb_wb_sel = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reg_id2wb_regfile_we_en = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_id2wb_regfile_we_addr = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  reg_ex2wb_result_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_mem2wb_memory_data = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_WBU(
  input         io__prev_valid,
  input         io__prev_bits_id2wb_intr_exce_ret,
  input         io__prev_bits_id2wb_fencei,
  input         io__prev_bits_id2wb_wb_sel,
  input         io__prev_bits_id2wb_regfile_we_en,
  input  [4:0]  io__prev_bits_id2wb_regfile_we_addr,
  input  [63:0] io__prev_bits_ex2wb_result_data,
  input  [63:0] io__prev_bits_mem2wb_memory_data,
  output        io__regfile_en,
  output [4:0]  io__regfile_addr,
  output [63:0] io__regfile_data,
  output        io_prev_bits_id2wb_fencei,
  output        io_prev_bits_id2wb_intr_exce_ret
);
  assign io__regfile_en = io__prev_bits_id2wb_regfile_we_en & io__prev_valid; // @[WBU.scala 44:20]
  assign io__regfile_addr = io__prev_bits_id2wb_regfile_we_addr; // @[WBU.scala 45:11]
  assign io__regfile_data = io__prev_bits_id2wb_wb_sel ? io__prev_bits_mem2wb_memory_data :
    io__prev_bits_ex2wb_result_data; // @[WBU.scala 46:17]
  assign io_prev_bits_id2wb_fencei = io__prev_bits_id2wb_fencei;
  assign io_prev_bits_id2wb_intr_exce_ret = io__prev_bits_id2wb_intr_exce_ret;
endmodule
module ysyx_040978_FWU(
  output [63:0] io_idu_fw_src1_data,
  output [63:0] io_idu_fw_src2_data,
  output        io_idu_fw_ready,
  input         io_idu_optype_Itype,
  input  [4:0]  io_idu_src1_addr,
  input  [4:0]  io_idu_src2_addr,
  input  [63:0] io_idu_src1_data,
  input  [63:0] io_idu_src2_data,
  input         io_exu_is_load,
  input  [4:0]  io_exu_dst_addr,
  input  [63:0] io_exu_dst_data,
  input         io_memu_is_load_1,
  input  [4:0]  io_memu_dst_addr_1,
  input  [63:0] io_memu_dst_data_1,
  input  [4:0]  io_memu_dst_addr_2,
  input  [4:0]  io_wbu_dst_addr,
  input  [63:0] io_wbu_dst_data
);
  wire  ex_zero_n = io_exu_dst_addr != 5'h0; // @[FWU.scala 62:30]
  wire  mem1_zero_n = io_memu_dst_addr_1 != 5'h0; // @[FWU.scala 63:32]
  wire  mem2_zero_n = io_memu_dst_addr_2 != 5'h0; // @[FWU.scala 64:32]
  wire  wb_zero_n = io_wbu_dst_addr != 5'h0; // @[FWU.scala 65:30]
  wire  eq1_ex = io_idu_src1_addr == io_exu_dst_addr & ex_zero_n; // @[FWU.scala 68:43]
  wire  eq1_mem1 = io_idu_src1_addr == io_memu_dst_addr_1 & mem1_zero_n; // @[FWU.scala 69:43]
  wire  eq1_mem2 = io_idu_src1_addr == io_memu_dst_addr_2 & mem2_zero_n; // @[FWU.scala 70:43]
  wire  eq1_wb = io_idu_src1_addr == io_wbu_dst_addr & wb_zero_n; // @[FWU.scala 71:43]
  wire  eq2_ex = io_idu_src2_addr == io_exu_dst_addr & ex_zero_n; // @[FWU.scala 72:43]
  wire  eq2_mem1 = io_idu_src2_addr == io_memu_dst_addr_1 & mem1_zero_n; // @[FWU.scala 73:43]
  wire  eq2_mem2 = io_idu_src2_addr == io_memu_dst_addr_2 & mem2_zero_n; // @[FWU.scala 74:43]
  wire  eq2_wb = io_idu_src2_addr == io_wbu_dst_addr & wb_zero_n; // @[FWU.scala 75:43]
  wire  pre_is_load = (eq1_ex | eq2_ex) & io_exu_is_load | io_memu_is_load_1 | eq1_mem2 | eq2_mem2; // @[FWU.scala 77:82]
  wire [63:0] _io_idu_fw_src1_data_T = eq1_wb ? io_wbu_dst_data : io_idu_src1_data; // @[Mux.scala 98:16]
  wire [63:0] _io_idu_fw_src1_data_T_1 = eq1_mem1 ? io_memu_dst_data_1 : _io_idu_fw_src1_data_T; // @[Mux.scala 98:16]
  wire [63:0] _io_idu_fw_src2_data_T = eq2_wb ? io_wbu_dst_data : io_idu_src2_data; // @[Mux.scala 98:16]
  wire [63:0] _io_idu_fw_src2_data_T_1 = eq2_mem1 ? io_memu_dst_data_1 : _io_idu_fw_src2_data_T; // @[Mux.scala 98:16]
  wire [63:0] _io_idu_fw_src2_data_T_2 = eq2_ex ? io_exu_dst_data : _io_idu_fw_src2_data_T_1; // @[Mux.scala 98:16]
  assign io_idu_fw_src1_data = eq1_ex ? io_exu_dst_data : _io_idu_fw_src1_data_T_1; // @[Mux.scala 98:16]
  assign io_idu_fw_src2_data = io_idu_optype_Itype ? io_idu_src2_data : _io_idu_fw_src2_data_T_2; // @[Mux.scala 98:16]
  assign io_idu_fw_ready = ~pre_is_load; // @[FWU.scala 96:22]
endmodule
module ysyx_040978_BRU(
  input         clock,
  input         reset,
  input         io_idu_brh,
  input         io_idu_jal,
  input         io_idu_jalr,
  input  [63:0] io_idu_pc,
  input  [63:0] io_idu_src1,
  input  [63:0] io_idu_src2,
  input  [63:0] io_idu_imm,
  output        io_ifu_jump,
  output [63:0] io_ifu_npc,
  output        io_ifu_jump0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _jump_T = io_idu_brh | io_idu_jal; // @[BRU.scala 37:18]
  wire  jump = io_idu_brh | io_idu_jal | io_idu_jalr; // @[BRU.scala 37:24]
  reg  prev_jump; // @[BRU.scala 41:26]
  wire [63:0] _io_ifu_npc_T_2 = io_idu_pc + io_idu_imm; // @[BRU.scala 47:26]
  wire [63:0] _io_ifu_npc_T_4 = io_idu_src1 + io_idu_src2; // @[BRU.scala 48:32]
  wire [62:0] io_ifu_npc_hi = _io_ifu_npc_T_4[63:1]; // @[BRU.scala 48:39]
  wire [63:0] _io_ifu_npc_T_5 = {io_ifu_npc_hi,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _io_ifu_npc_T_7 = io_idu_jalr ? _io_ifu_npc_T_5 : 64'h0; // @[Mux.scala 98:16]
  assign io_ifu_jump = io_idu_brh | io_idu_jal | io_idu_jalr; // @[BRU.scala 37:24]
  assign io_ifu_npc = _jump_T ? _io_ifu_npc_T_2 : _io_ifu_npc_T_7; // @[Mux.scala 98:16]
  assign io_ifu_jump0 = ~prev_jump & jump; // @[BRU.scala 42:27]
  always @(posedge clock) begin
    if (reset) begin // @[BRU.scala 41:26]
      prev_jump <= 1'h0; // @[BRU.scala 41:26]
    end else begin
      prev_jump <= jump; // @[BRU.scala 41:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prev_jump = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_RegFile(
  input         clock,
  input         reset,
  input         io_wbu_en,
  input  [4:0]  io_wbu_addr,
  input  [63:0] io_wbu_data,
  input  [4:0]  io_idu_addr1,
  output [63:0] io_idu_data1,
  input  [4:0]  io_idu_addr2,
  output [63:0] io_idu_data2
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] gpr_1; // @[RegFile.scala 22:20]
  reg [63:0] gpr_2; // @[RegFile.scala 22:20]
  reg [63:0] gpr_3; // @[RegFile.scala 22:20]
  reg [63:0] gpr_4; // @[RegFile.scala 22:20]
  reg [63:0] gpr_5; // @[RegFile.scala 22:20]
  reg [63:0] gpr_6; // @[RegFile.scala 22:20]
  reg [63:0] gpr_7; // @[RegFile.scala 22:20]
  reg [63:0] gpr_8; // @[RegFile.scala 22:20]
  reg [63:0] gpr_9; // @[RegFile.scala 22:20]
  reg [63:0] gpr_10; // @[RegFile.scala 22:20]
  reg [63:0] gpr_11; // @[RegFile.scala 22:20]
  reg [63:0] gpr_12; // @[RegFile.scala 22:20]
  reg [63:0] gpr_13; // @[RegFile.scala 22:20]
  reg [63:0] gpr_14; // @[RegFile.scala 22:20]
  reg [63:0] gpr_15; // @[RegFile.scala 22:20]
  reg [63:0] gpr_16; // @[RegFile.scala 22:20]
  reg [63:0] gpr_17; // @[RegFile.scala 22:20]
  reg [63:0] gpr_18; // @[RegFile.scala 22:20]
  reg [63:0] gpr_19; // @[RegFile.scala 22:20]
  reg [63:0] gpr_20; // @[RegFile.scala 22:20]
  reg [63:0] gpr_21; // @[RegFile.scala 22:20]
  reg [63:0] gpr_22; // @[RegFile.scala 22:20]
  reg [63:0] gpr_23; // @[RegFile.scala 22:20]
  reg [63:0] gpr_24; // @[RegFile.scala 22:20]
  reg [63:0] gpr_25; // @[RegFile.scala 22:20]
  reg [63:0] gpr_26; // @[RegFile.scala 22:20]
  reg [63:0] gpr_27; // @[RegFile.scala 22:20]
  reg [63:0] gpr_28; // @[RegFile.scala 22:20]
  reg [63:0] gpr_29; // @[RegFile.scala 22:20]
  reg [63:0] gpr_30; // @[RegFile.scala 22:20]
  reg [63:0] gpr_31; // @[RegFile.scala 22:20]
  wire [63:0] _GEN_1 = 5'h1 == io_idu_addr1 ? gpr_1 : 64'h0; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_2 = 5'h2 == io_idu_addr1 ? gpr_2 : _GEN_1; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_3 = 5'h3 == io_idu_addr1 ? gpr_3 : _GEN_2; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_4 = 5'h4 == io_idu_addr1 ? gpr_4 : _GEN_3; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_5 = 5'h5 == io_idu_addr1 ? gpr_5 : _GEN_4; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_6 = 5'h6 == io_idu_addr1 ? gpr_6 : _GEN_5; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_7 = 5'h7 == io_idu_addr1 ? gpr_7 : _GEN_6; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_8 = 5'h8 == io_idu_addr1 ? gpr_8 : _GEN_7; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_9 = 5'h9 == io_idu_addr1 ? gpr_9 : _GEN_8; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_10 = 5'ha == io_idu_addr1 ? gpr_10 : _GEN_9; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_11 = 5'hb == io_idu_addr1 ? gpr_11 : _GEN_10; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_12 = 5'hc == io_idu_addr1 ? gpr_12 : _GEN_11; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_13 = 5'hd == io_idu_addr1 ? gpr_13 : _GEN_12; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_14 = 5'he == io_idu_addr1 ? gpr_14 : _GEN_13; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_15 = 5'hf == io_idu_addr1 ? gpr_15 : _GEN_14; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_16 = 5'h10 == io_idu_addr1 ? gpr_16 : _GEN_15; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_17 = 5'h11 == io_idu_addr1 ? gpr_17 : _GEN_16; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_18 = 5'h12 == io_idu_addr1 ? gpr_18 : _GEN_17; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_19 = 5'h13 == io_idu_addr1 ? gpr_19 : _GEN_18; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_20 = 5'h14 == io_idu_addr1 ? gpr_20 : _GEN_19; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_21 = 5'h15 == io_idu_addr1 ? gpr_21 : _GEN_20; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_22 = 5'h16 == io_idu_addr1 ? gpr_22 : _GEN_21; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_23 = 5'h17 == io_idu_addr1 ? gpr_23 : _GEN_22; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_24 = 5'h18 == io_idu_addr1 ? gpr_24 : _GEN_23; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_25 = 5'h19 == io_idu_addr1 ? gpr_25 : _GEN_24; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_26 = 5'h1a == io_idu_addr1 ? gpr_26 : _GEN_25; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_27 = 5'h1b == io_idu_addr1 ? gpr_27 : _GEN_26; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_28 = 5'h1c == io_idu_addr1 ? gpr_28 : _GEN_27; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_29 = 5'h1d == io_idu_addr1 ? gpr_29 : _GEN_28; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_30 = 5'h1e == io_idu_addr1 ? gpr_30 : _GEN_29; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  wire [63:0] _GEN_33 = 5'h1 == io_idu_addr2 ? gpr_1 : 64'h0; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_34 = 5'h2 == io_idu_addr2 ? gpr_2 : _GEN_33; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_35 = 5'h3 == io_idu_addr2 ? gpr_3 : _GEN_34; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_36 = 5'h4 == io_idu_addr2 ? gpr_4 : _GEN_35; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_37 = 5'h5 == io_idu_addr2 ? gpr_5 : _GEN_36; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_38 = 5'h6 == io_idu_addr2 ? gpr_6 : _GEN_37; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_39 = 5'h7 == io_idu_addr2 ? gpr_7 : _GEN_38; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_40 = 5'h8 == io_idu_addr2 ? gpr_8 : _GEN_39; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_41 = 5'h9 == io_idu_addr2 ? gpr_9 : _GEN_40; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_42 = 5'ha == io_idu_addr2 ? gpr_10 : _GEN_41; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_43 = 5'hb == io_idu_addr2 ? gpr_11 : _GEN_42; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_44 = 5'hc == io_idu_addr2 ? gpr_12 : _GEN_43; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_45 = 5'hd == io_idu_addr2 ? gpr_13 : _GEN_44; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_46 = 5'he == io_idu_addr2 ? gpr_14 : _GEN_45; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_47 = 5'hf == io_idu_addr2 ? gpr_15 : _GEN_46; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_48 = 5'h10 == io_idu_addr2 ? gpr_16 : _GEN_47; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_49 = 5'h11 == io_idu_addr2 ? gpr_17 : _GEN_48; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_50 = 5'h12 == io_idu_addr2 ? gpr_18 : _GEN_49; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_51 = 5'h13 == io_idu_addr2 ? gpr_19 : _GEN_50; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_52 = 5'h14 == io_idu_addr2 ? gpr_20 : _GEN_51; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_53 = 5'h15 == io_idu_addr2 ? gpr_21 : _GEN_52; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_54 = 5'h16 == io_idu_addr2 ? gpr_22 : _GEN_53; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_55 = 5'h17 == io_idu_addr2 ? gpr_23 : _GEN_54; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_56 = 5'h18 == io_idu_addr2 ? gpr_24 : _GEN_55; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_57 = 5'h19 == io_idu_addr2 ? gpr_25 : _GEN_56; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_58 = 5'h1a == io_idu_addr2 ? gpr_26 : _GEN_57; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_59 = 5'h1b == io_idu_addr2 ? gpr_27 : _GEN_58; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_60 = 5'h1c == io_idu_addr2 ? gpr_28 : _GEN_59; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_61 = 5'h1d == io_idu_addr2 ? gpr_29 : _GEN_60; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_62 = 5'h1e == io_idu_addr2 ? gpr_30 : _GEN_61; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  wire [63:0] _GEN_65 = 5'h1 == io_wbu_addr ? gpr_1 : 64'h0; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_66 = 5'h2 == io_wbu_addr ? gpr_2 : _GEN_65; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_67 = 5'h3 == io_wbu_addr ? gpr_3 : _GEN_66; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_68 = 5'h4 == io_wbu_addr ? gpr_4 : _GEN_67; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_69 = 5'h5 == io_wbu_addr ? gpr_5 : _GEN_68; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_70 = 5'h6 == io_wbu_addr ? gpr_6 : _GEN_69; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_71 = 5'h7 == io_wbu_addr ? gpr_7 : _GEN_70; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_72 = 5'h8 == io_wbu_addr ? gpr_8 : _GEN_71; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_73 = 5'h9 == io_wbu_addr ? gpr_9 : _GEN_72; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_74 = 5'ha == io_wbu_addr ? gpr_10 : _GEN_73; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_75 = 5'hb == io_wbu_addr ? gpr_11 : _GEN_74; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_76 = 5'hc == io_wbu_addr ? gpr_12 : _GEN_75; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_77 = 5'hd == io_wbu_addr ? gpr_13 : _GEN_76; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_78 = 5'he == io_wbu_addr ? gpr_14 : _GEN_77; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_79 = 5'hf == io_wbu_addr ? gpr_15 : _GEN_78; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_80 = 5'h10 == io_wbu_addr ? gpr_16 : _GEN_79; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_81 = 5'h11 == io_wbu_addr ? gpr_17 : _GEN_80; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_82 = 5'h12 == io_wbu_addr ? gpr_18 : _GEN_81; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_83 = 5'h13 == io_wbu_addr ? gpr_19 : _GEN_82; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_84 = 5'h14 == io_wbu_addr ? gpr_20 : _GEN_83; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_85 = 5'h15 == io_wbu_addr ? gpr_21 : _GEN_84; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_86 = 5'h16 == io_wbu_addr ? gpr_22 : _GEN_85; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_87 = 5'h17 == io_wbu_addr ? gpr_23 : _GEN_86; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_88 = 5'h18 == io_wbu_addr ? gpr_24 : _GEN_87; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_89 = 5'h19 == io_wbu_addr ? gpr_25 : _GEN_88; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_90 = 5'h1a == io_wbu_addr ? gpr_26 : _GEN_89; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_91 = 5'h1b == io_wbu_addr ? gpr_27 : _GEN_90; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_92 = 5'h1c == io_wbu_addr ? gpr_28 : _GEN_91; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_93 = 5'h1d == io_wbu_addr ? gpr_29 : _GEN_92; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  wire [63:0] _GEN_94 = 5'h1e == io_wbu_addr ? gpr_30 : _GEN_93; // @[RegFile.scala 26:26 RegFile.scala 26:26]
  assign io_idu_data1 = 5'h1f == io_idu_addr1 ? gpr_31 : _GEN_30; // @[RegFile.scala 23:16 RegFile.scala 23:16]
  assign io_idu_data2 = 5'h1f == io_idu_addr2 ? gpr_31 : _GEN_62; // @[RegFile.scala 24:16 RegFile.scala 24:16]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_1 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_1 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_1 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_1 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_2 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h2 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_2 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_2 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_2 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_3 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h3 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_3 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_3 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_3 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_4 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h4 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_4 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_4 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_4 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_5 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h5 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_5 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_5 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_5 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_6 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h6 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_6 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_6 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_6 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_7 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h7 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_7 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_7 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_7 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_8 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h8 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_8 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_8 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_8 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_9 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h9 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_9 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_9 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_9 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_10 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'ha == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_10 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_10 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_10 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_11 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'hb == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_11 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_11 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_11 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_12 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'hc == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_12 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_12 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_12 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_13 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'hd == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_13 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_13 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_13 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_14 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'he == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_14 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_14 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_14 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_15 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'hf == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_15 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_15 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_15 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_16 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h10 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_16 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_16 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_16 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_17 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h11 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_17 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_17 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_17 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_18 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h12 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_18 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_18 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_18 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_19 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h13 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_19 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_19 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_19 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_20 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h14 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_20 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_20 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_20 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_21 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h15 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_21 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_21 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_21 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_22 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h16 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_22 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_22 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_22 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_23 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h17 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_23 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_23 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_23 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_24 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h18 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_24 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_24 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_24 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_25 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h19 == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_25 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_25 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_25 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_26 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1a == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_26 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_26 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_26 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_27 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1b == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_27 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_27 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_27 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_28 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1c == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_28 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_28 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_28 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_29 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1d == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_29 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_29 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_29 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_30 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1e == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_30 <= io_wbu_data;
      end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:26]
        gpr_30 <= gpr_31; // @[RegFile.scala 26:26]
      end else begin
        gpr_30 <= _GEN_94;
      end
    end
    if (reset) begin // @[RegFile.scala 22:20]
      gpr_31 <= 64'h0; // @[RegFile.scala 22:20]
    end else if (5'h1f == io_wbu_addr) begin // @[RegFile.scala 26:20]
      if (io_wbu_en) begin // @[RegFile.scala 26:26]
        gpr_31 <= io_wbu_data;
      end else if (!(5'h1f == io_wbu_addr)) begin // @[RegFile.scala 26:26]
        gpr_31 <= _GEN_94;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  gpr_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  gpr_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  gpr_3 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  gpr_4 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  gpr_5 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  gpr_6 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  gpr_7 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  gpr_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  gpr_9 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  gpr_10 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  gpr_11 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  gpr_12 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  gpr_13 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  gpr_14 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  gpr_15 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  gpr_16 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  gpr_17 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  gpr_18 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  gpr_19 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  gpr_20 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  gpr_21 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  gpr_22 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  gpr_23 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  gpr_24 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  gpr_25 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  gpr_26 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  gpr_27 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  gpr_28 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  gpr_29 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  gpr_30 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  gpr_31 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_SparkCore(
  input          clock,
  input          reset,
  input          io_maxi4_ar_ready,
  output         io_maxi4_ar_valid,
  output [31:0]  io_maxi4_ar_bits_addr,
  output [1:0]   io_maxi4_ar_bits_burst,
  output [3:0]   io_maxi4_ar_bits_id,
  output [7:0]   io_maxi4_ar_bits_len,
  output [2:0]   io_maxi4_ar_bits_size,
  output         io_maxi4_r_ready,
  input          io_maxi4_r_valid,
  input  [63:0]  io_maxi4_r_bits_data,
  input  [3:0]   io_maxi4_r_bits_id,
  input          io_maxi4_r_bits_last,
  input  [1:0]   io_maxi4_r_bits_resp,
  input          io_maxi4_aw_ready,
  output         io_maxi4_aw_valid,
  output [31:0]  io_maxi4_aw_bits_addr,
  output [1:0]   io_maxi4_aw_bits_burst,
  output [3:0]   io_maxi4_aw_bits_id,
  output [7:0]   io_maxi4_aw_bits_len,
  output [2:0]   io_maxi4_aw_bits_size,
  input          io_maxi4_w_ready,
  output         io_maxi4_w_valid,
  output [63:0]  io_maxi4_w_bits_data,
  output [7:0]   io_maxi4_w_bits_strb,
  output         io_maxi4_w_bits_last,
  output         io_maxi4_b_ready,
  input          io_maxi4_b_valid,
  input  [3:0]   io_maxi4_b_bits_id,
  input  [1:0]   io_maxi4_b_bits_resp,
  input          io_sideband_clint_msip,
  input          io_sideband_clint_mtip,
  input  [63:0]  io_sideband_clint_mtime,
  input          io_sideband_meip,
  output [5:0]   io_sram0_addr,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,
  output         clint_we,
  output [31:0]  _T_24,
  input  [63:0]  clint_rdata,
  output [63:0]  clint_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  icon_clock; // @[AXI.scala 285:30]
  wire  icon_reset; // @[AXI.scala 285:30]
  wire  icon_io_maxi_ar_ready; // @[AXI.scala 285:30]
  wire  icon_io_maxi_ar_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_maxi_ar_bits_addr; // @[AXI.scala 285:30]
  wire [3:0] icon_io_maxi_ar_bits_id; // @[AXI.scala 285:30]
  wire [7:0] icon_io_maxi_ar_bits_len; // @[AXI.scala 285:30]
  wire [2:0] icon_io_maxi_ar_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_maxi_r_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_maxi_r_bits_data; // @[AXI.scala 285:30]
  wire [3:0] icon_io_maxi_r_bits_id; // @[AXI.scala 285:30]
  wire  icon_io_maxi_r_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_maxi_aw_ready; // @[AXI.scala 285:30]
  wire  icon_io_maxi_aw_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_maxi_aw_bits_addr; // @[AXI.scala 285:30]
  wire [3:0] icon_io_maxi_aw_bits_id; // @[AXI.scala 285:30]
  wire [7:0] icon_io_maxi_aw_bits_len; // @[AXI.scala 285:30]
  wire [2:0] icon_io_maxi_aw_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_maxi_w_ready; // @[AXI.scala 285:30]
  wire  icon_io_maxi_w_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_maxi_w_bits_data; // @[AXI.scala 285:30]
  wire [7:0] icon_io_maxi_w_bits_strb; // @[AXI.scala 285:30]
  wire  icon_io_maxi_w_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_maxi_b_valid; // @[AXI.scala 285:30]
  wire [3:0] icon_io_maxi_b_bits_id; // @[AXI.scala 285:30]
  wire  icon_io_ifu_ar_ready; // @[AXI.scala 285:30]
  wire  icon_io_ifu_ar_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_ifu_ar_bits_addr; // @[AXI.scala 285:30]
  wire [7:0] icon_io_ifu_ar_bits_len; // @[AXI.scala 285:30]
  wire [2:0] icon_io_ifu_ar_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_ifu_r_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_ifu_r_bits_data; // @[AXI.scala 285:30]
  wire  icon_io_ifu_r_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_memu_ar_ready; // @[AXI.scala 285:30]
  wire  icon_io_memu_ar_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_memu_ar_bits_addr; // @[AXI.scala 285:30]
  wire [7:0] icon_io_memu_ar_bits_len; // @[AXI.scala 285:30]
  wire [2:0] icon_io_memu_ar_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_memu_r_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_memu_r_bits_data; // @[AXI.scala 285:30]
  wire  icon_io_memu_r_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_memu_aw_ready; // @[AXI.scala 285:30]
  wire  icon_io_memu_aw_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_memu_aw_bits_addr; // @[AXI.scala 285:30]
  wire [7:0] icon_io_memu_aw_bits_len; // @[AXI.scala 285:30]
  wire [2:0] icon_io_memu_aw_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_memu_w_ready; // @[AXI.scala 285:30]
  wire  icon_io_memu_w_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_memu_w_bits_data; // @[AXI.scala 285:30]
  wire [7:0] icon_io_memu_w_bits_strb; // @[AXI.scala 285:30]
  wire  icon_io_memu_w_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_memu_b_valid; // @[AXI.scala 285:30]
  wire  icon_io_devu_ar_ready; // @[AXI.scala 285:30]
  wire  icon_io_devu_ar_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_devu_ar_bits_addr; // @[AXI.scala 285:30]
  wire [2:0] icon_io_devu_ar_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_devu_r_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_devu_r_bits_data; // @[AXI.scala 285:30]
  wire  icon_io_devu_r_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_devu_aw_ready; // @[AXI.scala 285:30]
  wire  icon_io_devu_aw_valid; // @[AXI.scala 285:30]
  wire [31:0] icon_io_devu_aw_bits_addr; // @[AXI.scala 285:30]
  wire [2:0] icon_io_devu_aw_bits_size; // @[AXI.scala 285:30]
  wire  icon_io_devu_w_ready; // @[AXI.scala 285:30]
  wire  icon_io_devu_w_valid; // @[AXI.scala 285:30]
  wire [63:0] icon_io_devu_w_bits_data; // @[AXI.scala 285:30]
  wire [7:0] icon_io_devu_w_bits_strb; // @[AXI.scala 285:30]
  wire  icon_io_devu_w_bits_last; // @[AXI.scala 285:30]
  wire  icon_io_devu_b_valid; // @[AXI.scala 285:30]
  wire  pc_clock; // @[IFU.scala 96:20]
  wire  pc_reset; // @[IFU.scala 96:20]
  wire  pc_io_jump0; // @[IFU.scala 96:20]
  wire  pc_io_jump; // @[IFU.scala 96:20]
  wire [63:0] pc_io_npc; // @[IFU.scala 96:20]
  wire  pc_io_sys_ready; // @[IFU.scala 96:20]
  wire  pc_io_next_ready; // @[IFU.scala 96:20]
  wire  pc_io_next_valid; // @[IFU.scala 96:20]
  wire [63:0] pc_io_next_bits_pc2if_pc; // @[IFU.scala 96:20]
  wire  ifu_clock; // @[IFU.scala 102:21]
  wire  ifu_reset; // @[IFU.scala 102:21]
  wire  ifu_io_cache_reset; // @[IFU.scala 102:21]
  wire  ifu_io_prev_ready; // @[IFU.scala 102:21]
  wire  ifu_io_prev_valid; // @[IFU.scala 102:21]
  wire [63:0] ifu_io_prev_bits_pc2if_pc; // @[IFU.scala 102:21]
  wire  ifu_io_maxi_ar_ready; // @[IFU.scala 102:21]
  wire  ifu_io_maxi_ar_valid; // @[IFU.scala 102:21]
  wire [31:0] ifu_io_maxi_ar_bits_addr; // @[IFU.scala 102:21]
  wire [7:0] ifu_io_maxi_ar_bits_len; // @[IFU.scala 102:21]
  wire [2:0] ifu_io_maxi_ar_bits_size; // @[IFU.scala 102:21]
  wire  ifu_io_maxi_r_valid; // @[IFU.scala 102:21]
  wire [63:0] ifu_io_maxi_r_bits_data; // @[IFU.scala 102:21]
  wire  ifu_io_maxi_r_bits_last; // @[IFU.scala 102:21]
  wire  ifu_io_next_ready; // @[IFU.scala 102:21]
  wire  ifu_io_next_valid; // @[IFU.scala 102:21]
  wire [31:0] ifu_io_next_bits_if2id_inst; // @[IFU.scala 102:21]
  wire [63:0] ifu_io_next_bits_if2id_pc; // @[IFU.scala 102:21]
  wire [5:0] ifu_io_sram0_addr; // @[IFU.scala 102:21]
  wire  ifu_io_sram0_wen; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram0_wmask; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram0_wdata; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram0_rdata; // @[IFU.scala 102:21]
  wire [5:0] ifu_io_sram1_addr; // @[IFU.scala 102:21]
  wire  ifu_io_sram1_wen; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram1_wmask; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram1_wdata; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram1_rdata; // @[IFU.scala 102:21]
  wire [5:0] ifu_io_sram2_addr; // @[IFU.scala 102:21]
  wire  ifu_io_sram2_wen; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram2_wmask; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram2_wdata; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram2_rdata; // @[IFU.scala 102:21]
  wire [5:0] ifu_io_sram3_addr; // @[IFU.scala 102:21]
  wire  ifu_io_sram3_wen; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram3_wmask; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram3_wdata; // @[IFU.scala 102:21]
  wire [127:0] ifu_io_sram3_rdata; // @[IFU.scala 102:21]
  wire  ifu_fenceiing; // @[IFU.scala 102:21]
  wire  IF2IDReg_clock; // @[IDU.scala 286:26]
  wire  IF2IDReg_reset; // @[IDU.scala 286:26]
  wire  IF2IDReg_io_prev_ready; // @[IDU.scala 286:26]
  wire  IF2IDReg_io_prev_valid; // @[IDU.scala 286:26]
  wire [31:0] IF2IDReg_io_prev_bits_if2id_inst; // @[IDU.scala 286:26]
  wire [63:0] IF2IDReg_io_prev_bits_if2id_pc; // @[IDU.scala 286:26]
  wire  IF2IDReg_io_next_ready; // @[IDU.scala 286:26]
  wire  IF2IDReg_io_next_valid; // @[IDU.scala 286:26]
  wire [31:0] IF2IDReg_io_next_bits_if2id_inst; // @[IDU.scala 286:26]
  wire [63:0] IF2IDReg_io_next_bits_if2id_pc; // @[IDU.scala 286:26]
  wire  idu_clock; // @[IDU.scala 290:21]
  wire  idu_reset; // @[IDU.scala 290:21]
  wire [4:0] idu_io_regfile_addr1; // @[IDU.scala 290:21]
  wire [63:0] idu_io_regfile_data1; // @[IDU.scala 290:21]
  wire [4:0] idu_io_regfile_addr2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_regfile_data2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_fwu_fw_src1_data; // @[IDU.scala 290:21]
  wire [63:0] idu_io_fwu_fw_src2_data; // @[IDU.scala 290:21]
  wire  idu_io_fwu_optype_Itype; // @[IDU.scala 290:21]
  wire [4:0] idu_io_fwu_src1_addr; // @[IDU.scala 290:21]
  wire [4:0] idu_io_fwu_src2_addr; // @[IDU.scala 290:21]
  wire [63:0] idu_io_fwu_src1_data; // @[IDU.scala 290:21]
  wire [63:0] idu_io_fwu_src2_data; // @[IDU.scala 290:21]
  wire  idu_io_bru_brh; // @[IDU.scala 290:21]
  wire  idu_io_bru_jal; // @[IDU.scala 290:21]
  wire  idu_io_bru_jalr; // @[IDU.scala 290:21]
  wire [63:0] idu_io_bru_pc; // @[IDU.scala 290:21]
  wire [63:0] idu_io_bru_src1; // @[IDU.scala 290:21]
  wire [63:0] idu_io_bru_src2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_bru_imm; // @[IDU.scala 290:21]
  wire [63:0] idu_io_csr_out_mepc; // @[IDU.scala 290:21]
  wire [63:0] idu_io_csr_out_mtvec; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_mie; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_mtie; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_msie; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_meie; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_mtip; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_msip; // @[IDU.scala 290:21]
  wire  idu_io_csr_out_meip; // @[IDU.scala 290:21]
  wire  idu_io_prev_ready; // @[IDU.scala 290:21]
  wire  idu_io_prev_valid; // @[IDU.scala 290:21]
  wire [31:0] idu_io_prev_bits_if2id_inst; // @[IDU.scala 290:21]
  wire [63:0] idu_io_prev_bits_if2id_pc; // @[IDU.scala 290:21]
  wire  idu_io_next_ready; // @[IDU.scala 290:21]
  wire  idu_io_next_valid; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_alu_src1; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_alu_src2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_salu_src1; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_salu_src2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_src1; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_src2; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_src3; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_auipc; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_lui; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_jal; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_jalr; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sb; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sh; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sw; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sd; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_add; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sub; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sll; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_slt; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sltu; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_xor; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_srl; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_sra; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_or; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_and; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_is_csr; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrw; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrs; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrc; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrwi; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrsi; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_operator_csr_csrrci; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_srcsize_byte; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_srcsize_hword; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_srcsize_word; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_srcsize_dword; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_is_load; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_is_save; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_div_inf; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_we; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mepc; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mtvec; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mstatus; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mie; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mcause; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mip; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mtime; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mcycle; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_csr_hit_is_mhartid; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mdu_op_mul_signed; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mdu_op_is_mu; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mdu_op_mul_32; // @[IDU.scala 290:21]
  wire [1:0] idu_io_next_bits_id2ex_mdu_op_div_signed; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mdu_op_is_div; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mdu_op_is_du; // @[IDU.scala 290:21]
  wire [4:0] idu_io_next_bits_id2ex_zimm; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_intr; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_exec; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_mret; // @[IDU.scala 290:21]
  wire [3:0] idu_io_next_bits_id2ex_exce_code; // @[IDU.scala 290:21]
  wire [63:0] idu_io_next_bits_id2ex_pc; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2ex_is_iem; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_fencei; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_size_byte; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_size_hword; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_size_word; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_size_dword; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_sext_flag; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_memory_rd_en; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2mem_memory_we_en; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2wb_intr_exce_ret; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2wb_fencei; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2wb_wb_sel; // @[IDU.scala 290:21]
  wire  idu_io_next_bits_id2wb_regfile_we_en; // @[IDU.scala 290:21]
  wire [4:0] idu_io_next_bits_id2wb_regfile_we_addr; // @[IDU.scala 290:21]
  wire  idu_wb_fencei_0; // @[IDU.scala 290:21]
  wire  idu_wb_intr_exce_ret_0; // @[IDU.scala 290:21]
  wire  idu_fenceiing_0; // @[IDU.scala 290:21]
  wire  ID2EXReg_clock; // @[EXU.scala 155:26]
  wire  ID2EXReg_reset; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_ready; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_valid; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_alu_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_alu_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_salu_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_salu_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_src3; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_auipc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_lui; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_jal; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_jalr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sb; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sh; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sw; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sd; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_add; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sub; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sll; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_slt; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sltu; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_xor; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_srl; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_sra; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_or; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_and; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_is_csr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_srcsize_byte; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_srcsize_hword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_srcsize_word; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_srcsize_dword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_is_load; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_is_save; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_div_inf; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_we; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 155:26]
  wire [1:0] ID2EXReg_io_prev_bits_id2ex_mdu_op_div_signed; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mdu_op_is_div; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mdu_op_is_du; // @[EXU.scala 155:26]
  wire [4:0] ID2EXReg_io_prev_bits_id2ex_zimm; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_intr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_exec; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_mret; // @[EXU.scala 155:26]
  wire [3:0] ID2EXReg_io_prev_bits_id2ex_exce_code; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_prev_bits_id2ex_pc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2ex_is_iem; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_fencei; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_size_byte; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_size_hword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_size_word; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_size_dword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_sext_flag; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_memory_rd_en; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2mem_memory_we_en; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2wb_intr_exce_ret; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2wb_fencei; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2wb_wb_sel; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_prev_bits_id2wb_regfile_we_en; // @[EXU.scala 155:26]
  wire [4:0] ID2EXReg_io_prev_bits_id2wb_regfile_we_addr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_ready; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_valid; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_alu_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_alu_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_salu_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_salu_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_src1; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_src2; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_src3; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_auipc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_lui; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_jal; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_jalr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sb; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sh; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sw; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sd; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_add; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sub; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sll; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_slt; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sltu; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_xor; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_srl; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_sra; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_or; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_and; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_is_csr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_srcsize_byte; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_srcsize_hword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_srcsize_word; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_srcsize_dword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_is_load; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_is_save; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_div_inf; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_we; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 155:26]
  wire [1:0] ID2EXReg_io_next_bits_id2ex_mdu_op_div_signed; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mdu_op_is_div; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mdu_op_is_du; // @[EXU.scala 155:26]
  wire [4:0] ID2EXReg_io_next_bits_id2ex_zimm; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_intr; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_exec; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_mret; // @[EXU.scala 155:26]
  wire [3:0] ID2EXReg_io_next_bits_id2ex_exce_code; // @[EXU.scala 155:26]
  wire [63:0] ID2EXReg_io_next_bits_id2ex_pc; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2ex_is_iem; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_fencei; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_size_byte; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_size_hword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_size_word; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_size_dword; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_sext_flag; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_memory_rd_en; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2mem_memory_we_en; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2wb_intr_exce_ret; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2wb_fencei; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2wb_wb_sel; // @[EXU.scala 155:26]
  wire  ID2EXReg_io_next_bits_id2wb_regfile_we_en; // @[EXU.scala 155:26]
  wire [4:0] ID2EXReg_io_next_bits_id2wb_regfile_we_addr; // @[EXU.scala 155:26]
  wire  exu_clock; // @[EXU.scala 158:21]
  wire  exu_reset; // @[EXU.scala 158:21]
  wire  exu_io_prev_ready; // @[EXU.scala 158:21]
  wire  exu_io_prev_valid; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_alu_src1; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_alu_src2; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_salu_src1; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_salu_src2; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_src1; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_src2; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_src3; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_auipc; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_lui; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_jal; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_jalr; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sb; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sh; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sw; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sd; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_add; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sub; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sll; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_slt; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sltu; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_xor; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_srl; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_sra; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_or; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_and; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_is_csr; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_srcsize_byte; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_srcsize_hword; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_srcsize_word; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_srcsize_dword; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_is_load; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_is_save; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_div_inf; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_we; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 158:21]
  wire [1:0] exu_io_prev_bits_id2ex_mdu_op_div_signed; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mdu_op_is_div; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mdu_op_is_du; // @[EXU.scala 158:21]
  wire [4:0] exu_io_prev_bits_id2ex_zimm; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_intr; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_exec; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_mret; // @[EXU.scala 158:21]
  wire [3:0] exu_io_prev_bits_id2ex_exce_code; // @[EXU.scala 158:21]
  wire [63:0] exu_io_prev_bits_id2ex_pc; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2ex_is_iem; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_fencei; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_size_byte; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_size_hword; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_size_word; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_size_dword; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_sext_flag; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_memory_rd_en; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2mem_memory_we_en; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2wb_intr_exce_ret; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2wb_fencei; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2wb_wb_sel; // @[EXU.scala 158:21]
  wire  exu_io_prev_bits_id2wb_regfile_we_en; // @[EXU.scala 158:21]
  wire [4:0] exu_io_prev_bits_id2wb_regfile_we_addr; // @[EXU.scala 158:21]
  wire  exu_io_next_ready; // @[EXU.scala 158:21]
  wire  exu_io_next_valid; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_fencei; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_size_byte; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_size_hword; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_size_word; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_size_dword; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_sext_flag; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_memory_rd_en; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2mem_memory_we_en; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2wb_intr_exce_ret; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2wb_fencei; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2wb_wb_sel; // @[EXU.scala 158:21]
  wire  exu_io_next_bits_id2wb_regfile_we_en; // @[EXU.scala 158:21]
  wire [4:0] exu_io_next_bits_id2wb_regfile_we_addr; // @[EXU.scala 158:21]
  wire [38:0] exu_io_next_bits_ex2mem_addr; // @[EXU.scala 158:21]
  wire [63:0] exu_io_next_bits_ex2mem_we_data; // @[EXU.scala 158:21]
  wire [7:0] exu_io_next_bits_ex2mem_we_mask; // @[EXU.scala 158:21]
  wire [63:0] exu_io_next_bits_ex2wb_result_data; // @[EXU.scala 158:21]
  wire [63:0] exu_io_csr2ctrl_out_mepc; // @[EXU.scala 158:21]
  wire [63:0] exu_io_csr2ctrl_out_mtvec; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_mie; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_mtie; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_msie; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_meie; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_mtip; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_msip; // @[EXU.scala 158:21]
  wire  exu_io_csr2ctrl_out_meip; // @[EXU.scala 158:21]
  wire  exu_io_sb_clint_msip; // @[EXU.scala 158:21]
  wire  exu_io_sb_clint_mtip; // @[EXU.scala 158:21]
  wire [63:0] exu_io_sb_clint_mtime; // @[EXU.scala 158:21]
  wire  exu_io_sb_meip; // @[EXU.scala 158:21]
  wire  EX2MEMReg_clock; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_reset; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_ready; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_valid; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_fencei; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_size_byte; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_size_hword; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_size_word; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_size_dword; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_sext_flag; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_memory_rd_en; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2mem_memory_we_en; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2wb_intr_exce_ret; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2wb_fencei; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2wb_wb_sel; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_prev_bits_id2wb_regfile_we_en; // @[MEMU.scala 84:27]
  wire [4:0] EX2MEMReg_io_prev_bits_id2wb_regfile_we_addr; // @[MEMU.scala 84:27]
  wire [38:0] EX2MEMReg_io_prev_bits_ex2mem_addr; // @[MEMU.scala 84:27]
  wire [63:0] EX2MEMReg_io_prev_bits_ex2mem_we_data; // @[MEMU.scala 84:27]
  wire [7:0] EX2MEMReg_io_prev_bits_ex2mem_we_mask; // @[MEMU.scala 84:27]
  wire [63:0] EX2MEMReg_io_prev_bits_ex2wb_result_data; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_ready; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_valid; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_fencei; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_size_byte; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_size_hword; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_size_word; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_size_dword; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_sext_flag; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_memory_rd_en; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2mem_memory_we_en; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2wb_intr_exce_ret; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2wb_fencei; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2wb_wb_sel; // @[MEMU.scala 84:27]
  wire  EX2MEMReg_io_next_bits_id2wb_regfile_we_en; // @[MEMU.scala 84:27]
  wire [4:0] EX2MEMReg_io_next_bits_id2wb_regfile_we_addr; // @[MEMU.scala 84:27]
  wire [38:0] EX2MEMReg_io_next_bits_ex2mem_addr; // @[MEMU.scala 84:27]
  wire [63:0] EX2MEMReg_io_next_bits_ex2mem_we_data; // @[MEMU.scala 84:27]
  wire [7:0] EX2MEMReg_io_next_bits_ex2mem_we_mask; // @[MEMU.scala 84:27]
  wire [63:0] EX2MEMReg_io_next_bits_ex2wb_result_data; // @[MEMU.scala 84:27]
  wire  memu_clock; // @[MEMU.scala 87:22]
  wire  memu_reset; // @[MEMU.scala 87:22]
  wire  memu_io_prev_ready; // @[MEMU.scala 87:22]
  wire  memu_io_prev_valid; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_fencei; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_size_byte; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_size_hword; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_size_word; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_size_dword; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_sext_flag; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_memory_rd_en; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2mem_memory_we_en; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2wb_intr_exce_ret; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2wb_fencei; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2wb_wb_sel; // @[MEMU.scala 87:22]
  wire  memu_io_prev_bits_id2wb_regfile_we_en; // @[MEMU.scala 87:22]
  wire [4:0] memu_io_prev_bits_id2wb_regfile_we_addr; // @[MEMU.scala 87:22]
  wire [38:0] memu_io_prev_bits_ex2mem_addr; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_prev_bits_ex2mem_we_data; // @[MEMU.scala 87:22]
  wire [7:0] memu_io_prev_bits_ex2mem_we_mask; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_prev_bits_ex2wb_result_data; // @[MEMU.scala 87:22]
  wire  memu_io_next_valid; // @[MEMU.scala 87:22]
  wire  memu_io_next_bits_id2wb_intr_exce_ret; // @[MEMU.scala 87:22]
  wire  memu_io_next_bits_id2wb_fencei; // @[MEMU.scala 87:22]
  wire  memu_io_next_bits_id2wb_wb_sel; // @[MEMU.scala 87:22]
  wire  memu_io_next_bits_id2wb_regfile_we_en; // @[MEMU.scala 87:22]
  wire [4:0] memu_io_next_bits_id2wb_regfile_we_addr; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_next_bits_ex2wb_result_data; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_next_bits_mem2wb_memory_data; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_ar_ready; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_ar_valid; // @[MEMU.scala 87:22]
  wire [31:0] memu_io_maxi_ar_bits_addr; // @[MEMU.scala 87:22]
  wire [7:0] memu_io_maxi_ar_bits_len; // @[MEMU.scala 87:22]
  wire [2:0] memu_io_maxi_ar_bits_size; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_r_valid; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_maxi_r_bits_data; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_r_bits_last; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_aw_ready; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_aw_valid; // @[MEMU.scala 87:22]
  wire [31:0] memu_io_maxi_aw_bits_addr; // @[MEMU.scala 87:22]
  wire [7:0] memu_io_maxi_aw_bits_len; // @[MEMU.scala 87:22]
  wire [2:0] memu_io_maxi_aw_bits_size; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_w_ready; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_w_valid; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_maxi_w_bits_data; // @[MEMU.scala 87:22]
  wire [7:0] memu_io_maxi_w_bits_strb; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_w_bits_last; // @[MEMU.scala 87:22]
  wire  memu_io_maxi_b_valid; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_ar_ready; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_ar_valid; // @[MEMU.scala 87:22]
  wire [31:0] memu_io_mmio_ar_bits_addr; // @[MEMU.scala 87:22]
  wire [2:0] memu_io_mmio_ar_bits_size; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_r_valid; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_mmio_r_bits_data; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_r_bits_last; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_aw_ready; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_aw_valid; // @[MEMU.scala 87:22]
  wire [31:0] memu_io_mmio_aw_bits_addr; // @[MEMU.scala 87:22]
  wire [2:0] memu_io_mmio_aw_bits_size; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_w_ready; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_w_valid; // @[MEMU.scala 87:22]
  wire [63:0] memu_io_mmio_w_bits_data; // @[MEMU.scala 87:22]
  wire [7:0] memu_io_mmio_w_bits_strb; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_w_bits_last; // @[MEMU.scala 87:22]
  wire  memu_io_mmio_b_valid; // @[MEMU.scala 87:22]
  wire [5:0] memu_io_sram4_addr; // @[MEMU.scala 87:22]
  wire  memu_io_sram4_wen; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram4_wmask; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram4_wdata; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram4_rdata; // @[MEMU.scala 87:22]
  wire [5:0] memu_io_sram5_addr; // @[MEMU.scala 87:22]
  wire  memu_io_sram5_wen; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram5_wmask; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram5_wdata; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram5_rdata; // @[MEMU.scala 87:22]
  wire [5:0] memu_io_sram6_addr; // @[MEMU.scala 87:22]
  wire  memu_io_sram6_wen; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram6_wmask; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram6_wdata; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram6_rdata; // @[MEMU.scala 87:22]
  wire [5:0] memu_io_sram7_addr; // @[MEMU.scala 87:22]
  wire  memu_io_sram7_wen; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram7_wmask; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram7_wdata; // @[MEMU.scala 87:22]
  wire [127:0] memu_io_sram7_rdata; // @[MEMU.scala 87:22]
  wire  memu_clint_we; // @[MEMU.scala 87:22]
  wire [31:0] memu__T_24; // @[MEMU.scala 87:22]
  wire [63:0] memu_clint_rdata; // @[MEMU.scala 87:22]
  wire [63:0] memu_clint_wdata; // @[MEMU.scala 87:22]
  wire  MEM2WBReg_clock; // @[WBU.scala 77:27]
  wire  MEM2WBReg_reset; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_prev_valid; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_prev_bits_id2wb_intr_exce_ret; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_prev_bits_id2wb_fencei; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_prev_bits_id2wb_wb_sel; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_prev_bits_id2wb_regfile_we_en; // @[WBU.scala 77:27]
  wire [4:0] MEM2WBReg_io_prev_bits_id2wb_regfile_we_addr; // @[WBU.scala 77:27]
  wire [63:0] MEM2WBReg_io_prev_bits_ex2wb_result_data; // @[WBU.scala 77:27]
  wire [63:0] MEM2WBReg_io_prev_bits_mem2wb_memory_data; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_next_valid; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_next_bits_id2wb_intr_exce_ret; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_next_bits_id2wb_fencei; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_next_bits_id2wb_wb_sel; // @[WBU.scala 77:27]
  wire  MEM2WBReg_io_next_bits_id2wb_regfile_we_en; // @[WBU.scala 77:27]
  wire [4:0] MEM2WBReg_io_next_bits_id2wb_regfile_we_addr; // @[WBU.scala 77:27]
  wire [63:0] MEM2WBReg_io_next_bits_ex2wb_result_data; // @[WBU.scala 77:27]
  wire [63:0] MEM2WBReg_io_next_bits_mem2wb_memory_data; // @[WBU.scala 77:27]
  wire  wbu_io__prev_valid; // @[WBU.scala 80:21]
  wire  wbu_io__prev_bits_id2wb_intr_exce_ret; // @[WBU.scala 80:21]
  wire  wbu_io__prev_bits_id2wb_fencei; // @[WBU.scala 80:21]
  wire  wbu_io__prev_bits_id2wb_wb_sel; // @[WBU.scala 80:21]
  wire  wbu_io__prev_bits_id2wb_regfile_we_en; // @[WBU.scala 80:21]
  wire [4:0] wbu_io__prev_bits_id2wb_regfile_we_addr; // @[WBU.scala 80:21]
  wire [63:0] wbu_io__prev_bits_ex2wb_result_data; // @[WBU.scala 80:21]
  wire [63:0] wbu_io__prev_bits_mem2wb_memory_data; // @[WBU.scala 80:21]
  wire  wbu_io__regfile_en; // @[WBU.scala 80:21]
  wire [4:0] wbu_io__regfile_addr; // @[WBU.scala 80:21]
  wire [63:0] wbu_io__regfile_data; // @[WBU.scala 80:21]
  wire  wbu_io_prev_bits_id2wb_fencei; // @[WBU.scala 80:21]
  wire  wbu_io_prev_bits_id2wb_intr_exce_ret; // @[WBU.scala 80:21]
  wire [63:0] fwu_io_idu_fw_src1_data; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_idu_fw_src2_data; // @[FWU.scala 102:21]
  wire  fwu_io_idu_fw_ready; // @[FWU.scala 102:21]
  wire  fwu_io_idu_optype_Itype; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_idu_src1_addr; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_idu_src2_addr; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_idu_src1_data; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_idu_src2_data; // @[FWU.scala 102:21]
  wire  fwu_io_exu_is_load; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_exu_dst_addr; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_exu_dst_data; // @[FWU.scala 102:21]
  wire  fwu_io_memu_is_load_1; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_memu_dst_addr_1; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_memu_dst_data_1; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_memu_dst_addr_2; // @[FWU.scala 102:21]
  wire [4:0] fwu_io_wbu_dst_addr; // @[FWU.scala 102:21]
  wire [63:0] fwu_io_wbu_dst_data; // @[FWU.scala 102:21]
  wire  bru_clock; // @[BRU.scala 56:21]
  wire  bru_reset; // @[BRU.scala 56:21]
  wire  bru_io_idu_brh; // @[BRU.scala 56:21]
  wire  bru_io_idu_jal; // @[BRU.scala 56:21]
  wire  bru_io_idu_jalr; // @[BRU.scala 56:21]
  wire [63:0] bru_io_idu_pc; // @[BRU.scala 56:21]
  wire [63:0] bru_io_idu_src1; // @[BRU.scala 56:21]
  wire [63:0] bru_io_idu_src2; // @[BRU.scala 56:21]
  wire [63:0] bru_io_idu_imm; // @[BRU.scala 56:21]
  wire  bru_io_ifu_jump; // @[BRU.scala 56:21]
  wire [63:0] bru_io_ifu_npc; // @[BRU.scala 56:21]
  wire  bru_io_ifu_jump0; // @[BRU.scala 56:21]
  wire  regfile_clock; // @[Top.scala 53:31]
  wire  regfile_reset; // @[Top.scala 53:31]
  wire  regfile_io_wbu_en; // @[Top.scala 53:31]
  wire [4:0] regfile_io_wbu_addr; // @[Top.scala 53:31]
  wire [63:0] regfile_io_wbu_data; // @[Top.scala 53:31]
  wire [4:0] regfile_io_idu_addr1; // @[Top.scala 53:31]
  wire [63:0] regfile_io_idu_data1; // @[Top.scala 53:31]
  wire [4:0] regfile_io_idu_addr2; // @[Top.scala 53:31]
  wire [63:0] regfile_io_idu_data2; // @[Top.scala 53:31]
  reg  sram_init_reg; // @[Top.scala 42:38]
  reg [5:0] sram_init_cnt; // @[Counter.scala 60:40]
  wire  wrap_wrap = sram_init_cnt == 6'h3f; // @[Counter.scala 72:24]
  wire [5:0] _wrap_value_T_1 = sram_init_cnt + 6'h1; // @[Counter.scala 76:24]
  wire  BRIFBdl_jump = bru_io_ifu_jump; // @[Top.scala 23:29 BRU.scala 57:16]
  wire  IDUOut_ready = ID2EXReg_io_prev_ready; // @[Top.scala 26:29 EXU.scala 156:22]
  wire  IDFWBdl_fw_ready = fwu_io_idu_fw_ready; // @[Top.scala 29:29 FWU.scala 103:16]
  wire  _GEN_52 = wrap_wrap ? 1'h0 : sram_init_reg; // @[Top.scala 76:31 Top.scala 77:19 Top.scala 42:38]
  ysyx_040978_Interconnect3x1 icon ( // @[AXI.scala 285:30]
    .clock(icon_clock),
    .reset(icon_reset),
    .io_maxi_ar_ready(icon_io_maxi_ar_ready),
    .io_maxi_ar_valid(icon_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(icon_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_id(icon_io_maxi_ar_bits_id),
    .io_maxi_ar_bits_len(icon_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(icon_io_maxi_ar_bits_size),
    .io_maxi_r_valid(icon_io_maxi_r_valid),
    .io_maxi_r_bits_data(icon_io_maxi_r_bits_data),
    .io_maxi_r_bits_id(icon_io_maxi_r_bits_id),
    .io_maxi_r_bits_last(icon_io_maxi_r_bits_last),
    .io_maxi_aw_ready(icon_io_maxi_aw_ready),
    .io_maxi_aw_valid(icon_io_maxi_aw_valid),
    .io_maxi_aw_bits_addr(icon_io_maxi_aw_bits_addr),
    .io_maxi_aw_bits_id(icon_io_maxi_aw_bits_id),
    .io_maxi_aw_bits_len(icon_io_maxi_aw_bits_len),
    .io_maxi_aw_bits_size(icon_io_maxi_aw_bits_size),
    .io_maxi_w_ready(icon_io_maxi_w_ready),
    .io_maxi_w_valid(icon_io_maxi_w_valid),
    .io_maxi_w_bits_data(icon_io_maxi_w_bits_data),
    .io_maxi_w_bits_strb(icon_io_maxi_w_bits_strb),
    .io_maxi_w_bits_last(icon_io_maxi_w_bits_last),
    .io_maxi_b_valid(icon_io_maxi_b_valid),
    .io_maxi_b_bits_id(icon_io_maxi_b_bits_id),
    .io_ifu_ar_ready(icon_io_ifu_ar_ready),
    .io_ifu_ar_valid(icon_io_ifu_ar_valid),
    .io_ifu_ar_bits_addr(icon_io_ifu_ar_bits_addr),
    .io_ifu_ar_bits_len(icon_io_ifu_ar_bits_len),
    .io_ifu_ar_bits_size(icon_io_ifu_ar_bits_size),
    .io_ifu_r_valid(icon_io_ifu_r_valid),
    .io_ifu_r_bits_data(icon_io_ifu_r_bits_data),
    .io_ifu_r_bits_last(icon_io_ifu_r_bits_last),
    .io_memu_ar_ready(icon_io_memu_ar_ready),
    .io_memu_ar_valid(icon_io_memu_ar_valid),
    .io_memu_ar_bits_addr(icon_io_memu_ar_bits_addr),
    .io_memu_ar_bits_len(icon_io_memu_ar_bits_len),
    .io_memu_ar_bits_size(icon_io_memu_ar_bits_size),
    .io_memu_r_valid(icon_io_memu_r_valid),
    .io_memu_r_bits_data(icon_io_memu_r_bits_data),
    .io_memu_r_bits_last(icon_io_memu_r_bits_last),
    .io_memu_aw_ready(icon_io_memu_aw_ready),
    .io_memu_aw_valid(icon_io_memu_aw_valid),
    .io_memu_aw_bits_addr(icon_io_memu_aw_bits_addr),
    .io_memu_aw_bits_len(icon_io_memu_aw_bits_len),
    .io_memu_aw_bits_size(icon_io_memu_aw_bits_size),
    .io_memu_w_ready(icon_io_memu_w_ready),
    .io_memu_w_valid(icon_io_memu_w_valid),
    .io_memu_w_bits_data(icon_io_memu_w_bits_data),
    .io_memu_w_bits_strb(icon_io_memu_w_bits_strb),
    .io_memu_w_bits_last(icon_io_memu_w_bits_last),
    .io_memu_b_valid(icon_io_memu_b_valid),
    .io_devu_ar_ready(icon_io_devu_ar_ready),
    .io_devu_ar_valid(icon_io_devu_ar_valid),
    .io_devu_ar_bits_addr(icon_io_devu_ar_bits_addr),
    .io_devu_ar_bits_size(icon_io_devu_ar_bits_size),
    .io_devu_r_valid(icon_io_devu_r_valid),
    .io_devu_r_bits_data(icon_io_devu_r_bits_data),
    .io_devu_r_bits_last(icon_io_devu_r_bits_last),
    .io_devu_aw_ready(icon_io_devu_aw_ready),
    .io_devu_aw_valid(icon_io_devu_aw_valid),
    .io_devu_aw_bits_addr(icon_io_devu_aw_bits_addr),
    .io_devu_aw_bits_size(icon_io_devu_aw_bits_size),
    .io_devu_w_ready(icon_io_devu_w_ready),
    .io_devu_w_valid(icon_io_devu_w_valid),
    .io_devu_w_bits_data(icon_io_devu_w_bits_data),
    .io_devu_w_bits_strb(icon_io_devu_w_bits_strb),
    .io_devu_w_bits_last(icon_io_devu_w_bits_last),
    .io_devu_b_valid(icon_io_devu_b_valid)
  );
  ysyx_040978_PC pc ( // @[IFU.scala 96:20]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_jump0(pc_io_jump0),
    .io_jump(pc_io_jump),
    .io_npc(pc_io_npc),
    .io_sys_ready(pc_io_sys_ready),
    .io_next_ready(pc_io_next_ready),
    .io_next_valid(pc_io_next_valid),
    .io_next_bits_pc2if_pc(pc_io_next_bits_pc2if_pc)
  );
  ysyx_040978_IFU ifu ( // @[IFU.scala 102:21]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_cache_reset(ifu_io_cache_reset),
    .io_prev_ready(ifu_io_prev_ready),
    .io_prev_valid(ifu_io_prev_valid),
    .io_prev_bits_pc2if_pc(ifu_io_prev_bits_pc2if_pc),
    .io_maxi_ar_ready(ifu_io_maxi_ar_ready),
    .io_maxi_ar_valid(ifu_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(ifu_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(ifu_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(ifu_io_maxi_ar_bits_size),
    .io_maxi_r_valid(ifu_io_maxi_r_valid),
    .io_maxi_r_bits_data(ifu_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(ifu_io_maxi_r_bits_last),
    .io_next_ready(ifu_io_next_ready),
    .io_next_valid(ifu_io_next_valid),
    .io_next_bits_if2id_inst(ifu_io_next_bits_if2id_inst),
    .io_next_bits_if2id_pc(ifu_io_next_bits_if2id_pc),
    .io_sram0_addr(ifu_io_sram0_addr),
    .io_sram0_wen(ifu_io_sram0_wen),
    .io_sram0_wmask(ifu_io_sram0_wmask),
    .io_sram0_wdata(ifu_io_sram0_wdata),
    .io_sram0_rdata(ifu_io_sram0_rdata),
    .io_sram1_addr(ifu_io_sram1_addr),
    .io_sram1_wen(ifu_io_sram1_wen),
    .io_sram1_wmask(ifu_io_sram1_wmask),
    .io_sram1_wdata(ifu_io_sram1_wdata),
    .io_sram1_rdata(ifu_io_sram1_rdata),
    .io_sram2_addr(ifu_io_sram2_addr),
    .io_sram2_wen(ifu_io_sram2_wen),
    .io_sram2_wmask(ifu_io_sram2_wmask),
    .io_sram2_wdata(ifu_io_sram2_wdata),
    .io_sram2_rdata(ifu_io_sram2_rdata),
    .io_sram3_addr(ifu_io_sram3_addr),
    .io_sram3_wen(ifu_io_sram3_wen),
    .io_sram3_wmask(ifu_io_sram3_wmask),
    .io_sram3_wdata(ifu_io_sram3_wdata),
    .io_sram3_rdata(ifu_io_sram3_rdata),
    .fenceiing(ifu_fenceiing)
  );
  ysyx_040978_IDReg IF2IDReg ( // @[IDU.scala 286:26]
    .clock(IF2IDReg_clock),
    .reset(IF2IDReg_reset),
    .io_prev_ready(IF2IDReg_io_prev_ready),
    .io_prev_valid(IF2IDReg_io_prev_valid),
    .io_prev_bits_if2id_inst(IF2IDReg_io_prev_bits_if2id_inst),
    .io_prev_bits_if2id_pc(IF2IDReg_io_prev_bits_if2id_pc),
    .io_next_ready(IF2IDReg_io_next_ready),
    .io_next_valid(IF2IDReg_io_next_valid),
    .io_next_bits_if2id_inst(IF2IDReg_io_next_bits_if2id_inst),
    .io_next_bits_if2id_pc(IF2IDReg_io_next_bits_if2id_pc)
  );
  ysyx_040978_IDU idu ( // @[IDU.scala 290:21]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_regfile_addr1(idu_io_regfile_addr1),
    .io_regfile_data1(idu_io_regfile_data1),
    .io_regfile_addr2(idu_io_regfile_addr2),
    .io_regfile_data2(idu_io_regfile_data2),
    .io_fwu_fw_src1_data(idu_io_fwu_fw_src1_data),
    .io_fwu_fw_src2_data(idu_io_fwu_fw_src2_data),
    .io_fwu_optype_Itype(idu_io_fwu_optype_Itype),
    .io_fwu_src1_addr(idu_io_fwu_src1_addr),
    .io_fwu_src2_addr(idu_io_fwu_src2_addr),
    .io_fwu_src1_data(idu_io_fwu_src1_data),
    .io_fwu_src2_data(idu_io_fwu_src2_data),
    .io_bru_brh(idu_io_bru_brh),
    .io_bru_jal(idu_io_bru_jal),
    .io_bru_jalr(idu_io_bru_jalr),
    .io_bru_pc(idu_io_bru_pc),
    .io_bru_src1(idu_io_bru_src1),
    .io_bru_src2(idu_io_bru_src2),
    .io_bru_imm(idu_io_bru_imm),
    .io_csr_out_mepc(idu_io_csr_out_mepc),
    .io_csr_out_mtvec(idu_io_csr_out_mtvec),
    .io_csr_out_mie(idu_io_csr_out_mie),
    .io_csr_out_mtie(idu_io_csr_out_mtie),
    .io_csr_out_msie(idu_io_csr_out_msie),
    .io_csr_out_meie(idu_io_csr_out_meie),
    .io_csr_out_mtip(idu_io_csr_out_mtip),
    .io_csr_out_msip(idu_io_csr_out_msip),
    .io_csr_out_meip(idu_io_csr_out_meip),
    .io_prev_ready(idu_io_prev_ready),
    .io_prev_valid(idu_io_prev_valid),
    .io_prev_bits_if2id_inst(idu_io_prev_bits_if2id_inst),
    .io_prev_bits_if2id_pc(idu_io_prev_bits_if2id_pc),
    .io_next_ready(idu_io_next_ready),
    .io_next_valid(idu_io_next_valid),
    .io_next_bits_id2ex_alu_src1(idu_io_next_bits_id2ex_alu_src1),
    .io_next_bits_id2ex_alu_src2(idu_io_next_bits_id2ex_alu_src2),
    .io_next_bits_id2ex_salu_src1(idu_io_next_bits_id2ex_salu_src1),
    .io_next_bits_id2ex_salu_src2(idu_io_next_bits_id2ex_salu_src2),
    .io_next_bits_id2ex_src1(idu_io_next_bits_id2ex_src1),
    .io_next_bits_id2ex_src2(idu_io_next_bits_id2ex_src2),
    .io_next_bits_id2ex_src3(idu_io_next_bits_id2ex_src3),
    .io_next_bits_id2ex_operator_auipc(idu_io_next_bits_id2ex_operator_auipc),
    .io_next_bits_id2ex_operator_lui(idu_io_next_bits_id2ex_operator_lui),
    .io_next_bits_id2ex_operator_jal(idu_io_next_bits_id2ex_operator_jal),
    .io_next_bits_id2ex_operator_jalr(idu_io_next_bits_id2ex_operator_jalr),
    .io_next_bits_id2ex_operator_sb(idu_io_next_bits_id2ex_operator_sb),
    .io_next_bits_id2ex_operator_sh(idu_io_next_bits_id2ex_operator_sh),
    .io_next_bits_id2ex_operator_sw(idu_io_next_bits_id2ex_operator_sw),
    .io_next_bits_id2ex_operator_sd(idu_io_next_bits_id2ex_operator_sd),
    .io_next_bits_id2ex_operator_add(idu_io_next_bits_id2ex_operator_add),
    .io_next_bits_id2ex_operator_sub(idu_io_next_bits_id2ex_operator_sub),
    .io_next_bits_id2ex_operator_sll(idu_io_next_bits_id2ex_operator_sll),
    .io_next_bits_id2ex_operator_slt(idu_io_next_bits_id2ex_operator_slt),
    .io_next_bits_id2ex_operator_sltu(idu_io_next_bits_id2ex_operator_sltu),
    .io_next_bits_id2ex_operator_xor(idu_io_next_bits_id2ex_operator_xor),
    .io_next_bits_id2ex_operator_srl(idu_io_next_bits_id2ex_operator_srl),
    .io_next_bits_id2ex_operator_sra(idu_io_next_bits_id2ex_operator_sra),
    .io_next_bits_id2ex_operator_or(idu_io_next_bits_id2ex_operator_or),
    .io_next_bits_id2ex_operator_and(idu_io_next_bits_id2ex_operator_and),
    .io_next_bits_id2ex_operator_csr_is_csr(idu_io_next_bits_id2ex_operator_csr_is_csr),
    .io_next_bits_id2ex_operator_csr_csrrw(idu_io_next_bits_id2ex_operator_csr_csrrw),
    .io_next_bits_id2ex_operator_csr_csrrs(idu_io_next_bits_id2ex_operator_csr_csrrs),
    .io_next_bits_id2ex_operator_csr_csrrc(idu_io_next_bits_id2ex_operator_csr_csrrc),
    .io_next_bits_id2ex_operator_csr_csrrwi(idu_io_next_bits_id2ex_operator_csr_csrrwi),
    .io_next_bits_id2ex_operator_csr_csrrsi(idu_io_next_bits_id2ex_operator_csr_csrrsi),
    .io_next_bits_id2ex_operator_csr_csrrci(idu_io_next_bits_id2ex_operator_csr_csrrci),
    .io_next_bits_id2ex_srcsize_byte(idu_io_next_bits_id2ex_srcsize_byte),
    .io_next_bits_id2ex_srcsize_hword(idu_io_next_bits_id2ex_srcsize_hword),
    .io_next_bits_id2ex_srcsize_word(idu_io_next_bits_id2ex_srcsize_word),
    .io_next_bits_id2ex_srcsize_dword(idu_io_next_bits_id2ex_srcsize_dword),
    .io_next_bits_id2ex_is_load(idu_io_next_bits_id2ex_is_load),
    .io_next_bits_id2ex_is_save(idu_io_next_bits_id2ex_is_save),
    .io_next_bits_id2ex_div_inf(idu_io_next_bits_id2ex_div_inf),
    .io_next_bits_id2ex_csr_we(idu_io_next_bits_id2ex_csr_we),
    .io_next_bits_id2ex_csr_hit_is_mepc(idu_io_next_bits_id2ex_csr_hit_is_mepc),
    .io_next_bits_id2ex_csr_hit_is_mtvec(idu_io_next_bits_id2ex_csr_hit_is_mtvec),
    .io_next_bits_id2ex_csr_hit_is_mstatus(idu_io_next_bits_id2ex_csr_hit_is_mstatus),
    .io_next_bits_id2ex_csr_hit_is_mie(idu_io_next_bits_id2ex_csr_hit_is_mie),
    .io_next_bits_id2ex_csr_hit_is_mcause(idu_io_next_bits_id2ex_csr_hit_is_mcause),
    .io_next_bits_id2ex_csr_hit_is_mip(idu_io_next_bits_id2ex_csr_hit_is_mip),
    .io_next_bits_id2ex_csr_hit_is_mtime(idu_io_next_bits_id2ex_csr_hit_is_mtime),
    .io_next_bits_id2ex_csr_hit_is_mcycle(idu_io_next_bits_id2ex_csr_hit_is_mcycle),
    .io_next_bits_id2ex_csr_hit_is_mhartid(idu_io_next_bits_id2ex_csr_hit_is_mhartid),
    .io_next_bits_id2ex_mdu_op_mul_signed(idu_io_next_bits_id2ex_mdu_op_mul_signed),
    .io_next_bits_id2ex_mdu_op_is_mu(idu_io_next_bits_id2ex_mdu_op_is_mu),
    .io_next_bits_id2ex_mdu_op_mul_32(idu_io_next_bits_id2ex_mdu_op_mul_32),
    .io_next_bits_id2ex_mdu_op_div_signed(idu_io_next_bits_id2ex_mdu_op_div_signed),
    .io_next_bits_id2ex_mdu_op_is_div(idu_io_next_bits_id2ex_mdu_op_is_div),
    .io_next_bits_id2ex_mdu_op_is_du(idu_io_next_bits_id2ex_mdu_op_is_du),
    .io_next_bits_id2ex_zimm(idu_io_next_bits_id2ex_zimm),
    .io_next_bits_id2ex_intr(idu_io_next_bits_id2ex_intr),
    .io_next_bits_id2ex_exec(idu_io_next_bits_id2ex_exec),
    .io_next_bits_id2ex_mret(idu_io_next_bits_id2ex_mret),
    .io_next_bits_id2ex_exce_code(idu_io_next_bits_id2ex_exce_code),
    .io_next_bits_id2ex_pc(idu_io_next_bits_id2ex_pc),
    .io_next_bits_id2ex_is_iem(idu_io_next_bits_id2ex_is_iem),
    .io_next_bits_id2mem_fencei(idu_io_next_bits_id2mem_fencei),
    .io_next_bits_id2mem_size_byte(idu_io_next_bits_id2mem_size_byte),
    .io_next_bits_id2mem_size_hword(idu_io_next_bits_id2mem_size_hword),
    .io_next_bits_id2mem_size_word(idu_io_next_bits_id2mem_size_word),
    .io_next_bits_id2mem_size_dword(idu_io_next_bits_id2mem_size_dword),
    .io_next_bits_id2mem_sext_flag(idu_io_next_bits_id2mem_sext_flag),
    .io_next_bits_id2mem_memory_rd_en(idu_io_next_bits_id2mem_memory_rd_en),
    .io_next_bits_id2mem_memory_we_en(idu_io_next_bits_id2mem_memory_we_en),
    .io_next_bits_id2wb_intr_exce_ret(idu_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(idu_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(idu_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(idu_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(idu_io_next_bits_id2wb_regfile_we_addr),
    .wb_fencei_0(idu_wb_fencei_0),
    .wb_intr_exce_ret_0(idu_wb_intr_exce_ret_0),
    .fenceiing_0(idu_fenceiing_0)
  );
  ysyx_040978_EXReg ID2EXReg ( // @[EXU.scala 155:26]
    .clock(ID2EXReg_clock),
    .reset(ID2EXReg_reset),
    .io_prev_ready(ID2EXReg_io_prev_ready),
    .io_prev_valid(ID2EXReg_io_prev_valid),
    .io_prev_bits_id2ex_alu_src1(ID2EXReg_io_prev_bits_id2ex_alu_src1),
    .io_prev_bits_id2ex_alu_src2(ID2EXReg_io_prev_bits_id2ex_alu_src2),
    .io_prev_bits_id2ex_salu_src1(ID2EXReg_io_prev_bits_id2ex_salu_src1),
    .io_prev_bits_id2ex_salu_src2(ID2EXReg_io_prev_bits_id2ex_salu_src2),
    .io_prev_bits_id2ex_src1(ID2EXReg_io_prev_bits_id2ex_src1),
    .io_prev_bits_id2ex_src2(ID2EXReg_io_prev_bits_id2ex_src2),
    .io_prev_bits_id2ex_src3(ID2EXReg_io_prev_bits_id2ex_src3),
    .io_prev_bits_id2ex_operator_auipc(ID2EXReg_io_prev_bits_id2ex_operator_auipc),
    .io_prev_bits_id2ex_operator_lui(ID2EXReg_io_prev_bits_id2ex_operator_lui),
    .io_prev_bits_id2ex_operator_jal(ID2EXReg_io_prev_bits_id2ex_operator_jal),
    .io_prev_bits_id2ex_operator_jalr(ID2EXReg_io_prev_bits_id2ex_operator_jalr),
    .io_prev_bits_id2ex_operator_sb(ID2EXReg_io_prev_bits_id2ex_operator_sb),
    .io_prev_bits_id2ex_operator_sh(ID2EXReg_io_prev_bits_id2ex_operator_sh),
    .io_prev_bits_id2ex_operator_sw(ID2EXReg_io_prev_bits_id2ex_operator_sw),
    .io_prev_bits_id2ex_operator_sd(ID2EXReg_io_prev_bits_id2ex_operator_sd),
    .io_prev_bits_id2ex_operator_add(ID2EXReg_io_prev_bits_id2ex_operator_add),
    .io_prev_bits_id2ex_operator_sub(ID2EXReg_io_prev_bits_id2ex_operator_sub),
    .io_prev_bits_id2ex_operator_sll(ID2EXReg_io_prev_bits_id2ex_operator_sll),
    .io_prev_bits_id2ex_operator_slt(ID2EXReg_io_prev_bits_id2ex_operator_slt),
    .io_prev_bits_id2ex_operator_sltu(ID2EXReg_io_prev_bits_id2ex_operator_sltu),
    .io_prev_bits_id2ex_operator_xor(ID2EXReg_io_prev_bits_id2ex_operator_xor),
    .io_prev_bits_id2ex_operator_srl(ID2EXReg_io_prev_bits_id2ex_operator_srl),
    .io_prev_bits_id2ex_operator_sra(ID2EXReg_io_prev_bits_id2ex_operator_sra),
    .io_prev_bits_id2ex_operator_or(ID2EXReg_io_prev_bits_id2ex_operator_or),
    .io_prev_bits_id2ex_operator_and(ID2EXReg_io_prev_bits_id2ex_operator_and),
    .io_prev_bits_id2ex_operator_csr_is_csr(ID2EXReg_io_prev_bits_id2ex_operator_csr_is_csr),
    .io_prev_bits_id2ex_operator_csr_csrrw(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrw),
    .io_prev_bits_id2ex_operator_csr_csrrs(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrs),
    .io_prev_bits_id2ex_operator_csr_csrrc(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrc),
    .io_prev_bits_id2ex_operator_csr_csrrwi(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrwi),
    .io_prev_bits_id2ex_operator_csr_csrrsi(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrsi),
    .io_prev_bits_id2ex_operator_csr_csrrci(ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrci),
    .io_prev_bits_id2ex_srcsize_byte(ID2EXReg_io_prev_bits_id2ex_srcsize_byte),
    .io_prev_bits_id2ex_srcsize_hword(ID2EXReg_io_prev_bits_id2ex_srcsize_hword),
    .io_prev_bits_id2ex_srcsize_word(ID2EXReg_io_prev_bits_id2ex_srcsize_word),
    .io_prev_bits_id2ex_srcsize_dword(ID2EXReg_io_prev_bits_id2ex_srcsize_dword),
    .io_prev_bits_id2ex_is_load(ID2EXReg_io_prev_bits_id2ex_is_load),
    .io_prev_bits_id2ex_is_save(ID2EXReg_io_prev_bits_id2ex_is_save),
    .io_prev_bits_id2ex_div_inf(ID2EXReg_io_prev_bits_id2ex_div_inf),
    .io_prev_bits_id2ex_csr_we(ID2EXReg_io_prev_bits_id2ex_csr_we),
    .io_prev_bits_id2ex_csr_hit_is_mepc(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mepc),
    .io_prev_bits_id2ex_csr_hit_is_mtvec(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtvec),
    .io_prev_bits_id2ex_csr_hit_is_mstatus(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mstatus),
    .io_prev_bits_id2ex_csr_hit_is_mie(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mie),
    .io_prev_bits_id2ex_csr_hit_is_mcause(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcause),
    .io_prev_bits_id2ex_csr_hit_is_mip(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mip),
    .io_prev_bits_id2ex_csr_hit_is_mtime(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtime),
    .io_prev_bits_id2ex_csr_hit_is_mcycle(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcycle),
    .io_prev_bits_id2ex_csr_hit_is_mhartid(ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mhartid),
    .io_prev_bits_id2ex_mdu_op_mul_signed(ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_signed),
    .io_prev_bits_id2ex_mdu_op_is_mu(ID2EXReg_io_prev_bits_id2ex_mdu_op_is_mu),
    .io_prev_bits_id2ex_mdu_op_mul_32(ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_32),
    .io_prev_bits_id2ex_mdu_op_div_signed(ID2EXReg_io_prev_bits_id2ex_mdu_op_div_signed),
    .io_prev_bits_id2ex_mdu_op_is_div(ID2EXReg_io_prev_bits_id2ex_mdu_op_is_div),
    .io_prev_bits_id2ex_mdu_op_is_du(ID2EXReg_io_prev_bits_id2ex_mdu_op_is_du),
    .io_prev_bits_id2ex_zimm(ID2EXReg_io_prev_bits_id2ex_zimm),
    .io_prev_bits_id2ex_intr(ID2EXReg_io_prev_bits_id2ex_intr),
    .io_prev_bits_id2ex_exec(ID2EXReg_io_prev_bits_id2ex_exec),
    .io_prev_bits_id2ex_mret(ID2EXReg_io_prev_bits_id2ex_mret),
    .io_prev_bits_id2ex_exce_code(ID2EXReg_io_prev_bits_id2ex_exce_code),
    .io_prev_bits_id2ex_pc(ID2EXReg_io_prev_bits_id2ex_pc),
    .io_prev_bits_id2ex_is_iem(ID2EXReg_io_prev_bits_id2ex_is_iem),
    .io_prev_bits_id2mem_fencei(ID2EXReg_io_prev_bits_id2mem_fencei),
    .io_prev_bits_id2mem_size_byte(ID2EXReg_io_prev_bits_id2mem_size_byte),
    .io_prev_bits_id2mem_size_hword(ID2EXReg_io_prev_bits_id2mem_size_hword),
    .io_prev_bits_id2mem_size_word(ID2EXReg_io_prev_bits_id2mem_size_word),
    .io_prev_bits_id2mem_size_dword(ID2EXReg_io_prev_bits_id2mem_size_dword),
    .io_prev_bits_id2mem_sext_flag(ID2EXReg_io_prev_bits_id2mem_sext_flag),
    .io_prev_bits_id2mem_memory_rd_en(ID2EXReg_io_prev_bits_id2mem_memory_rd_en),
    .io_prev_bits_id2mem_memory_we_en(ID2EXReg_io_prev_bits_id2mem_memory_we_en),
    .io_prev_bits_id2wb_intr_exce_ret(ID2EXReg_io_prev_bits_id2wb_intr_exce_ret),
    .io_prev_bits_id2wb_fencei(ID2EXReg_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_wb_sel(ID2EXReg_io_prev_bits_id2wb_wb_sel),
    .io_prev_bits_id2wb_regfile_we_en(ID2EXReg_io_prev_bits_id2wb_regfile_we_en),
    .io_prev_bits_id2wb_regfile_we_addr(ID2EXReg_io_prev_bits_id2wb_regfile_we_addr),
    .io_next_ready(ID2EXReg_io_next_ready),
    .io_next_valid(ID2EXReg_io_next_valid),
    .io_next_bits_id2ex_alu_src1(ID2EXReg_io_next_bits_id2ex_alu_src1),
    .io_next_bits_id2ex_alu_src2(ID2EXReg_io_next_bits_id2ex_alu_src2),
    .io_next_bits_id2ex_salu_src1(ID2EXReg_io_next_bits_id2ex_salu_src1),
    .io_next_bits_id2ex_salu_src2(ID2EXReg_io_next_bits_id2ex_salu_src2),
    .io_next_bits_id2ex_src1(ID2EXReg_io_next_bits_id2ex_src1),
    .io_next_bits_id2ex_src2(ID2EXReg_io_next_bits_id2ex_src2),
    .io_next_bits_id2ex_src3(ID2EXReg_io_next_bits_id2ex_src3),
    .io_next_bits_id2ex_operator_auipc(ID2EXReg_io_next_bits_id2ex_operator_auipc),
    .io_next_bits_id2ex_operator_lui(ID2EXReg_io_next_bits_id2ex_operator_lui),
    .io_next_bits_id2ex_operator_jal(ID2EXReg_io_next_bits_id2ex_operator_jal),
    .io_next_bits_id2ex_operator_jalr(ID2EXReg_io_next_bits_id2ex_operator_jalr),
    .io_next_bits_id2ex_operator_sb(ID2EXReg_io_next_bits_id2ex_operator_sb),
    .io_next_bits_id2ex_operator_sh(ID2EXReg_io_next_bits_id2ex_operator_sh),
    .io_next_bits_id2ex_operator_sw(ID2EXReg_io_next_bits_id2ex_operator_sw),
    .io_next_bits_id2ex_operator_sd(ID2EXReg_io_next_bits_id2ex_operator_sd),
    .io_next_bits_id2ex_operator_add(ID2EXReg_io_next_bits_id2ex_operator_add),
    .io_next_bits_id2ex_operator_sub(ID2EXReg_io_next_bits_id2ex_operator_sub),
    .io_next_bits_id2ex_operator_sll(ID2EXReg_io_next_bits_id2ex_operator_sll),
    .io_next_bits_id2ex_operator_slt(ID2EXReg_io_next_bits_id2ex_operator_slt),
    .io_next_bits_id2ex_operator_sltu(ID2EXReg_io_next_bits_id2ex_operator_sltu),
    .io_next_bits_id2ex_operator_xor(ID2EXReg_io_next_bits_id2ex_operator_xor),
    .io_next_bits_id2ex_operator_srl(ID2EXReg_io_next_bits_id2ex_operator_srl),
    .io_next_bits_id2ex_operator_sra(ID2EXReg_io_next_bits_id2ex_operator_sra),
    .io_next_bits_id2ex_operator_or(ID2EXReg_io_next_bits_id2ex_operator_or),
    .io_next_bits_id2ex_operator_and(ID2EXReg_io_next_bits_id2ex_operator_and),
    .io_next_bits_id2ex_operator_csr_is_csr(ID2EXReg_io_next_bits_id2ex_operator_csr_is_csr),
    .io_next_bits_id2ex_operator_csr_csrrw(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrw),
    .io_next_bits_id2ex_operator_csr_csrrs(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrs),
    .io_next_bits_id2ex_operator_csr_csrrc(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrc),
    .io_next_bits_id2ex_operator_csr_csrrwi(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrwi),
    .io_next_bits_id2ex_operator_csr_csrrsi(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrsi),
    .io_next_bits_id2ex_operator_csr_csrrci(ID2EXReg_io_next_bits_id2ex_operator_csr_csrrci),
    .io_next_bits_id2ex_srcsize_byte(ID2EXReg_io_next_bits_id2ex_srcsize_byte),
    .io_next_bits_id2ex_srcsize_hword(ID2EXReg_io_next_bits_id2ex_srcsize_hword),
    .io_next_bits_id2ex_srcsize_word(ID2EXReg_io_next_bits_id2ex_srcsize_word),
    .io_next_bits_id2ex_srcsize_dword(ID2EXReg_io_next_bits_id2ex_srcsize_dword),
    .io_next_bits_id2ex_is_load(ID2EXReg_io_next_bits_id2ex_is_load),
    .io_next_bits_id2ex_is_save(ID2EXReg_io_next_bits_id2ex_is_save),
    .io_next_bits_id2ex_div_inf(ID2EXReg_io_next_bits_id2ex_div_inf),
    .io_next_bits_id2ex_csr_we(ID2EXReg_io_next_bits_id2ex_csr_we),
    .io_next_bits_id2ex_csr_hit_is_mepc(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mepc),
    .io_next_bits_id2ex_csr_hit_is_mtvec(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtvec),
    .io_next_bits_id2ex_csr_hit_is_mstatus(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mstatus),
    .io_next_bits_id2ex_csr_hit_is_mie(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mie),
    .io_next_bits_id2ex_csr_hit_is_mcause(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcause),
    .io_next_bits_id2ex_csr_hit_is_mip(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mip),
    .io_next_bits_id2ex_csr_hit_is_mtime(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtime),
    .io_next_bits_id2ex_csr_hit_is_mcycle(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcycle),
    .io_next_bits_id2ex_csr_hit_is_mhartid(ID2EXReg_io_next_bits_id2ex_csr_hit_is_mhartid),
    .io_next_bits_id2ex_mdu_op_mul_signed(ID2EXReg_io_next_bits_id2ex_mdu_op_mul_signed),
    .io_next_bits_id2ex_mdu_op_is_mu(ID2EXReg_io_next_bits_id2ex_mdu_op_is_mu),
    .io_next_bits_id2ex_mdu_op_mul_32(ID2EXReg_io_next_bits_id2ex_mdu_op_mul_32),
    .io_next_bits_id2ex_mdu_op_div_signed(ID2EXReg_io_next_bits_id2ex_mdu_op_div_signed),
    .io_next_bits_id2ex_mdu_op_is_div(ID2EXReg_io_next_bits_id2ex_mdu_op_is_div),
    .io_next_bits_id2ex_mdu_op_is_du(ID2EXReg_io_next_bits_id2ex_mdu_op_is_du),
    .io_next_bits_id2ex_zimm(ID2EXReg_io_next_bits_id2ex_zimm),
    .io_next_bits_id2ex_intr(ID2EXReg_io_next_bits_id2ex_intr),
    .io_next_bits_id2ex_exec(ID2EXReg_io_next_bits_id2ex_exec),
    .io_next_bits_id2ex_mret(ID2EXReg_io_next_bits_id2ex_mret),
    .io_next_bits_id2ex_exce_code(ID2EXReg_io_next_bits_id2ex_exce_code),
    .io_next_bits_id2ex_pc(ID2EXReg_io_next_bits_id2ex_pc),
    .io_next_bits_id2ex_is_iem(ID2EXReg_io_next_bits_id2ex_is_iem),
    .io_next_bits_id2mem_fencei(ID2EXReg_io_next_bits_id2mem_fencei),
    .io_next_bits_id2mem_size_byte(ID2EXReg_io_next_bits_id2mem_size_byte),
    .io_next_bits_id2mem_size_hword(ID2EXReg_io_next_bits_id2mem_size_hword),
    .io_next_bits_id2mem_size_word(ID2EXReg_io_next_bits_id2mem_size_word),
    .io_next_bits_id2mem_size_dword(ID2EXReg_io_next_bits_id2mem_size_dword),
    .io_next_bits_id2mem_sext_flag(ID2EXReg_io_next_bits_id2mem_sext_flag),
    .io_next_bits_id2mem_memory_rd_en(ID2EXReg_io_next_bits_id2mem_memory_rd_en),
    .io_next_bits_id2mem_memory_we_en(ID2EXReg_io_next_bits_id2mem_memory_we_en),
    .io_next_bits_id2wb_intr_exce_ret(ID2EXReg_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(ID2EXReg_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(ID2EXReg_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(ID2EXReg_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(ID2EXReg_io_next_bits_id2wb_regfile_we_addr)
  );
  ysyx_040978_EXU exu ( // @[EXU.scala 158:21]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_prev_ready(exu_io_prev_ready),
    .io_prev_valid(exu_io_prev_valid),
    .io_prev_bits_id2ex_alu_src1(exu_io_prev_bits_id2ex_alu_src1),
    .io_prev_bits_id2ex_alu_src2(exu_io_prev_bits_id2ex_alu_src2),
    .io_prev_bits_id2ex_salu_src1(exu_io_prev_bits_id2ex_salu_src1),
    .io_prev_bits_id2ex_salu_src2(exu_io_prev_bits_id2ex_salu_src2),
    .io_prev_bits_id2ex_src1(exu_io_prev_bits_id2ex_src1),
    .io_prev_bits_id2ex_src2(exu_io_prev_bits_id2ex_src2),
    .io_prev_bits_id2ex_src3(exu_io_prev_bits_id2ex_src3),
    .io_prev_bits_id2ex_operator_auipc(exu_io_prev_bits_id2ex_operator_auipc),
    .io_prev_bits_id2ex_operator_lui(exu_io_prev_bits_id2ex_operator_lui),
    .io_prev_bits_id2ex_operator_jal(exu_io_prev_bits_id2ex_operator_jal),
    .io_prev_bits_id2ex_operator_jalr(exu_io_prev_bits_id2ex_operator_jalr),
    .io_prev_bits_id2ex_operator_sb(exu_io_prev_bits_id2ex_operator_sb),
    .io_prev_bits_id2ex_operator_sh(exu_io_prev_bits_id2ex_operator_sh),
    .io_prev_bits_id2ex_operator_sw(exu_io_prev_bits_id2ex_operator_sw),
    .io_prev_bits_id2ex_operator_sd(exu_io_prev_bits_id2ex_operator_sd),
    .io_prev_bits_id2ex_operator_add(exu_io_prev_bits_id2ex_operator_add),
    .io_prev_bits_id2ex_operator_sub(exu_io_prev_bits_id2ex_operator_sub),
    .io_prev_bits_id2ex_operator_sll(exu_io_prev_bits_id2ex_operator_sll),
    .io_prev_bits_id2ex_operator_slt(exu_io_prev_bits_id2ex_operator_slt),
    .io_prev_bits_id2ex_operator_sltu(exu_io_prev_bits_id2ex_operator_sltu),
    .io_prev_bits_id2ex_operator_xor(exu_io_prev_bits_id2ex_operator_xor),
    .io_prev_bits_id2ex_operator_srl(exu_io_prev_bits_id2ex_operator_srl),
    .io_prev_bits_id2ex_operator_sra(exu_io_prev_bits_id2ex_operator_sra),
    .io_prev_bits_id2ex_operator_or(exu_io_prev_bits_id2ex_operator_or),
    .io_prev_bits_id2ex_operator_and(exu_io_prev_bits_id2ex_operator_and),
    .io_prev_bits_id2ex_operator_csr_is_csr(exu_io_prev_bits_id2ex_operator_csr_is_csr),
    .io_prev_bits_id2ex_operator_csr_csrrw(exu_io_prev_bits_id2ex_operator_csr_csrrw),
    .io_prev_bits_id2ex_operator_csr_csrrs(exu_io_prev_bits_id2ex_operator_csr_csrrs),
    .io_prev_bits_id2ex_operator_csr_csrrc(exu_io_prev_bits_id2ex_operator_csr_csrrc),
    .io_prev_bits_id2ex_operator_csr_csrrwi(exu_io_prev_bits_id2ex_operator_csr_csrrwi),
    .io_prev_bits_id2ex_operator_csr_csrrsi(exu_io_prev_bits_id2ex_operator_csr_csrrsi),
    .io_prev_bits_id2ex_operator_csr_csrrci(exu_io_prev_bits_id2ex_operator_csr_csrrci),
    .io_prev_bits_id2ex_srcsize_byte(exu_io_prev_bits_id2ex_srcsize_byte),
    .io_prev_bits_id2ex_srcsize_hword(exu_io_prev_bits_id2ex_srcsize_hword),
    .io_prev_bits_id2ex_srcsize_word(exu_io_prev_bits_id2ex_srcsize_word),
    .io_prev_bits_id2ex_srcsize_dword(exu_io_prev_bits_id2ex_srcsize_dword),
    .io_prev_bits_id2ex_is_load(exu_io_prev_bits_id2ex_is_load),
    .io_prev_bits_id2ex_is_save(exu_io_prev_bits_id2ex_is_save),
    .io_prev_bits_id2ex_div_inf(exu_io_prev_bits_id2ex_div_inf),
    .io_prev_bits_id2ex_csr_we(exu_io_prev_bits_id2ex_csr_we),
    .io_prev_bits_id2ex_csr_hit_is_mepc(exu_io_prev_bits_id2ex_csr_hit_is_mepc),
    .io_prev_bits_id2ex_csr_hit_is_mtvec(exu_io_prev_bits_id2ex_csr_hit_is_mtvec),
    .io_prev_bits_id2ex_csr_hit_is_mstatus(exu_io_prev_bits_id2ex_csr_hit_is_mstatus),
    .io_prev_bits_id2ex_csr_hit_is_mie(exu_io_prev_bits_id2ex_csr_hit_is_mie),
    .io_prev_bits_id2ex_csr_hit_is_mcause(exu_io_prev_bits_id2ex_csr_hit_is_mcause),
    .io_prev_bits_id2ex_csr_hit_is_mip(exu_io_prev_bits_id2ex_csr_hit_is_mip),
    .io_prev_bits_id2ex_csr_hit_is_mtime(exu_io_prev_bits_id2ex_csr_hit_is_mtime),
    .io_prev_bits_id2ex_csr_hit_is_mcycle(exu_io_prev_bits_id2ex_csr_hit_is_mcycle),
    .io_prev_bits_id2ex_csr_hit_is_mhartid(exu_io_prev_bits_id2ex_csr_hit_is_mhartid),
    .io_prev_bits_id2ex_mdu_op_mul_signed(exu_io_prev_bits_id2ex_mdu_op_mul_signed),
    .io_prev_bits_id2ex_mdu_op_is_mu(exu_io_prev_bits_id2ex_mdu_op_is_mu),
    .io_prev_bits_id2ex_mdu_op_mul_32(exu_io_prev_bits_id2ex_mdu_op_mul_32),
    .io_prev_bits_id2ex_mdu_op_div_signed(exu_io_prev_bits_id2ex_mdu_op_div_signed),
    .io_prev_bits_id2ex_mdu_op_is_div(exu_io_prev_bits_id2ex_mdu_op_is_div),
    .io_prev_bits_id2ex_mdu_op_is_du(exu_io_prev_bits_id2ex_mdu_op_is_du),
    .io_prev_bits_id2ex_zimm(exu_io_prev_bits_id2ex_zimm),
    .io_prev_bits_id2ex_intr(exu_io_prev_bits_id2ex_intr),
    .io_prev_bits_id2ex_exec(exu_io_prev_bits_id2ex_exec),
    .io_prev_bits_id2ex_mret(exu_io_prev_bits_id2ex_mret),
    .io_prev_bits_id2ex_exce_code(exu_io_prev_bits_id2ex_exce_code),
    .io_prev_bits_id2ex_pc(exu_io_prev_bits_id2ex_pc),
    .io_prev_bits_id2ex_is_iem(exu_io_prev_bits_id2ex_is_iem),
    .io_prev_bits_id2mem_fencei(exu_io_prev_bits_id2mem_fencei),
    .io_prev_bits_id2mem_size_byte(exu_io_prev_bits_id2mem_size_byte),
    .io_prev_bits_id2mem_size_hword(exu_io_prev_bits_id2mem_size_hword),
    .io_prev_bits_id2mem_size_word(exu_io_prev_bits_id2mem_size_word),
    .io_prev_bits_id2mem_size_dword(exu_io_prev_bits_id2mem_size_dword),
    .io_prev_bits_id2mem_sext_flag(exu_io_prev_bits_id2mem_sext_flag),
    .io_prev_bits_id2mem_memory_rd_en(exu_io_prev_bits_id2mem_memory_rd_en),
    .io_prev_bits_id2mem_memory_we_en(exu_io_prev_bits_id2mem_memory_we_en),
    .io_prev_bits_id2wb_intr_exce_ret(exu_io_prev_bits_id2wb_intr_exce_ret),
    .io_prev_bits_id2wb_fencei(exu_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_wb_sel(exu_io_prev_bits_id2wb_wb_sel),
    .io_prev_bits_id2wb_regfile_we_en(exu_io_prev_bits_id2wb_regfile_we_en),
    .io_prev_bits_id2wb_regfile_we_addr(exu_io_prev_bits_id2wb_regfile_we_addr),
    .io_next_ready(exu_io_next_ready),
    .io_next_valid(exu_io_next_valid),
    .io_next_bits_id2mem_fencei(exu_io_next_bits_id2mem_fencei),
    .io_next_bits_id2mem_size_byte(exu_io_next_bits_id2mem_size_byte),
    .io_next_bits_id2mem_size_hword(exu_io_next_bits_id2mem_size_hword),
    .io_next_bits_id2mem_size_word(exu_io_next_bits_id2mem_size_word),
    .io_next_bits_id2mem_size_dword(exu_io_next_bits_id2mem_size_dword),
    .io_next_bits_id2mem_sext_flag(exu_io_next_bits_id2mem_sext_flag),
    .io_next_bits_id2mem_memory_rd_en(exu_io_next_bits_id2mem_memory_rd_en),
    .io_next_bits_id2mem_memory_we_en(exu_io_next_bits_id2mem_memory_we_en),
    .io_next_bits_id2wb_intr_exce_ret(exu_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(exu_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(exu_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(exu_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(exu_io_next_bits_id2wb_regfile_we_addr),
    .io_next_bits_ex2mem_addr(exu_io_next_bits_ex2mem_addr),
    .io_next_bits_ex2mem_we_data(exu_io_next_bits_ex2mem_we_data),
    .io_next_bits_ex2mem_we_mask(exu_io_next_bits_ex2mem_we_mask),
    .io_next_bits_ex2wb_result_data(exu_io_next_bits_ex2wb_result_data),
    .io_csr2ctrl_out_mepc(exu_io_csr2ctrl_out_mepc),
    .io_csr2ctrl_out_mtvec(exu_io_csr2ctrl_out_mtvec),
    .io_csr2ctrl_out_mie(exu_io_csr2ctrl_out_mie),
    .io_csr2ctrl_out_mtie(exu_io_csr2ctrl_out_mtie),
    .io_csr2ctrl_out_msie(exu_io_csr2ctrl_out_msie),
    .io_csr2ctrl_out_meie(exu_io_csr2ctrl_out_meie),
    .io_csr2ctrl_out_mtip(exu_io_csr2ctrl_out_mtip),
    .io_csr2ctrl_out_msip(exu_io_csr2ctrl_out_msip),
    .io_csr2ctrl_out_meip(exu_io_csr2ctrl_out_meip),
    .io_sb_clint_msip(exu_io_sb_clint_msip),
    .io_sb_clint_mtip(exu_io_sb_clint_mtip),
    .io_sb_clint_mtime(exu_io_sb_clint_mtime),
    .io_sb_meip(exu_io_sb_meip)
  );
  ysyx_040978_MEMReg EX2MEMReg ( // @[MEMU.scala 84:27]
    .clock(EX2MEMReg_clock),
    .reset(EX2MEMReg_reset),
    .io_prev_ready(EX2MEMReg_io_prev_ready),
    .io_prev_valid(EX2MEMReg_io_prev_valid),
    .io_prev_bits_id2mem_fencei(EX2MEMReg_io_prev_bits_id2mem_fencei),
    .io_prev_bits_id2mem_size_byte(EX2MEMReg_io_prev_bits_id2mem_size_byte),
    .io_prev_bits_id2mem_size_hword(EX2MEMReg_io_prev_bits_id2mem_size_hword),
    .io_prev_bits_id2mem_size_word(EX2MEMReg_io_prev_bits_id2mem_size_word),
    .io_prev_bits_id2mem_size_dword(EX2MEMReg_io_prev_bits_id2mem_size_dword),
    .io_prev_bits_id2mem_sext_flag(EX2MEMReg_io_prev_bits_id2mem_sext_flag),
    .io_prev_bits_id2mem_memory_rd_en(EX2MEMReg_io_prev_bits_id2mem_memory_rd_en),
    .io_prev_bits_id2mem_memory_we_en(EX2MEMReg_io_prev_bits_id2mem_memory_we_en),
    .io_prev_bits_id2wb_intr_exce_ret(EX2MEMReg_io_prev_bits_id2wb_intr_exce_ret),
    .io_prev_bits_id2wb_fencei(EX2MEMReg_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_wb_sel(EX2MEMReg_io_prev_bits_id2wb_wb_sel),
    .io_prev_bits_id2wb_regfile_we_en(EX2MEMReg_io_prev_bits_id2wb_regfile_we_en),
    .io_prev_bits_id2wb_regfile_we_addr(EX2MEMReg_io_prev_bits_id2wb_regfile_we_addr),
    .io_prev_bits_ex2mem_addr(EX2MEMReg_io_prev_bits_ex2mem_addr),
    .io_prev_bits_ex2mem_we_data(EX2MEMReg_io_prev_bits_ex2mem_we_data),
    .io_prev_bits_ex2mem_we_mask(EX2MEMReg_io_prev_bits_ex2mem_we_mask),
    .io_prev_bits_ex2wb_result_data(EX2MEMReg_io_prev_bits_ex2wb_result_data),
    .io_next_ready(EX2MEMReg_io_next_ready),
    .io_next_valid(EX2MEMReg_io_next_valid),
    .io_next_bits_id2mem_fencei(EX2MEMReg_io_next_bits_id2mem_fencei),
    .io_next_bits_id2mem_size_byte(EX2MEMReg_io_next_bits_id2mem_size_byte),
    .io_next_bits_id2mem_size_hword(EX2MEMReg_io_next_bits_id2mem_size_hword),
    .io_next_bits_id2mem_size_word(EX2MEMReg_io_next_bits_id2mem_size_word),
    .io_next_bits_id2mem_size_dword(EX2MEMReg_io_next_bits_id2mem_size_dword),
    .io_next_bits_id2mem_sext_flag(EX2MEMReg_io_next_bits_id2mem_sext_flag),
    .io_next_bits_id2mem_memory_rd_en(EX2MEMReg_io_next_bits_id2mem_memory_rd_en),
    .io_next_bits_id2mem_memory_we_en(EX2MEMReg_io_next_bits_id2mem_memory_we_en),
    .io_next_bits_id2wb_intr_exce_ret(EX2MEMReg_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(EX2MEMReg_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(EX2MEMReg_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(EX2MEMReg_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(EX2MEMReg_io_next_bits_id2wb_regfile_we_addr),
    .io_next_bits_ex2mem_addr(EX2MEMReg_io_next_bits_ex2mem_addr),
    .io_next_bits_ex2mem_we_data(EX2MEMReg_io_next_bits_ex2mem_we_data),
    .io_next_bits_ex2mem_we_mask(EX2MEMReg_io_next_bits_ex2mem_we_mask),
    .io_next_bits_ex2wb_result_data(EX2MEMReg_io_next_bits_ex2wb_result_data)
  );
  ysyx_040978_MEMU memu ( // @[MEMU.scala 87:22]
    .clock(memu_clock),
    .reset(memu_reset),
    .io_prev_ready(memu_io_prev_ready),
    .io_prev_valid(memu_io_prev_valid),
    .io_prev_bits_id2mem_fencei(memu_io_prev_bits_id2mem_fencei),
    .io_prev_bits_id2mem_size_byte(memu_io_prev_bits_id2mem_size_byte),
    .io_prev_bits_id2mem_size_hword(memu_io_prev_bits_id2mem_size_hword),
    .io_prev_bits_id2mem_size_word(memu_io_prev_bits_id2mem_size_word),
    .io_prev_bits_id2mem_size_dword(memu_io_prev_bits_id2mem_size_dword),
    .io_prev_bits_id2mem_sext_flag(memu_io_prev_bits_id2mem_sext_flag),
    .io_prev_bits_id2mem_memory_rd_en(memu_io_prev_bits_id2mem_memory_rd_en),
    .io_prev_bits_id2mem_memory_we_en(memu_io_prev_bits_id2mem_memory_we_en),
    .io_prev_bits_id2wb_intr_exce_ret(memu_io_prev_bits_id2wb_intr_exce_ret),
    .io_prev_bits_id2wb_fencei(memu_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_wb_sel(memu_io_prev_bits_id2wb_wb_sel),
    .io_prev_bits_id2wb_regfile_we_en(memu_io_prev_bits_id2wb_regfile_we_en),
    .io_prev_bits_id2wb_regfile_we_addr(memu_io_prev_bits_id2wb_regfile_we_addr),
    .io_prev_bits_ex2mem_addr(memu_io_prev_bits_ex2mem_addr),
    .io_prev_bits_ex2mem_we_data(memu_io_prev_bits_ex2mem_we_data),
    .io_prev_bits_ex2mem_we_mask(memu_io_prev_bits_ex2mem_we_mask),
    .io_prev_bits_ex2wb_result_data(memu_io_prev_bits_ex2wb_result_data),
    .io_next_valid(memu_io_next_valid),
    .io_next_bits_id2wb_intr_exce_ret(memu_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(memu_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(memu_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(memu_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(memu_io_next_bits_id2wb_regfile_we_addr),
    .io_next_bits_ex2wb_result_data(memu_io_next_bits_ex2wb_result_data),
    .io_next_bits_mem2wb_memory_data(memu_io_next_bits_mem2wb_memory_data),
    .io_maxi_ar_ready(memu_io_maxi_ar_ready),
    .io_maxi_ar_valid(memu_io_maxi_ar_valid),
    .io_maxi_ar_bits_addr(memu_io_maxi_ar_bits_addr),
    .io_maxi_ar_bits_len(memu_io_maxi_ar_bits_len),
    .io_maxi_ar_bits_size(memu_io_maxi_ar_bits_size),
    .io_maxi_r_valid(memu_io_maxi_r_valid),
    .io_maxi_r_bits_data(memu_io_maxi_r_bits_data),
    .io_maxi_r_bits_last(memu_io_maxi_r_bits_last),
    .io_maxi_aw_ready(memu_io_maxi_aw_ready),
    .io_maxi_aw_valid(memu_io_maxi_aw_valid),
    .io_maxi_aw_bits_addr(memu_io_maxi_aw_bits_addr),
    .io_maxi_aw_bits_len(memu_io_maxi_aw_bits_len),
    .io_maxi_aw_bits_size(memu_io_maxi_aw_bits_size),
    .io_maxi_w_ready(memu_io_maxi_w_ready),
    .io_maxi_w_valid(memu_io_maxi_w_valid),
    .io_maxi_w_bits_data(memu_io_maxi_w_bits_data),
    .io_maxi_w_bits_strb(memu_io_maxi_w_bits_strb),
    .io_maxi_w_bits_last(memu_io_maxi_w_bits_last),
    .io_maxi_b_valid(memu_io_maxi_b_valid),
    .io_mmio_ar_ready(memu_io_mmio_ar_ready),
    .io_mmio_ar_valid(memu_io_mmio_ar_valid),
    .io_mmio_ar_bits_addr(memu_io_mmio_ar_bits_addr),
    .io_mmio_ar_bits_size(memu_io_mmio_ar_bits_size),
    .io_mmio_r_valid(memu_io_mmio_r_valid),
    .io_mmio_r_bits_data(memu_io_mmio_r_bits_data),
    .io_mmio_r_bits_last(memu_io_mmio_r_bits_last),
    .io_mmio_aw_ready(memu_io_mmio_aw_ready),
    .io_mmio_aw_valid(memu_io_mmio_aw_valid),
    .io_mmio_aw_bits_addr(memu_io_mmio_aw_bits_addr),
    .io_mmio_aw_bits_size(memu_io_mmio_aw_bits_size),
    .io_mmio_w_ready(memu_io_mmio_w_ready),
    .io_mmio_w_valid(memu_io_mmio_w_valid),
    .io_mmio_w_bits_data(memu_io_mmio_w_bits_data),
    .io_mmio_w_bits_strb(memu_io_mmio_w_bits_strb),
    .io_mmio_w_bits_last(memu_io_mmio_w_bits_last),
    .io_mmio_b_valid(memu_io_mmio_b_valid),
    .io_sram4_addr(memu_io_sram4_addr),
    .io_sram4_wen(memu_io_sram4_wen),
    .io_sram4_wmask(memu_io_sram4_wmask),
    .io_sram4_wdata(memu_io_sram4_wdata),
    .io_sram4_rdata(memu_io_sram4_rdata),
    .io_sram5_addr(memu_io_sram5_addr),
    .io_sram5_wen(memu_io_sram5_wen),
    .io_sram5_wmask(memu_io_sram5_wmask),
    .io_sram5_wdata(memu_io_sram5_wdata),
    .io_sram5_rdata(memu_io_sram5_rdata),
    .io_sram6_addr(memu_io_sram6_addr),
    .io_sram6_wen(memu_io_sram6_wen),
    .io_sram6_wmask(memu_io_sram6_wmask),
    .io_sram6_wdata(memu_io_sram6_wdata),
    .io_sram6_rdata(memu_io_sram6_rdata),
    .io_sram7_addr(memu_io_sram7_addr),
    .io_sram7_wen(memu_io_sram7_wen),
    .io_sram7_wmask(memu_io_sram7_wmask),
    .io_sram7_wdata(memu_io_sram7_wdata),
    .io_sram7_rdata(memu_io_sram7_rdata),
    .clint_we(memu_clint_we),
    ._T_24(memu__T_24),
    .clint_rdata(memu_clint_rdata),
    .clint_wdata(memu_clint_wdata)
  );
  ysyx_040978_WBReg MEM2WBReg ( // @[WBU.scala 77:27]
    .clock(MEM2WBReg_clock),
    .reset(MEM2WBReg_reset),
    .io_prev_valid(MEM2WBReg_io_prev_valid),
    .io_prev_bits_id2wb_intr_exce_ret(MEM2WBReg_io_prev_bits_id2wb_intr_exce_ret),
    .io_prev_bits_id2wb_fencei(MEM2WBReg_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_wb_sel(MEM2WBReg_io_prev_bits_id2wb_wb_sel),
    .io_prev_bits_id2wb_regfile_we_en(MEM2WBReg_io_prev_bits_id2wb_regfile_we_en),
    .io_prev_bits_id2wb_regfile_we_addr(MEM2WBReg_io_prev_bits_id2wb_regfile_we_addr),
    .io_prev_bits_ex2wb_result_data(MEM2WBReg_io_prev_bits_ex2wb_result_data),
    .io_prev_bits_mem2wb_memory_data(MEM2WBReg_io_prev_bits_mem2wb_memory_data),
    .io_next_valid(MEM2WBReg_io_next_valid),
    .io_next_bits_id2wb_intr_exce_ret(MEM2WBReg_io_next_bits_id2wb_intr_exce_ret),
    .io_next_bits_id2wb_fencei(MEM2WBReg_io_next_bits_id2wb_fencei),
    .io_next_bits_id2wb_wb_sel(MEM2WBReg_io_next_bits_id2wb_wb_sel),
    .io_next_bits_id2wb_regfile_we_en(MEM2WBReg_io_next_bits_id2wb_regfile_we_en),
    .io_next_bits_id2wb_regfile_we_addr(MEM2WBReg_io_next_bits_id2wb_regfile_we_addr),
    .io_next_bits_ex2wb_result_data(MEM2WBReg_io_next_bits_ex2wb_result_data),
    .io_next_bits_mem2wb_memory_data(MEM2WBReg_io_next_bits_mem2wb_memory_data)
  );
  ysyx_040978_WBU wbu ( // @[WBU.scala 80:21]
    .io__prev_valid(wbu_io__prev_valid),
    .io__prev_bits_id2wb_intr_exce_ret(wbu_io__prev_bits_id2wb_intr_exce_ret),
    .io__prev_bits_id2wb_fencei(wbu_io__prev_bits_id2wb_fencei),
    .io__prev_bits_id2wb_wb_sel(wbu_io__prev_bits_id2wb_wb_sel),
    .io__prev_bits_id2wb_regfile_we_en(wbu_io__prev_bits_id2wb_regfile_we_en),
    .io__prev_bits_id2wb_regfile_we_addr(wbu_io__prev_bits_id2wb_regfile_we_addr),
    .io__prev_bits_ex2wb_result_data(wbu_io__prev_bits_ex2wb_result_data),
    .io__prev_bits_mem2wb_memory_data(wbu_io__prev_bits_mem2wb_memory_data),
    .io__regfile_en(wbu_io__regfile_en),
    .io__regfile_addr(wbu_io__regfile_addr),
    .io__regfile_data(wbu_io__regfile_data),
    .io_prev_bits_id2wb_fencei(wbu_io_prev_bits_id2wb_fencei),
    .io_prev_bits_id2wb_intr_exce_ret(wbu_io_prev_bits_id2wb_intr_exce_ret)
  );
  ysyx_040978_FWU fwu ( // @[FWU.scala 102:21]
    .io_idu_fw_src1_data(fwu_io_idu_fw_src1_data),
    .io_idu_fw_src2_data(fwu_io_idu_fw_src2_data),
    .io_idu_fw_ready(fwu_io_idu_fw_ready),
    .io_idu_optype_Itype(fwu_io_idu_optype_Itype),
    .io_idu_src1_addr(fwu_io_idu_src1_addr),
    .io_idu_src2_addr(fwu_io_idu_src2_addr),
    .io_idu_src1_data(fwu_io_idu_src1_data),
    .io_idu_src2_data(fwu_io_idu_src2_data),
    .io_exu_is_load(fwu_io_exu_is_load),
    .io_exu_dst_addr(fwu_io_exu_dst_addr),
    .io_exu_dst_data(fwu_io_exu_dst_data),
    .io_memu_is_load_1(fwu_io_memu_is_load_1),
    .io_memu_dst_addr_1(fwu_io_memu_dst_addr_1),
    .io_memu_dst_data_1(fwu_io_memu_dst_data_1),
    .io_memu_dst_addr_2(fwu_io_memu_dst_addr_2),
    .io_wbu_dst_addr(fwu_io_wbu_dst_addr),
    .io_wbu_dst_data(fwu_io_wbu_dst_data)
  );
  ysyx_040978_BRU bru ( // @[BRU.scala 56:21]
    .clock(bru_clock),
    .reset(bru_reset),
    .io_idu_brh(bru_io_idu_brh),
    .io_idu_jal(bru_io_idu_jal),
    .io_idu_jalr(bru_io_idu_jalr),
    .io_idu_pc(bru_io_idu_pc),
    .io_idu_src1(bru_io_idu_src1),
    .io_idu_src2(bru_io_idu_src2),
    .io_idu_imm(bru_io_idu_imm),
    .io_ifu_jump(bru_io_ifu_jump),
    .io_ifu_npc(bru_io_ifu_npc),
    .io_ifu_jump0(bru_io_ifu_jump0)
  );
  ysyx_040978_RegFile regfile ( // @[Top.scala 53:31]
    .clock(regfile_clock),
    .reset(regfile_reset),
    .io_wbu_en(regfile_io_wbu_en),
    .io_wbu_addr(regfile_io_wbu_addr),
    .io_wbu_data(regfile_io_wbu_data),
    .io_idu_addr1(regfile_io_idu_addr1),
    .io_idu_data1(regfile_io_idu_data1),
    .io_idu_addr2(regfile_io_idu_addr2),
    .io_idu_data2(regfile_io_idu_data2)
  );
  assign io_maxi4_ar_valid = icon_io_maxi_ar_valid; // @[AXI.scala 286:27]
  assign io_maxi4_ar_bits_addr = icon_io_maxi_ar_bits_addr; // @[AXI.scala 286:27]
  assign io_maxi4_ar_bits_burst = 2'h1; // @[AXI.scala 286:27]
  assign io_maxi4_ar_bits_id = icon_io_maxi_ar_bits_id; // @[AXI.scala 286:27]
  assign io_maxi4_ar_bits_len = icon_io_maxi_ar_bits_len; // @[AXI.scala 286:27]
  assign io_maxi4_ar_bits_size = icon_io_maxi_ar_bits_size; // @[AXI.scala 286:27]
  assign io_maxi4_r_ready = 1'h1; // @[AXI.scala 286:27]
  assign io_maxi4_aw_valid = icon_io_maxi_aw_valid; // @[AXI.scala 286:27]
  assign io_maxi4_aw_bits_addr = icon_io_maxi_aw_bits_addr; // @[AXI.scala 286:27]
  assign io_maxi4_aw_bits_burst = 2'h1; // @[AXI.scala 286:27]
  assign io_maxi4_aw_bits_id = icon_io_maxi_aw_bits_id; // @[AXI.scala 286:27]
  assign io_maxi4_aw_bits_len = icon_io_maxi_aw_bits_len; // @[AXI.scala 286:27]
  assign io_maxi4_aw_bits_size = icon_io_maxi_aw_bits_size; // @[AXI.scala 286:27]
  assign io_maxi4_w_valid = icon_io_maxi_w_valid; // @[AXI.scala 286:27]
  assign io_maxi4_w_bits_data = icon_io_maxi_w_bits_data; // @[AXI.scala 286:27]
  assign io_maxi4_w_bits_strb = icon_io_maxi_w_bits_strb; // @[AXI.scala 286:27]
  assign io_maxi4_w_bits_last = icon_io_maxi_w_bits_last; // @[AXI.scala 286:27]
  assign io_maxi4_b_ready = 1'h1; // @[AXI.scala 286:27]
  assign io_sram0_addr = sram_init_reg ? sram_init_cnt : ifu_io_sram0_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 58:17]
  assign io_sram0_wen = sram_init_reg ? 1'h0 : ifu_io_sram0_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 58:17]
  assign io_sram0_wmask = sram_init_reg ? 128'h0 : ifu_io_sram0_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 58:17]
  assign io_sram0_wdata = sram_init_reg ? 128'h0 : ifu_io_sram0_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 58:17]
  assign io_sram1_addr = sram_init_reg ? sram_init_cnt : ifu_io_sram1_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 59:17]
  assign io_sram1_wen = sram_init_reg ? 1'h0 : ifu_io_sram1_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 59:17]
  assign io_sram1_wmask = sram_init_reg ? 128'h0 : ifu_io_sram1_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 59:17]
  assign io_sram1_wdata = sram_init_reg ? 128'h0 : ifu_io_sram1_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 59:17]
  assign io_sram2_addr = sram_init_reg ? sram_init_cnt : ifu_io_sram2_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 60:17]
  assign io_sram2_wen = sram_init_reg ? 1'h0 : ifu_io_sram2_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 60:17]
  assign io_sram2_wmask = sram_init_reg ? 128'h0 : ifu_io_sram2_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 60:17]
  assign io_sram2_wdata = sram_init_reg ? 128'h0 : ifu_io_sram2_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 60:17]
  assign io_sram3_addr = sram_init_reg ? sram_init_cnt : ifu_io_sram3_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 61:17]
  assign io_sram3_wen = sram_init_reg ? 1'h0 : ifu_io_sram3_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 61:17]
  assign io_sram3_wmask = sram_init_reg ? 128'h0 : ifu_io_sram3_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 61:17]
  assign io_sram3_wdata = sram_init_reg ? 128'h0 : ifu_io_sram3_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 61:17]
  assign io_sram4_addr = sram_init_reg ? sram_init_cnt : memu_io_sram4_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 62:17]
  assign io_sram4_wen = sram_init_reg ? 1'h0 : memu_io_sram4_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 62:17]
  assign io_sram4_wmask = sram_init_reg ? 128'h0 : memu_io_sram4_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 62:17]
  assign io_sram4_wdata = sram_init_reg ? 128'h0 : memu_io_sram4_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 62:17]
  assign io_sram5_addr = sram_init_reg ? sram_init_cnt : memu_io_sram5_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 63:17]
  assign io_sram5_wen = sram_init_reg ? 1'h0 : memu_io_sram5_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 63:17]
  assign io_sram5_wmask = sram_init_reg ? 128'h0 : memu_io_sram5_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 63:17]
  assign io_sram5_wdata = sram_init_reg ? 128'h0 : memu_io_sram5_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 63:17]
  assign io_sram6_addr = sram_init_reg ? sram_init_cnt : memu_io_sram6_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 64:17]
  assign io_sram6_wen = sram_init_reg ? 1'h0 : memu_io_sram6_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 64:17]
  assign io_sram6_wmask = sram_init_reg ? 128'h0 : memu_io_sram6_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 64:17]
  assign io_sram6_wdata = sram_init_reg ? 128'h0 : memu_io_sram6_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 64:17]
  assign io_sram7_addr = sram_init_reg ? sram_init_cnt : memu_io_sram7_addr; // @[Top.scala 66:22 CacheBase.scala 73:14 Top.scala 65:17]
  assign io_sram7_wen = sram_init_reg ? 1'h0 : memu_io_sram7_wen; // @[Top.scala 66:22 CacheBase.scala 72:13 Top.scala 65:17]
  assign io_sram7_wmask = sram_init_reg ? 128'h0 : memu_io_sram7_wmask; // @[Top.scala 66:22 CacheBase.scala 75:15 Top.scala 65:17]
  assign io_sram7_wdata = sram_init_reg ? 128'h0 : memu_io_sram7_wdata; // @[Top.scala 66:22 CacheBase.scala 74:15 Top.scala 65:17]
  assign clint_we = memu_clint_we;
  assign _T_24 = memu__T_24;
  assign clint_wdata = memu_clint_wdata;
  assign icon_clock = clock;
  assign icon_reset = reset;
  assign icon_io_maxi_ar_ready = io_maxi4_ar_ready; // @[AXI.scala 286:27]
  assign icon_io_maxi_r_valid = io_maxi4_r_valid; // @[AXI.scala 286:27]
  assign icon_io_maxi_r_bits_data = io_maxi4_r_bits_data; // @[AXI.scala 286:27]
  assign icon_io_maxi_r_bits_id = io_maxi4_r_bits_id; // @[AXI.scala 286:27]
  assign icon_io_maxi_r_bits_last = io_maxi4_r_bits_last; // @[AXI.scala 286:27]
  assign icon_io_maxi_aw_ready = io_maxi4_aw_ready; // @[AXI.scala 286:27]
  assign icon_io_maxi_w_ready = io_maxi4_w_ready; // @[AXI.scala 286:27]
  assign icon_io_maxi_b_valid = io_maxi4_b_valid; // @[AXI.scala 286:27]
  assign icon_io_maxi_b_bits_id = io_maxi4_b_bits_id; // @[AXI.scala 286:27]
  assign icon_io_ifu_ar_valid = ifu_io_maxi_ar_valid; // @[Top.scala 38:27 IFU.scala 110:10]
  assign icon_io_ifu_ar_bits_addr = ifu_io_maxi_ar_bits_addr; // @[Top.scala 38:27 IFU.scala 110:10]
  assign icon_io_ifu_ar_bits_len = ifu_io_maxi_ar_bits_len; // @[Top.scala 38:27 IFU.scala 110:10]
  assign icon_io_ifu_ar_bits_size = ifu_io_maxi_ar_bits_size; // @[Top.scala 38:27 IFU.scala 110:10]
  assign icon_io_memu_ar_valid = memu_io_maxi_ar_valid; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_ar_bits_addr = memu_io_maxi_ar_bits_addr; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_ar_bits_len = memu_io_maxi_ar_bits_len; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_ar_bits_size = memu_io_maxi_ar_bits_size; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_aw_valid = memu_io_maxi_aw_valid; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_aw_bits_addr = memu_io_maxi_aw_bits_addr; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_aw_bits_len = memu_io_maxi_aw_bits_len; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_aw_bits_size = memu_io_maxi_aw_bits_size; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_w_valid = memu_io_maxi_w_valid; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_w_bits_data = memu_io_maxi_w_bits_data; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_w_bits_strb = memu_io_maxi_w_bits_strb; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_memu_w_bits_last = memu_io_maxi_w_bits_last; // @[Top.scala 39:28 MEMU.scala 89:18]
  assign icon_io_devu_ar_valid = memu_io_mmio_ar_valid; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_ar_bits_addr = memu_io_mmio_ar_bits_addr; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_ar_bits_size = memu_io_mmio_ar_bits_size; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_aw_valid = memu_io_mmio_aw_valid; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_aw_bits_addr = memu_io_mmio_aw_bits_addr; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_aw_bits_size = memu_io_mmio_aw_bits_size; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_w_valid = memu_io_mmio_w_valid; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_w_bits_data = memu_io_mmio_w_bits_data; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_w_bits_strb = memu_io_mmio_w_bits_strb; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign icon_io_devu_w_bits_last = memu_io_mmio_w_bits_last; // @[Top.scala 40:29 MEMU.scala 90:18]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_jump0 = bru_io_ifu_jump0; // @[Top.scala 23:29 BRU.scala 57:16]
  assign pc_io_jump = bru_io_ifu_jump; // @[Top.scala 23:29 BRU.scala 57:16]
  assign pc_io_npc = bru_io_ifu_npc; // @[Top.scala 23:29 BRU.scala 57:16]
  assign pc_io_sys_ready = ~sram_init_reg; // @[Top.scala 45:81]
  assign pc_io_next_ready = ifu_io_prev_ready; // @[IFU.scala 103:17]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_cache_reset = bru_io_ifu_jump0; // @[Top.scala 23:29 BRU.scala 57:16]
  assign ifu_io_prev_valid = pc_io_next_valid; // @[IFU.scala 103:17]
  assign ifu_io_prev_bits_pc2if_pc = pc_io_next_bits_pc2if_pc; // @[IFU.scala 103:17]
  assign ifu_io_maxi_ar_ready = icon_io_ifu_ar_ready; // @[Top.scala 38:27 AXI.scala 287:27]
  assign ifu_io_maxi_r_valid = icon_io_ifu_r_valid; // @[Top.scala 38:27 AXI.scala 287:27]
  assign ifu_io_maxi_r_bits_data = icon_io_ifu_r_bits_data; // @[Top.scala 38:27 AXI.scala 287:27]
  assign ifu_io_maxi_r_bits_last = icon_io_ifu_r_bits_last; // @[Top.scala 38:27 AXI.scala 287:27]
  assign ifu_io_next_ready = IF2IDReg_io_prev_ready; // @[Top.scala 25:29 IDU.scala 288:22]
  assign ifu_io_sram0_rdata = io_sram0_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 58:17]
  assign ifu_io_sram1_rdata = io_sram1_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 59:17]
  assign ifu_io_sram2_rdata = io_sram2_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 60:17]
  assign ifu_io_sram3_rdata = io_sram3_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 61:17]
  assign ifu_fenceiing = idu_fenceiing_0;
  assign IF2IDReg_clock = clock;
  assign IF2IDReg_reset = BRIFBdl_jump | reset; // @[IDU.scala 287:17 IDU.scala 287:34]
  assign IF2IDReg_io_prev_valid = ifu_io_next_valid; // @[Top.scala 25:29 IFU.scala 109:10]
  assign IF2IDReg_io_prev_bits_if2id_inst = ifu_io_next_bits_if2id_inst; // @[Top.scala 25:29 IFU.scala 109:10]
  assign IF2IDReg_io_prev_bits_if2id_pc = ifu_io_next_bits_if2id_pc; // @[Top.scala 25:29 IFU.scala 109:10]
  assign IF2IDReg_io_next_ready = idu_io_prev_ready; // @[IDU.scala 294:17]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_regfile_data1 = regfile_io_idu_data1; // @[Top.scala 35:34 Top.scala 55:18]
  assign idu_io_regfile_data2 = regfile_io_idu_data2; // @[Top.scala 35:34 Top.scala 55:18]
  assign idu_io_fwu_fw_src1_data = fwu_io_idu_fw_src1_data; // @[Top.scala 29:29 FWU.scala 103:16]
  assign idu_io_fwu_fw_src2_data = fwu_io_idu_fw_src2_data; // @[Top.scala 29:29 FWU.scala 103:16]
  assign idu_io_csr_out_mepc = exu_io_csr2ctrl_out_mepc; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_mtvec = exu_io_csr2ctrl_out_mtvec; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_mie = exu_io_csr2ctrl_out_mie; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_mtie = exu_io_csr2ctrl_out_mtie; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_msie = exu_io_csr2ctrl_out_msie; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_meie = exu_io_csr2ctrl_out_meie; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_mtip = exu_io_csr2ctrl_out_mtip; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_msip = exu_io_csr2ctrl_out_msip; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_csr_out_meip = exu_io_csr2ctrl_out_meip; // @[Top.scala 33:32 EXU.scala 160:21]
  assign idu_io_prev_valid = IF2IDReg_io_next_valid; // @[IDU.scala 294:17]
  assign idu_io_prev_bits_if2id_inst = IF2IDReg_io_next_bits_if2id_inst; // @[IDU.scala 294:17]
  assign idu_io_prev_bits_if2id_pc = IF2IDReg_io_next_bits_if2id_pc; // @[IDU.scala 294:17]
  assign idu_io_next_ready = IDUOut_ready & IDFWBdl_fw_ready; // @[IDU.scala 298:37]
  assign idu_wb_fencei_0 = wbu_io_prev_bits_id2wb_fencei;
  assign idu_wb_intr_exce_ret_0 = wbu_io_prev_bits_id2wb_intr_exce_ret;
  assign ID2EXReg_clock = clock;
  assign ID2EXReg_reset = reset;
  assign ID2EXReg_io_prev_valid = idu_io_next_valid & IDFWBdl_fw_ready; // @[IDU.scala 299:37]
  assign ID2EXReg_io_prev_bits_id2ex_alu_src1 = idu_io_next_bits_id2ex_alu_src1; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_alu_src2 = idu_io_next_bits_id2ex_alu_src2; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_salu_src1 = idu_io_next_bits_id2ex_salu_src1; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_salu_src2 = idu_io_next_bits_id2ex_salu_src2; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_src1 = idu_io_next_bits_id2ex_src1; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_src2 = idu_io_next_bits_id2ex_src2; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_src3 = idu_io_next_bits_id2ex_src3; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_auipc = idu_io_next_bits_id2ex_operator_auipc; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_lui = idu_io_next_bits_id2ex_operator_lui; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_jal = idu_io_next_bits_id2ex_operator_jal; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_jalr = idu_io_next_bits_id2ex_operator_jalr; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sb = idu_io_next_bits_id2ex_operator_sb; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sh = idu_io_next_bits_id2ex_operator_sh; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sw = idu_io_next_bits_id2ex_operator_sw; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sd = idu_io_next_bits_id2ex_operator_sd; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_add = idu_io_next_bits_id2ex_operator_add; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sub = idu_io_next_bits_id2ex_operator_sub; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sll = idu_io_next_bits_id2ex_operator_sll; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_slt = idu_io_next_bits_id2ex_operator_slt; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sltu = idu_io_next_bits_id2ex_operator_sltu; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_xor = idu_io_next_bits_id2ex_operator_xor; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_srl = idu_io_next_bits_id2ex_operator_srl; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_sra = idu_io_next_bits_id2ex_operator_sra; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_or = idu_io_next_bits_id2ex_operator_or; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_and = idu_io_next_bits_id2ex_operator_and; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_is_csr = idu_io_next_bits_id2ex_operator_csr_is_csr; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrw = idu_io_next_bits_id2ex_operator_csr_csrrw; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrs = idu_io_next_bits_id2ex_operator_csr_csrrs; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrc = idu_io_next_bits_id2ex_operator_csr_csrrc; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrwi = idu_io_next_bits_id2ex_operator_csr_csrrwi; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrsi = idu_io_next_bits_id2ex_operator_csr_csrrsi; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_operator_csr_csrrci = idu_io_next_bits_id2ex_operator_csr_csrrci; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_srcsize_byte = idu_io_next_bits_id2ex_srcsize_byte; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_srcsize_hword = idu_io_next_bits_id2ex_srcsize_hword; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_srcsize_word = idu_io_next_bits_id2ex_srcsize_word; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_srcsize_dword = idu_io_next_bits_id2ex_srcsize_dword; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_is_load = idu_io_next_bits_id2ex_is_load; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_is_save = idu_io_next_bits_id2ex_is_save; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_div_inf = idu_io_next_bits_id2ex_div_inf; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_we = idu_io_next_bits_id2ex_csr_we; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mepc = idu_io_next_bits_id2ex_csr_hit_is_mepc; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtvec = idu_io_next_bits_id2ex_csr_hit_is_mtvec; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mstatus = idu_io_next_bits_id2ex_csr_hit_is_mstatus; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mie = idu_io_next_bits_id2ex_csr_hit_is_mie; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcause = idu_io_next_bits_id2ex_csr_hit_is_mcause; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mip = idu_io_next_bits_id2ex_csr_hit_is_mip; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mtime = idu_io_next_bits_id2ex_csr_hit_is_mtime; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mcycle = idu_io_next_bits_id2ex_csr_hit_is_mcycle; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_csr_hit_is_mhartid = idu_io_next_bits_id2ex_csr_hit_is_mhartid; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_signed = idu_io_next_bits_id2ex_mdu_op_mul_signed; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_is_mu = idu_io_next_bits_id2ex_mdu_op_is_mu; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_mul_32 = idu_io_next_bits_id2ex_mdu_op_mul_32; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_div_signed = idu_io_next_bits_id2ex_mdu_op_div_signed; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_is_div = idu_io_next_bits_id2ex_mdu_op_is_div; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mdu_op_is_du = idu_io_next_bits_id2ex_mdu_op_is_du; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_zimm = idu_io_next_bits_id2ex_zimm; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_intr = idu_io_next_bits_id2ex_intr; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_exec = idu_io_next_bits_id2ex_exec; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_mret = idu_io_next_bits_id2ex_mret; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_exce_code = idu_io_next_bits_id2ex_exce_code; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_pc = idu_io_next_bits_id2ex_pc; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2ex_is_iem = idu_io_next_bits_id2ex_is_iem; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_fencei = idu_io_next_bits_id2mem_fencei; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_size_byte = idu_io_next_bits_id2mem_size_byte; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_size_hword = idu_io_next_bits_id2mem_size_hword; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_size_word = idu_io_next_bits_id2mem_size_word; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_size_dword = idu_io_next_bits_id2mem_size_dword; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_sext_flag = idu_io_next_bits_id2mem_sext_flag; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_memory_rd_en = idu_io_next_bits_id2mem_memory_rd_en; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2mem_memory_we_en = idu_io_next_bits_id2mem_memory_we_en; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2wb_intr_exce_ret = idu_io_next_bits_id2wb_intr_exce_ret; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2wb_fencei = idu_io_next_bits_id2wb_fencei; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2wb_wb_sel = idu_io_next_bits_id2wb_wb_sel; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2wb_regfile_we_en = idu_io_next_bits_id2wb_regfile_we_en; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_prev_bits_id2wb_regfile_we_addr = idu_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 26:29 IDU.scala 296:10]
  assign ID2EXReg_io_next_ready = exu_io_prev_ready; // @[EXU.scala 161:17]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_prev_valid = ID2EXReg_io_next_valid; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_alu_src1 = ID2EXReg_io_next_bits_id2ex_alu_src1; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_alu_src2 = ID2EXReg_io_next_bits_id2ex_alu_src2; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_salu_src1 = ID2EXReg_io_next_bits_id2ex_salu_src1; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_salu_src2 = ID2EXReg_io_next_bits_id2ex_salu_src2; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_src1 = ID2EXReg_io_next_bits_id2ex_src1; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_src2 = ID2EXReg_io_next_bits_id2ex_src2; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_src3 = ID2EXReg_io_next_bits_id2ex_src3; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_auipc = ID2EXReg_io_next_bits_id2ex_operator_auipc; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_lui = ID2EXReg_io_next_bits_id2ex_operator_lui; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_jal = ID2EXReg_io_next_bits_id2ex_operator_jal; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_jalr = ID2EXReg_io_next_bits_id2ex_operator_jalr; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sb = ID2EXReg_io_next_bits_id2ex_operator_sb; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sh = ID2EXReg_io_next_bits_id2ex_operator_sh; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sw = ID2EXReg_io_next_bits_id2ex_operator_sw; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sd = ID2EXReg_io_next_bits_id2ex_operator_sd; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_add = ID2EXReg_io_next_bits_id2ex_operator_add; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sub = ID2EXReg_io_next_bits_id2ex_operator_sub; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sll = ID2EXReg_io_next_bits_id2ex_operator_sll; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_slt = ID2EXReg_io_next_bits_id2ex_operator_slt; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sltu = ID2EXReg_io_next_bits_id2ex_operator_sltu; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_xor = ID2EXReg_io_next_bits_id2ex_operator_xor; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_srl = ID2EXReg_io_next_bits_id2ex_operator_srl; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_sra = ID2EXReg_io_next_bits_id2ex_operator_sra; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_or = ID2EXReg_io_next_bits_id2ex_operator_or; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_and = ID2EXReg_io_next_bits_id2ex_operator_and; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_is_csr = ID2EXReg_io_next_bits_id2ex_operator_csr_is_csr; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrw = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrw; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrs = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrs; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrc = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrc; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrwi = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrwi; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrsi = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrsi; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_operator_csr_csrrci = ID2EXReg_io_next_bits_id2ex_operator_csr_csrrci; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_srcsize_byte = ID2EXReg_io_next_bits_id2ex_srcsize_byte; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_srcsize_hword = ID2EXReg_io_next_bits_id2ex_srcsize_hword; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_srcsize_word = ID2EXReg_io_next_bits_id2ex_srcsize_word; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_srcsize_dword = ID2EXReg_io_next_bits_id2ex_srcsize_dword; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_is_load = ID2EXReg_io_next_bits_id2ex_is_load; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_is_save = ID2EXReg_io_next_bits_id2ex_is_save; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_div_inf = ID2EXReg_io_next_bits_id2ex_div_inf; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_we = ID2EXReg_io_next_bits_id2ex_csr_we; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mepc = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mepc; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mtvec = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtvec; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mstatus = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mstatus; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mie = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mie; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mcause = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcause; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mip = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mip; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mtime = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mtime; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mcycle = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mcycle; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_csr_hit_is_mhartid = ID2EXReg_io_next_bits_id2ex_csr_hit_is_mhartid; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_mul_signed = ID2EXReg_io_next_bits_id2ex_mdu_op_mul_signed; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_is_mu = ID2EXReg_io_next_bits_id2ex_mdu_op_is_mu; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_mul_32 = ID2EXReg_io_next_bits_id2ex_mdu_op_mul_32; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_div_signed = ID2EXReg_io_next_bits_id2ex_mdu_op_div_signed; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_is_div = ID2EXReg_io_next_bits_id2ex_mdu_op_is_div; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mdu_op_is_du = ID2EXReg_io_next_bits_id2ex_mdu_op_is_du; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_zimm = ID2EXReg_io_next_bits_id2ex_zimm; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_intr = ID2EXReg_io_next_bits_id2ex_intr; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_exec = ID2EXReg_io_next_bits_id2ex_exec; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_mret = ID2EXReg_io_next_bits_id2ex_mret; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_exce_code = ID2EXReg_io_next_bits_id2ex_exce_code; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_pc = ID2EXReg_io_next_bits_id2ex_pc; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2ex_is_iem = ID2EXReg_io_next_bits_id2ex_is_iem; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_fencei = ID2EXReg_io_next_bits_id2mem_fencei; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_size_byte = ID2EXReg_io_next_bits_id2mem_size_byte; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_size_hword = ID2EXReg_io_next_bits_id2mem_size_hword; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_size_word = ID2EXReg_io_next_bits_id2mem_size_word; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_size_dword = ID2EXReg_io_next_bits_id2mem_size_dword; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_sext_flag = ID2EXReg_io_next_bits_id2mem_sext_flag; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_memory_rd_en = ID2EXReg_io_next_bits_id2mem_memory_rd_en; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2mem_memory_we_en = ID2EXReg_io_next_bits_id2mem_memory_we_en; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2wb_intr_exce_ret = ID2EXReg_io_next_bits_id2wb_intr_exce_ret; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2wb_fencei = ID2EXReg_io_next_bits_id2wb_fencei; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2wb_wb_sel = ID2EXReg_io_next_bits_id2wb_wb_sel; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2wb_regfile_we_en = ID2EXReg_io_next_bits_id2wb_regfile_we_en; // @[EXU.scala 161:17]
  assign exu_io_prev_bits_id2wb_regfile_we_addr = ID2EXReg_io_next_bits_id2wb_regfile_we_addr; // @[EXU.scala 161:17]
  assign exu_io_next_ready = EX2MEMReg_io_prev_ready; // @[Top.scala 27:29 MEMU.scala 85:23]
  assign exu_io_sb_clint_msip = io_sideband_clint_msip; // @[EXU.scala 159:15]
  assign exu_io_sb_clint_mtip = io_sideband_clint_mtip; // @[EXU.scala 159:15]
  assign exu_io_sb_clint_mtime = io_sideband_clint_mtime; // @[EXU.scala 159:15]
  assign exu_io_sb_meip = io_sideband_meip; // @[EXU.scala 159:15]
  assign EX2MEMReg_clock = clock;
  assign EX2MEMReg_reset = reset;
  assign EX2MEMReg_io_prev_valid = exu_io_next_valid; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_fencei = exu_io_next_bits_id2mem_fencei; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_size_byte = exu_io_next_bits_id2mem_size_byte; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_size_hword = exu_io_next_bits_id2mem_size_hword; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_size_word = exu_io_next_bits_id2mem_size_word; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_size_dword = exu_io_next_bits_id2mem_size_dword; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_sext_flag = exu_io_next_bits_id2mem_sext_flag; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_memory_rd_en = exu_io_next_bits_id2mem_memory_rd_en; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2mem_memory_we_en = exu_io_next_bits_id2mem_memory_we_en; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2wb_intr_exce_ret = exu_io_next_bits_id2wb_intr_exce_ret; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2wb_fencei = exu_io_next_bits_id2wb_fencei; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2wb_wb_sel = exu_io_next_bits_id2wb_wb_sel; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2wb_regfile_we_en = exu_io_next_bits_id2wb_regfile_we_en; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_id2wb_regfile_we_addr = exu_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_ex2mem_addr = exu_io_next_bits_ex2mem_addr; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_ex2mem_we_data = exu_io_next_bits_ex2mem_we_data; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_ex2mem_we_mask = exu_io_next_bits_ex2mem_we_mask; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_prev_bits_ex2wb_result_data = exu_io_next_bits_ex2wb_result_data; // @[Top.scala 27:29 EXU.scala 162:10]
  assign EX2MEMReg_io_next_ready = memu_io_prev_ready; // @[MEMU.scala 88:18]
  assign memu_clock = clock;
  assign memu_reset = reset;
  assign memu_io_prev_valid = EX2MEMReg_io_next_valid; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_fencei = EX2MEMReg_io_next_bits_id2mem_fencei; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_size_byte = EX2MEMReg_io_next_bits_id2mem_size_byte; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_size_hword = EX2MEMReg_io_next_bits_id2mem_size_hword; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_size_word = EX2MEMReg_io_next_bits_id2mem_size_word; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_size_dword = EX2MEMReg_io_next_bits_id2mem_size_dword; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_sext_flag = EX2MEMReg_io_next_bits_id2mem_sext_flag; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_memory_rd_en = EX2MEMReg_io_next_bits_id2mem_memory_rd_en; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2mem_memory_we_en = EX2MEMReg_io_next_bits_id2mem_memory_we_en; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2wb_intr_exce_ret = EX2MEMReg_io_next_bits_id2wb_intr_exce_ret; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2wb_fencei = EX2MEMReg_io_next_bits_id2wb_fencei; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2wb_wb_sel = EX2MEMReg_io_next_bits_id2wb_wb_sel; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2wb_regfile_we_en = EX2MEMReg_io_next_bits_id2wb_regfile_we_en; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_id2wb_regfile_we_addr = EX2MEMReg_io_next_bits_id2wb_regfile_we_addr; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_ex2mem_addr = EX2MEMReg_io_next_bits_ex2mem_addr; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_ex2mem_we_data = EX2MEMReg_io_next_bits_ex2mem_we_data; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_ex2mem_we_mask = EX2MEMReg_io_next_bits_ex2mem_we_mask; // @[MEMU.scala 88:18]
  assign memu_io_prev_bits_ex2wb_result_data = EX2MEMReg_io_next_bits_ex2wb_result_data; // @[MEMU.scala 88:18]
  assign memu_io_maxi_ar_ready = icon_io_memu_ar_ready; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_r_valid = icon_io_memu_r_valid; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_r_bits_data = icon_io_memu_r_bits_data; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_r_bits_last = icon_io_memu_r_bits_last; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_aw_ready = icon_io_memu_aw_ready; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_w_ready = icon_io_memu_w_ready; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_maxi_b_valid = icon_io_memu_b_valid; // @[Top.scala 39:28 AXI.scala 288:27]
  assign memu_io_mmio_ar_ready = icon_io_devu_ar_ready; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_r_valid = icon_io_devu_r_valid; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_r_bits_data = icon_io_devu_r_bits_data; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_r_bits_last = icon_io_devu_r_bits_last; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_aw_ready = icon_io_devu_aw_ready; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_w_ready = icon_io_devu_w_ready; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_mmio_b_valid = icon_io_devu_b_valid; // @[Top.scala 40:29 AXI.scala 289:27]
  assign memu_io_sram4_rdata = io_sram4_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 62:17]
  assign memu_io_sram5_rdata = io_sram5_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 63:17]
  assign memu_io_sram6_rdata = io_sram6_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 64:17]
  assign memu_io_sram7_rdata = io_sram7_rdata; // @[Top.scala 66:22 CacheBase.scala 76:11 Top.scala 65:17]
  assign memu_clint_rdata = clint_rdata;
  assign MEM2WBReg_clock = clock;
  assign MEM2WBReg_reset = reset;
  assign MEM2WBReg_io_prev_valid = memu_io_next_valid; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_id2wb_intr_exce_ret = memu_io_next_bits_id2wb_intr_exce_ret; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_id2wb_fencei = memu_io_next_bits_id2wb_fencei; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_id2wb_wb_sel = memu_io_next_bits_id2wb_wb_sel; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_id2wb_regfile_we_en = memu_io_next_bits_id2wb_regfile_we_en; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_id2wb_regfile_we_addr = memu_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_ex2wb_result_data = memu_io_next_bits_ex2wb_result_data; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign MEM2WBReg_io_prev_bits_mem2wb_memory_data = memu_io_next_bits_mem2wb_memory_data; // @[Top.scala 28:29 MEMU.scala 91:10]
  assign wbu_io__prev_valid = MEM2WBReg_io_next_valid; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_id2wb_intr_exce_ret = MEM2WBReg_io_next_bits_id2wb_intr_exce_ret; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_id2wb_fencei = MEM2WBReg_io_next_bits_id2wb_fencei; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_id2wb_wb_sel = MEM2WBReg_io_next_bits_id2wb_wb_sel; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_id2wb_regfile_we_en = MEM2WBReg_io_next_bits_id2wb_regfile_we_en; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_id2wb_regfile_we_addr = MEM2WBReg_io_next_bits_id2wb_regfile_we_addr; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_ex2wb_result_data = MEM2WBReg_io_next_bits_ex2wb_result_data; // @[WBU.scala 81:17]
  assign wbu_io__prev_bits_mem2wb_memory_data = MEM2WBReg_io_next_bits_mem2wb_memory_data; // @[WBU.scala 81:17]
  assign fwu_io_idu_optype_Itype = idu_io_fwu_optype_Itype; // @[Top.scala 29:29 IDU.scala 291:16]
  assign fwu_io_idu_src1_addr = idu_io_fwu_src1_addr; // @[Top.scala 29:29 IDU.scala 291:16]
  assign fwu_io_idu_src2_addr = idu_io_fwu_src2_addr; // @[Top.scala 29:29 IDU.scala 291:16]
  assign fwu_io_idu_src1_data = idu_io_fwu_src1_data; // @[Top.scala 29:29 IDU.scala 291:16]
  assign fwu_io_idu_src2_data = idu_io_fwu_src2_data; // @[Top.scala 29:29 IDU.scala 291:16]
  assign fwu_io_exu_is_load = ID2EXReg_io_next_bits_id2mem_memory_rd_en; // @[Top.scala 30:29 EXU.scala 164:17]
  assign fwu_io_exu_dst_addr = ID2EXReg_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 30:29 EXU.scala 165:18]
  assign fwu_io_exu_dst_data = exu_io_next_bits_ex2wb_result_data; // @[Top.scala 30:29 EXU.scala 166:18]
  assign fwu_io_memu_is_load_1 = memu_io_prev_bits_id2wb_wb_sel; // @[Top.scala 31:30 MEMU.scala 97:19]
  assign fwu_io_memu_dst_addr_1 = memu_io_prev_bits_id2wb_regfile_we_addr; // @[Top.scala 31:30 MEMU.scala 94:20]
  assign fwu_io_memu_dst_data_1 = memu_io_prev_bits_ex2wb_result_data; // @[Top.scala 31:30 MEMU.scala 96:20]
  assign fwu_io_memu_dst_addr_2 = memu_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 31:30 MEMU.scala 99:20]
  assign fwu_io_wbu_dst_addr = MEM2WBReg_io_next_bits_id2wb_regfile_we_addr; // @[Top.scala 32:30 WBU.scala 84:18]
  assign fwu_io_wbu_dst_data = wbu_io__regfile_data; // @[Top.scala 32:30 WBU.scala 85:18]
  assign bru_clock = clock;
  assign bru_reset = reset;
  assign bru_io_idu_brh = idu_io_bru_brh; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_jal = idu_io_bru_jal; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_jalr = idu_io_bru_jalr; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_pc = idu_io_bru_pc; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_src1 = idu_io_bru_src1; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_src2 = idu_io_bru_src2; // @[Top.scala 24:29 IDU.scala 292:16]
  assign bru_io_idu_imm = idu_io_bru_imm; // @[Top.scala 24:29 IDU.scala 292:16]
  assign regfile_clock = clock;
  assign regfile_reset = reset;
  assign regfile_io_wbu_en = wbu_io__regfile_en; // @[Top.scala 36:34 WBU.scala 82:13]
  assign regfile_io_wbu_addr = wbu_io__regfile_addr; // @[Top.scala 36:34 WBU.scala 82:13]
  assign regfile_io_wbu_data = wbu_io__regfile_data; // @[Top.scala 36:34 WBU.scala 82:13]
  assign regfile_io_idu_addr1 = idu_io_regfile_addr1; // @[Top.scala 35:34 IDU.scala 293:20]
  assign regfile_io_idu_addr2 = idu_io_regfile_addr2; // @[Top.scala 35:34 IDU.scala 293:20]
  always @(posedge clock) begin
    sram_init_reg <= reset | _GEN_52; // @[Top.scala 42:38 Top.scala 42:38]
    if (reset) begin // @[Counter.scala 60:40]
      sram_init_cnt <= 6'h0; // @[Counter.scala 60:40]
    end else if (sram_init_reg) begin // @[Counter.scala 118:17]
      sram_init_cnt <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sram_init_reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sram_init_cnt = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978_CLINT(
  input         clock,
  input         reset,
  output        io_sideband_msip,
  output        io_sideband_mtip,
  output [63:0] io_sideband_mtime,
  input         clint_we_0,
  input  [31:0] clint_addr,
  output [63:0] clint_rdata_0,
  input  [63:0] clint_wdata_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[CLINT.scala 28:34]
  reg [63:0] mtimecmp; // @[CLINT.scala 29:34]
  reg [63:0] msip; // @[CLINT.scala 30:34]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[CLINT.scala 31:18]
  wire  _GEN_0 = ~(|clint_addr[2:0]) ? clint_addr[31:3] == 29'h4017ff : clint_addr[31:3] == 29'h4017ff; // @[CLINT.scala 51:33 CLINT.scala 52:18 CLINT.scala 48:16]
  wire  _GEN_1 = ~(|clint_addr[2:0]) ? clint_addr[31:3] == 29'h400800 : clint_addr[31:3] == 29'h400800; // @[CLINT.scala 51:33 CLINT.scala 53:18 CLINT.scala 49:16]
  wire  _GEN_2 = ~(|clint_addr[2:0]) ? clint_addr[31:3] == 29'h400000 : clint_addr[31:3] == 29'h400000; // @[CLINT.scala 51:33 CLINT.scala 54:18 CLINT.scala 50:16]
  wire [63:0] _GEN_4 = clint_we_0 ? 64'h0 : mtime; // @[CLINT.scala 62:19 CLINT.scala 65:19]
  wire [63:0] _GEN_6 = _GEN_0 ? _GEN_4 : 64'h0; // @[CLINT.scala 61:17]
  wire [63:0] _GEN_8 = clint_we_0 ? _GEN_6 : mtimecmp; // @[CLINT.scala 69:19 CLINT.scala 72:19]
  wire [63:0] _GEN_10 = _GEN_1 ? _GEN_8 : _GEN_6; // @[CLINT.scala 68:20]
  wire [63:0] _GEN_12 = clint_we_0 ? _GEN_10 : msip; // @[CLINT.scala 76:19 CLINT.scala 79:19]
  wire [63:0] clint_rdata = _GEN_2 ? _GEN_12 : _GEN_10; // @[CLINT.scala 75:17]
  assign io_sideband_msip = msip[0]; // @[CLINT.scala 33:20]
  assign io_sideband_mtip = mtime >= mtimecmp; // @[CLINT.scala 35:23]
  assign io_sideband_mtime = mtime; // @[CLINT.scala 34:13]
  assign clint_rdata_0 = clint_rdata;
  always @(posedge clock) begin
    if (reset) begin // @[CLINT.scala 28:34]
      mtime <= 64'h0; // @[CLINT.scala 28:34]
    end else if (_GEN_0) begin // @[CLINT.scala 61:17]
      if (clint_we_0) begin // @[CLINT.scala 62:19]
        mtime <= clint_wdata_1; // @[CLINT.scala 63:13]
      end else begin
        mtime <= _mtime_T_1; // @[CLINT.scala 31:9]
      end
    end else begin
      mtime <= _mtime_T_1; // @[CLINT.scala 31:9]
    end
    if (reset) begin // @[CLINT.scala 29:34]
      mtimecmp <= 64'h0; // @[CLINT.scala 29:34]
    end else if (_GEN_1) begin // @[CLINT.scala 68:20]
      if (clint_we_0) begin // @[CLINT.scala 69:19]
        mtimecmp <= clint_wdata_1; // @[CLINT.scala 70:16]
      end
    end
    if (reset) begin // @[CLINT.scala 30:34]
      msip <= 64'h0; // @[CLINT.scala 30:34]
    end else if (_GEN_2) begin // @[CLINT.scala 75:17]
      if (clint_we_0) begin // @[CLINT.scala 76:19]
        msip <= clint_wdata_1; // @[CLINT.scala 77:12]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  msip = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_040978(
  input          clock,
  input          reset,
  input          io_master_arready,
  output         io_master_arvalid,
  output [31:0]  io_master_araddr,
  output [3:0]   io_master_arid,
  output [7:0]   io_master_arlen,
  output [2:0]   io_master_arsize,
  output [1:0]   io_master_arburst,
  output         io_master_rready,
  input          io_master_rvalid,
  input  [1:0]   io_master_rresp,
  input  [63:0]  io_master_rdata,
  input          io_master_rlast,
  input  [3:0]   io_master_rid,
  input          io_master_awready,
  output         io_master_awvalid,
  output [31:0]  io_master_awaddr,
  output [3:0]   io_master_awid,
  output [7:0]   io_master_awlen,
  output [2:0]   io_master_awsize,
  output [1:0]   io_master_awburst,
  input          io_master_wready,
  output         io_master_wvalid,
  output [63:0]  io_master_wdata,
  output [7:0]   io_master_wstrb,
  output         io_master_wlast,
  output         io_master_bready,
  input          io_master_bvalid,
  input  [1:0]   io_master_bresp,
  input  [3:0]   io_master_bid,
  output         io_slave_arready,
  input          io_slave_arvalid,
  input  [31:0]  io_slave_araddr,
  input  [3:0]   io_slave_arid,
  input  [7:0]   io_slave_arlen,
  input  [2:0]   io_slave_arsize,
  input  [1:0]   io_slave_arburst,
  input          io_slave_rready,
  output         io_slave_rvalid,
  output [1:0]   io_slave_rresp,
  output [63:0]  io_slave_rdata,
  output         io_slave_rlast,
  output [3:0]   io_slave_rid,
  output         io_slave_awready,
  input          io_slave_awvalid,
  input  [31:0]  io_slave_awaddr,
  input  [3:0]   io_slave_awid,
  input  [7:0]   io_slave_awlen,
  input  [2:0]   io_slave_awsize,
  input  [1:0]   io_slave_awburst,
  output         io_slave_wready,
  input          io_slave_wvalid,
  input  [63:0]  io_slave_wdata,
  input  [7:0]   io_slave_wstrb,
  input          io_slave_wlast,
  input          io_slave_bready,
  output         io_slave_bvalid,
  output [1:0]   io_slave_bresp,
  output [3:0]   io_slave_bid,
  input          io_interrupt,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata
);
  wire  core_clock; // @[Top.scala 101:28]
  wire  core_reset; // @[Top.scala 101:28]
  wire  core_io_maxi4_ar_ready; // @[Top.scala 101:28]
  wire  core_io_maxi4_ar_valid; // @[Top.scala 101:28]
  wire [31:0] core_io_maxi4_ar_bits_addr; // @[Top.scala 101:28]
  wire [1:0] core_io_maxi4_ar_bits_burst; // @[Top.scala 101:28]
  wire [3:0] core_io_maxi4_ar_bits_id; // @[Top.scala 101:28]
  wire [7:0] core_io_maxi4_ar_bits_len; // @[Top.scala 101:28]
  wire [2:0] core_io_maxi4_ar_bits_size; // @[Top.scala 101:28]
  wire  core_io_maxi4_r_ready; // @[Top.scala 101:28]
  wire  core_io_maxi4_r_valid; // @[Top.scala 101:28]
  wire [63:0] core_io_maxi4_r_bits_data; // @[Top.scala 101:28]
  wire [3:0] core_io_maxi4_r_bits_id; // @[Top.scala 101:28]
  wire  core_io_maxi4_r_bits_last; // @[Top.scala 101:28]
  wire [1:0] core_io_maxi4_r_bits_resp; // @[Top.scala 101:28]
  wire  core_io_maxi4_aw_ready; // @[Top.scala 101:28]
  wire  core_io_maxi4_aw_valid; // @[Top.scala 101:28]
  wire [31:0] core_io_maxi4_aw_bits_addr; // @[Top.scala 101:28]
  wire [1:0] core_io_maxi4_aw_bits_burst; // @[Top.scala 101:28]
  wire [3:0] core_io_maxi4_aw_bits_id; // @[Top.scala 101:28]
  wire [7:0] core_io_maxi4_aw_bits_len; // @[Top.scala 101:28]
  wire [2:0] core_io_maxi4_aw_bits_size; // @[Top.scala 101:28]
  wire  core_io_maxi4_w_ready; // @[Top.scala 101:28]
  wire  core_io_maxi4_w_valid; // @[Top.scala 101:28]
  wire [63:0] core_io_maxi4_w_bits_data; // @[Top.scala 101:28]
  wire [7:0] core_io_maxi4_w_bits_strb; // @[Top.scala 101:28]
  wire  core_io_maxi4_w_bits_last; // @[Top.scala 101:28]
  wire  core_io_maxi4_b_ready; // @[Top.scala 101:28]
  wire  core_io_maxi4_b_valid; // @[Top.scala 101:28]
  wire [3:0] core_io_maxi4_b_bits_id; // @[Top.scala 101:28]
  wire [1:0] core_io_maxi4_b_bits_resp; // @[Top.scala 101:28]
  wire  core_io_sideband_clint_msip; // @[Top.scala 101:28]
  wire  core_io_sideband_clint_mtip; // @[Top.scala 101:28]
  wire [63:0] core_io_sideband_clint_mtime; // @[Top.scala 101:28]
  wire  core_io_sideband_meip; // @[Top.scala 101:28]
  wire [5:0] core_io_sram0_addr; // @[Top.scala 101:28]
  wire  core_io_sram0_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram0_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram0_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram0_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram1_addr; // @[Top.scala 101:28]
  wire  core_io_sram1_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram1_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram1_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram1_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram2_addr; // @[Top.scala 101:28]
  wire  core_io_sram2_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram2_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram2_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram2_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram3_addr; // @[Top.scala 101:28]
  wire  core_io_sram3_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram3_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram3_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram3_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram4_addr; // @[Top.scala 101:28]
  wire  core_io_sram4_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram4_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram4_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram4_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram5_addr; // @[Top.scala 101:28]
  wire  core_io_sram5_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram5_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram5_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram5_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram6_addr; // @[Top.scala 101:28]
  wire  core_io_sram6_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram6_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram6_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram6_rdata; // @[Top.scala 101:28]
  wire [5:0] core_io_sram7_addr; // @[Top.scala 101:28]
  wire  core_io_sram7_wen; // @[Top.scala 101:28]
  wire [127:0] core_io_sram7_wmask; // @[Top.scala 101:28]
  wire [127:0] core_io_sram7_wdata; // @[Top.scala 101:28]
  wire [127:0] core_io_sram7_rdata; // @[Top.scala 101:28]
  wire  core_clint_we; // @[Top.scala 101:28]
  wire [31:0] core__T_24; // @[Top.scala 101:28]
  wire [63:0] core_clint_rdata; // @[Top.scala 101:28]
  wire [63:0] core_clint_wdata; // @[Top.scala 101:28]
  wire  clint_clock; // @[Top.scala 149:29]
  wire  clint_reset; // @[Top.scala 149:29]
  wire  clint_io_sideband_msip; // @[Top.scala 149:29]
  wire  clint_io_sideband_mtip; // @[Top.scala 149:29]
  wire [63:0] clint_io_sideband_mtime; // @[Top.scala 149:29]
  wire  clint_clint_we_0; // @[Top.scala 149:29]
  wire [31:0] clint_clint_addr; // @[Top.scala 149:29]
  wire [63:0] clint_clint_rdata_0; // @[Top.scala 149:29]
  wire [63:0] clint_clint_wdata_1; // @[Top.scala 149:29]
  ysyx_040978_SparkCore core ( // @[Top.scala 101:28]
    .clock(core_clock),
    .reset(core_reset),
    .io_maxi4_ar_ready(core_io_maxi4_ar_ready),
    .io_maxi4_ar_valid(core_io_maxi4_ar_valid),
    .io_maxi4_ar_bits_addr(core_io_maxi4_ar_bits_addr),
    .io_maxi4_ar_bits_burst(core_io_maxi4_ar_bits_burst),
    .io_maxi4_ar_bits_id(core_io_maxi4_ar_bits_id),
    .io_maxi4_ar_bits_len(core_io_maxi4_ar_bits_len),
    .io_maxi4_ar_bits_size(core_io_maxi4_ar_bits_size),
    .io_maxi4_r_ready(core_io_maxi4_r_ready),
    .io_maxi4_r_valid(core_io_maxi4_r_valid),
    .io_maxi4_r_bits_data(core_io_maxi4_r_bits_data),
    .io_maxi4_r_bits_id(core_io_maxi4_r_bits_id),
    .io_maxi4_r_bits_last(core_io_maxi4_r_bits_last),
    .io_maxi4_r_bits_resp(core_io_maxi4_r_bits_resp),
    .io_maxi4_aw_ready(core_io_maxi4_aw_ready),
    .io_maxi4_aw_valid(core_io_maxi4_aw_valid),
    .io_maxi4_aw_bits_addr(core_io_maxi4_aw_bits_addr),
    .io_maxi4_aw_bits_burst(core_io_maxi4_aw_bits_burst),
    .io_maxi4_aw_bits_id(core_io_maxi4_aw_bits_id),
    .io_maxi4_aw_bits_len(core_io_maxi4_aw_bits_len),
    .io_maxi4_aw_bits_size(core_io_maxi4_aw_bits_size),
    .io_maxi4_w_ready(core_io_maxi4_w_ready),
    .io_maxi4_w_valid(core_io_maxi4_w_valid),
    .io_maxi4_w_bits_data(core_io_maxi4_w_bits_data),
    .io_maxi4_w_bits_strb(core_io_maxi4_w_bits_strb),
    .io_maxi4_w_bits_last(core_io_maxi4_w_bits_last),
    .io_maxi4_b_ready(core_io_maxi4_b_ready),
    .io_maxi4_b_valid(core_io_maxi4_b_valid),
    .io_maxi4_b_bits_id(core_io_maxi4_b_bits_id),
    .io_maxi4_b_bits_resp(core_io_maxi4_b_bits_resp),
    .io_sideband_clint_msip(core_io_sideband_clint_msip),
    .io_sideband_clint_mtip(core_io_sideband_clint_mtip),
    .io_sideband_clint_mtime(core_io_sideband_clint_mtime),
    .io_sideband_meip(core_io_sideband_meip),
    .io_sram0_addr(core_io_sram0_addr),
    .io_sram0_wen(core_io_sram0_wen),
    .io_sram0_wmask(core_io_sram0_wmask),
    .io_sram0_wdata(core_io_sram0_wdata),
    .io_sram0_rdata(core_io_sram0_rdata),
    .io_sram1_addr(core_io_sram1_addr),
    .io_sram1_wen(core_io_sram1_wen),
    .io_sram1_wmask(core_io_sram1_wmask),
    .io_sram1_wdata(core_io_sram1_wdata),
    .io_sram1_rdata(core_io_sram1_rdata),
    .io_sram2_addr(core_io_sram2_addr),
    .io_sram2_wen(core_io_sram2_wen),
    .io_sram2_wmask(core_io_sram2_wmask),
    .io_sram2_wdata(core_io_sram2_wdata),
    .io_sram2_rdata(core_io_sram2_rdata),
    .io_sram3_addr(core_io_sram3_addr),
    .io_sram3_wen(core_io_sram3_wen),
    .io_sram3_wmask(core_io_sram3_wmask),
    .io_sram3_wdata(core_io_sram3_wdata),
    .io_sram3_rdata(core_io_sram3_rdata),
    .io_sram4_addr(core_io_sram4_addr),
    .io_sram4_wen(core_io_sram4_wen),
    .io_sram4_wmask(core_io_sram4_wmask),
    .io_sram4_wdata(core_io_sram4_wdata),
    .io_sram4_rdata(core_io_sram4_rdata),
    .io_sram5_addr(core_io_sram5_addr),
    .io_sram5_wen(core_io_sram5_wen),
    .io_sram5_wmask(core_io_sram5_wmask),
    .io_sram5_wdata(core_io_sram5_wdata),
    .io_sram5_rdata(core_io_sram5_rdata),
    .io_sram6_addr(core_io_sram6_addr),
    .io_sram6_wen(core_io_sram6_wen),
    .io_sram6_wmask(core_io_sram6_wmask),
    .io_sram6_wdata(core_io_sram6_wdata),
    .io_sram6_rdata(core_io_sram6_rdata),
    .io_sram7_addr(core_io_sram7_addr),
    .io_sram7_wen(core_io_sram7_wen),
    .io_sram7_wmask(core_io_sram7_wmask),
    .io_sram7_wdata(core_io_sram7_wdata),
    .io_sram7_rdata(core_io_sram7_rdata),
    .clint_we(core_clint_we),
    ._T_24(core__T_24),
    .clint_rdata(core_clint_rdata),
    .clint_wdata(core_clint_wdata)
  );
  ysyx_040978_CLINT clint ( // @[Top.scala 149:29]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_sideband_msip(clint_io_sideband_msip),
    .io_sideband_mtip(clint_io_sideband_mtip),
    .io_sideband_mtime(clint_io_sideband_mtime),
    .clint_we_0(clint_clint_we_0),
    .clint_addr(clint_clint_addr),
    .clint_rdata_0(clint_clint_rdata_0),
    .clint_wdata_1(clint_clint_wdata_1)
  );
  assign io_master_arvalid = core_io_maxi4_ar_valid; // @[Top.scala 119:22]
  assign io_master_araddr = core_io_maxi4_ar_bits_addr; // @[Top.scala 116:22]
  assign io_master_arid = core_io_maxi4_ar_bits_id; // @[Top.scala 114:22]
  assign io_master_arlen = core_io_maxi4_ar_bits_len; // @[Top.scala 115:22]
  assign io_master_arsize = core_io_maxi4_ar_bits_size; // @[Top.scala 117:22]
  assign io_master_arburst = core_io_maxi4_ar_bits_burst; // @[Top.scala 118:22]
  assign io_master_rready = core_io_maxi4_r_ready; // @[Top.scala 126:26]
  assign io_master_awvalid = core_io_maxi4_aw_valid; // @[Top.scala 107:21]
  assign io_master_awaddr = core_io_maxi4_aw_bits_addr; // @[Top.scala 104:20]
  assign io_master_awid = core_io_maxi4_aw_bits_id; // @[Top.scala 102:18]
  assign io_master_awlen = core_io_maxi4_aw_bits_len; // @[Top.scala 103:19]
  assign io_master_awsize = core_io_maxi4_aw_bits_size; // @[Top.scala 105:20]
  assign io_master_awburst = core_io_maxi4_aw_bits_burst; // @[Top.scala 106:21]
  assign io_master_wvalid = core_io_maxi4_w_valid; // @[Top.scala 132:20]
  assign io_master_wdata = core_io_maxi4_w_bits_data; // @[Top.scala 129:19]
  assign io_master_wstrb = core_io_maxi4_w_bits_strb; // @[Top.scala 131:19]
  assign io_master_wlast = core_io_maxi4_w_bits_last; // @[Top.scala 130:19]
  assign io_master_bready = core_io_maxi4_b_ready; // @[Top.scala 138:20]
  assign io_slave_arready = 1'h0; // @[YSYXSoC3.scala 61:18]
  assign io_slave_rvalid = 1'h0; // @[YSYXSoC3.scala 84:18]
  assign io_slave_rresp = 2'h0; // @[YSYXSoC3.scala 85:18]
  assign io_slave_rdata = 64'h0; // @[YSYXSoC3.scala 86:18]
  assign io_slave_rlast = 1'h0; // @[YSYXSoC3.scala 87:18]
  assign io_slave_rid = 4'h0; // @[YSYXSoC3.scala 88:18]
  assign io_slave_awready = 1'h0; // @[YSYXSoC3.scala 71:18]
  assign io_slave_wready = 1'h0; // @[YSYXSoC3.scala 79:17]
  assign io_slave_bvalid = 1'h0; // @[YSYXSoC3.scala 93:18]
  assign io_slave_bresp = 2'h0; // @[YSYXSoC3.scala 94:18]
  assign io_slave_bid = 4'h0; // @[YSYXSoC3.scala 95:18]
  assign io_sram0_addr = core_io_sram0_addr; // @[Top.scala 140:17]
  assign io_sram0_cen = 1'h0; // @[Top.scala 140:17]
  assign io_sram0_wen = core_io_sram0_wen; // @[Top.scala 140:17]
  assign io_sram0_wmask = core_io_sram0_wmask; // @[Top.scala 140:17]
  assign io_sram0_wdata = core_io_sram0_wdata; // @[Top.scala 140:17]
  assign io_sram1_addr = core_io_sram1_addr; // @[Top.scala 141:17]
  assign io_sram1_cen = 1'h0; // @[Top.scala 141:17]
  assign io_sram1_wen = core_io_sram1_wen; // @[Top.scala 141:17]
  assign io_sram1_wmask = core_io_sram1_wmask; // @[Top.scala 141:17]
  assign io_sram1_wdata = core_io_sram1_wdata; // @[Top.scala 141:17]
  assign io_sram2_addr = core_io_sram2_addr; // @[Top.scala 142:17]
  assign io_sram2_cen = 1'h0; // @[Top.scala 142:17]
  assign io_sram2_wen = core_io_sram2_wen; // @[Top.scala 142:17]
  assign io_sram2_wmask = core_io_sram2_wmask; // @[Top.scala 142:17]
  assign io_sram2_wdata = core_io_sram2_wdata; // @[Top.scala 142:17]
  assign io_sram3_addr = core_io_sram3_addr; // @[Top.scala 143:17]
  assign io_sram3_cen = 1'h0; // @[Top.scala 143:17]
  assign io_sram3_wen = core_io_sram3_wen; // @[Top.scala 143:17]
  assign io_sram3_wmask = core_io_sram3_wmask; // @[Top.scala 143:17]
  assign io_sram3_wdata = core_io_sram3_wdata; // @[Top.scala 143:17]
  assign io_sram4_addr = core_io_sram4_addr; // @[Top.scala 144:17]
  assign io_sram4_cen = 1'h0; // @[Top.scala 144:17]
  assign io_sram4_wen = core_io_sram4_wen; // @[Top.scala 144:17]
  assign io_sram4_wmask = core_io_sram4_wmask; // @[Top.scala 144:17]
  assign io_sram4_wdata = core_io_sram4_wdata; // @[Top.scala 144:17]
  assign io_sram5_addr = core_io_sram5_addr; // @[Top.scala 145:17]
  assign io_sram5_cen = 1'h0; // @[Top.scala 145:17]
  assign io_sram5_wen = core_io_sram5_wen; // @[Top.scala 145:17]
  assign io_sram5_wmask = core_io_sram5_wmask; // @[Top.scala 145:17]
  assign io_sram5_wdata = core_io_sram5_wdata; // @[Top.scala 145:17]
  assign io_sram6_addr = core_io_sram6_addr; // @[Top.scala 146:17]
  assign io_sram6_cen = 1'h0; // @[Top.scala 146:17]
  assign io_sram6_wen = core_io_sram6_wen; // @[Top.scala 146:17]
  assign io_sram6_wmask = core_io_sram6_wmask; // @[Top.scala 146:17]
  assign io_sram6_wdata = core_io_sram6_wdata; // @[Top.scala 146:17]
  assign io_sram7_addr = core_io_sram7_addr; // @[Top.scala 147:17]
  assign io_sram7_cen = 1'h0; // @[Top.scala 147:17]
  assign io_sram7_wen = core_io_sram7_wen; // @[Top.scala 147:17]
  assign io_sram7_wmask = core_io_sram7_wmask; // @[Top.scala 147:17]
  assign io_sram7_wdata = core_io_sram7_wdata; // @[Top.scala 147:17]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_maxi4_ar_ready = io_master_arready; // @[Top.scala 120:26]
  assign core_io_maxi4_r_valid = io_master_rvalid; // @[Top.scala 127:29]
  assign core_io_maxi4_r_bits_data = io_master_rdata; // @[Top.scala 123:29]
  assign core_io_maxi4_r_bits_id = io_master_rid; // @[Top.scala 122:29]
  assign core_io_maxi4_r_bits_last = io_master_rlast; // @[Top.scala 125:29]
  assign core_io_maxi4_r_bits_resp = io_master_rresp; // @[Top.scala 124:29]
  assign core_io_maxi4_aw_ready = io_master_awready; // @[Top.scala 108:26]
  assign core_io_maxi4_w_ready = io_master_wready; // @[Top.scala 133:25]
  assign core_io_maxi4_b_valid = io_master_bvalid; // @[Top.scala 137:25]
  assign core_io_maxi4_b_bits_id = io_master_bid; // @[Top.scala 135:27]
  assign core_io_maxi4_b_bits_resp = io_master_bresp; // @[Top.scala 136:29]
  assign core_io_sideband_clint_msip = clint_io_sideband_msip; // @[Top.scala 150:26]
  assign core_io_sideband_clint_mtip = clint_io_sideband_mtip; // @[Top.scala 150:26]
  assign core_io_sideband_clint_mtime = clint_io_sideband_mtime; // @[Top.scala 150:26]
  assign core_io_sideband_meip = io_interrupt; // @[Top.scala 151:25]
  assign core_io_sram0_rdata = io_sram0_rdata; // @[Top.scala 140:17]
  assign core_io_sram1_rdata = io_sram1_rdata; // @[Top.scala 141:17]
  assign core_io_sram2_rdata = io_sram2_rdata; // @[Top.scala 142:17]
  assign core_io_sram3_rdata = io_sram3_rdata; // @[Top.scala 143:17]
  assign core_io_sram4_rdata = io_sram4_rdata; // @[Top.scala 144:17]
  assign core_io_sram5_rdata = io_sram5_rdata; // @[Top.scala 145:17]
  assign core_io_sram6_rdata = io_sram6_rdata; // @[Top.scala 146:17]
  assign core_io_sram7_rdata = io_sram7_rdata; // @[Top.scala 147:17]
  assign core_clint_rdata = clint_clint_rdata_0;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_clint_we_0 = core_clint_we;
  assign clint_clint_addr = core__T_24;
  assign clint_clint_wdata_1 = core_clint_wdata;
endmodule
`timescale 1ps/1ps

//MuxKey 模块实现了“键值选择”功能，即
//在一个 (键值，数据) 的列表 lut 中，
//根据给定的键值 key ，将 out 设置为与其匹配的数据。
//若列表中不存在键值为 key 的数据，则 out 为 0 。
//特别地， MuxKeyWithDefault 模块可以提供一个默认值 default_out ，
//当列表中不存在键值为 key 的数据，则 out 为 default_out 。
//实例化这两个模块时需要注意如下两点：
//
//  1.需要使用者提供键值对的数量 NR_KEY，键值的位宽 KEY_LEN 
//  以及数据的位宽 DATA_LEN 这三个参数，并保证端口的信号宽度与
//  提供的参数一致，否则将会输出错误的结果
//  2.若列表中存在多个键值为 key 的数据，则 out 的值是未定义的，
//  需要使用者来保证列表中的键值互不相同


module ysyx_040978_MuxKey #(NR_KEY = 2, KEY_LEN = 1, DATA_LEN = 1) (
  output [DATA_LEN-1:0] out,
  input [KEY_LEN-1:0] key,
  input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
);
  ysyx_040978_MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 0) i0 (out, key, {DATA_LEN{1'b0}}, lut);
endmodule`timescale 1ps/1ps

module ysyx_040978_MuxKeyWithDefault #(NR_KEY = 2, KEY_LEN = 1, DATA_LEN = 1) (
  output [DATA_LEN-1:0] out,
  input [KEY_LEN-1:0] key,
  input [DATA_LEN-1:0] default_out,
  input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
);
  ysyx_040978_MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 1) i0 (out, key, default_out, lut);
endmodule`timescale 1ps/1ps

//MuxKeyInternal 模块的实现中用到了很多高级的功能，
//如 generate 和 for 循环等，
//为了方便编写还使用了行为建模方式，在这里我们不展开介绍，
//通过结构化建模的抽象，使用者可以无需关心这些细节


module ysyx_040978_MuxKeyInternal #(NR_KEY = 2, KEY_LEN = 1, DATA_LEN = 1, HAS_DEFAULT = 0) (
  output reg [DATA_LEN-1:0] out,
  input [KEY_LEN-1:0] key,
  input [DATA_LEN-1:0] default_out,
  input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
);

  localparam PAIR_LEN = KEY_LEN + DATA_LEN;
  wire [PAIR_LEN-1:0] pair_list [NR_KEY-1:0];
  wire [KEY_LEN-1:0] key_list [NR_KEY-1:0];
  wire [DATA_LEN-1:0] data_list [NR_KEY-1:0];

  generate
    for (genvar n = 0; n < NR_KEY; n = n + 1) begin
      assign pair_list[n] = lut[PAIR_LEN*(n+1)-1 : PAIR_LEN*n];
      assign data_list[n] = pair_list[n][DATA_LEN-1:0];
      assign key_list[n]  = pair_list[n][PAIR_LEN-1:DATA_LEN];
    end
  endgenerate

  reg [DATA_LEN-1 : 0] lut_out;
  reg hit;
  integer i;
  always @(*) begin
    lut_out = 0;
    hit = 0;
    for (i = 0; i < NR_KEY; i = i + 1) begin
      lut_out = lut_out | ({DATA_LEN{key == key_list[i]}} & data_list[i]);
      hit = hit | (key == key_list[i]);
    end
    if (!HAS_DEFAULT) out = lut_out;
    else out = (hit ? lut_out : default_out);
  end

endmodule