module ysyx_040656_mul_YDecoder (
    input  yc,
    input  yb,
    input  ya,
    output negx,
    output x,
    output neg2x,
    output _2x
);
  assign negx  = (yc & yb & ~ya) | (yc & ~yb & ya);
  assign x     = (~yc & ~yb & ya) | (~yc & yb & ~ya);
  assign neg2x = (yc & ~yb & ~ya);
  assign _2x   = (~yc & yb & ya);
endmodule
module ysyx_040656_mul_BoothBase (
    input  negx,
    input  x,
    input  neg2x,
    input  _2x,
    input  InX,
    input  PosLastX,
    input  NegLastX,
    output PosNextX,
    output NegNextX,
    output OutX
);
  assign OutX     = (negx & ~InX) | (x & InX) | (neg2x & NegLastX) | (_2x & PosLastX);
  assign PosNextX = InX;
  assign NegNextX = ~InX;
endmodule
module ysyx_040656_mul_BoothInterBase (
    input [2:0] y,
    input [63:0] InX,
    output [63:0] OutX,
    output Carry
);
  wire negx, x, neg2x, _2x;
  wire [1:0] CarrySig[65];
  ysyx_040656_mul_YDecoder uu (
      .yc(y[2]),
      .yb(y[1]),
      .ya(y[0]),
      .negx(negx),
      .x(x),
      .neg2x(neg2x),
      ._2x(_2x)
  );
  ysyx_040656_mul_BoothBase fir (
      .negx(negx),
      .x(x),
      .neg2x(neg2x),
      ._2x(_2x),
      .InX(InX[0]),
      .PosLastX(1'b0),
      .NegLastX(1'b1),
      .PosNextX(CarrySig[1][0]),
      .NegNextX(CarrySig[1][1]),
      .OutX(OutX[0])
  );
  generate
    genvar i;
    for (i = 1; i < 64; i = i + 1) begin : g_for
      ysyx_040656_mul_BoothBase ui (
          .negx(negx),
          .x(x),
          .neg2x(neg2x),
          ._2x(_2x),
          .InX(InX[i]),
          .PosLastX(CarrySig[i][0]),
          .NegLastX(CarrySig[i][1]),
          .PosNextX(CarrySig[i+1][0]),
          .NegNextX(CarrySig[i+1][1]),
          .OutX(OutX[i])
      );
    end
  endgenerate
  assign Carry = negx || neg2x;
endmodule
module ysyx_040656_mul_addr (
    input  A,
    input  B,
    input  C,
    output Carry,
    output S
);
  assign S     = ~A & ~B & C | ~A & B & ~C | A & ~B & ~C | A & B & C;
  assign Carry = A & B | A & C | B & C;
endmodule
module ysyx_040656_mul_WallaceTreeBase (
    input [16:0] InData,
    input [13:0] CIn,
    output [13:0] COut,
    output C,
    output S
);
  wire [4:0] FirSig;
  ysyx_040656_mul_addr first1 (
      .A(InData[4]),
      .B(InData[3]),
      .C(InData[2]),
      .Carry(COut[0]),
      .S(FirSig[0])
  );
  ysyx_040656_mul_addr first2 (
      .A(InData[7]),
      .B(InData[6]),
      .C(InData[5]),
      .Carry(COut[1]),
      .S(FirSig[1])
  );
  ysyx_040656_mul_addr first3 (
      .A(InData[10]),
      .B(InData[9]),
      .C(InData[8]),
      .Carry(COut[2]),
      .S(FirSig[2])
  );
  ysyx_040656_mul_addr first4 (
      .A(InData[13]),
      .B(InData[12]),
      .C(InData[11]),
      .Carry(COut[3]),
      .S(FirSig[3])
  );
  ysyx_040656_mul_addr first5 (
      .A(InData[16]),
      .B(InData[15]),
      .C(InData[14]),
      .Carry(COut[4]),
      .S(FirSig[4])
  );
  wire [3:0] SecSig;
  ysyx_040656_mul_addr second1 (
      .A(CIn[2]),
      .B(CIn[1]),
      .C(CIn[0]),
      .Carry(COut[5]),
      .S(SecSig[0])
  );
  ysyx_040656_mul_addr second2 (
      .A(InData[0]),
      .B(CIn[4]),
      .C(CIn[3]),
      .Carry(COut[6]),
      .S(SecSig[1])
  );
  ysyx_040656_mul_addr second3 (
      .A(FirSig[1]),
      .B(FirSig[0]),
      .C(InData[1]),
      .Carry(COut[7]),
      .S(SecSig[2])
  );
  ysyx_040656_mul_addr second4 (
      .A(FirSig[4]),
      .B(FirSig[3]),
      .C(FirSig[2]),
      .Carry(COut[8]),
      .S(SecSig[3])
  );
  wire [1:0] ThiSig;
  ysyx_040656_mul_addr third1 (
      .A(SecSig[0]),
      .B(CIn[6]),
      .C(CIn[5]),
      .Carry(COut[9]),
      .S(ThiSig[0])
  );
  ysyx_040656_mul_addr third2 (
      .A(SecSig[3]),
      .B(SecSig[2]),
      .C(SecSig[1]),
      .Carry(COut[10]),
      .S(ThiSig[1])
  );
  wire [1:0] ForSig;
  ysyx_040656_mul_addr fourth1 (
      .A(CIn[9]),
      .B(CIn[8]),
      .C(CIn[7]),
      .Carry(COut[11]),
      .S(ForSig[0])
  );
  ysyx_040656_mul_addr fourth2 (
      .A(ThiSig[1]),
      .B(ThiSig[0]),
      .C(CIn[10]),
      .Carry(COut[12]),
      .S(ForSig[1])
  );
  wire FifSig;
  ysyx_040656_mul_addr fifth1 (
      .A(ForSig[1]),
      .B(ForSig[0]),
      .C(CIn[11]),
      .Carry(COut[13]),
      .S(FifSig)
  );
  ysyx_040656_mul_addr sixth1 (
      .A(FifSig),
      .B(CIn[13]),
      .C(CIn[12]),
      .Carry(C),
      .S(S)
  );
endmodule
module ysyx_040656_mul_mul (
    input clock,
    input reset,
    input sign,
    input [31:0] x,
    input [31:0] y,
    output [63:0] result
);
  wire [63:0] CalX;
  wire [32:0] CalY;
  assign CalX = sign ? {{32{x[31]}}, x} : {32'b0, x};
  assign CalY = sign ? {y[31], y} : {1'b0, y};
  wire [16:0] Carry;
  wire [63:0] BoothRes[17];
  ysyx_040656_mul_BoothInterBase fir (
      .y({CalY[1], CalY[0], 1'b0}),
      .InX(CalX),
      .OutX(BoothRes[0]),
      .Carry(Carry[0])
  );
  generate
    genvar i;
    for (i = 2; i < 32; i = i + 2) begin : g_boothfor
      ysyx_040656_mul_BoothInterBase ai (
          .y(CalY[i+1:i-1]),
          .InX(CalX << i),
          .OutX(BoothRes[i>>1]),
          .Carry(Carry[i>>1])
      );
    end
  endgenerate
  ysyx_040656_mul_BoothInterBase las (
      .y({CalY[32], CalY[32], CalY[31]}),
      .InX(CalX << 32),
      .OutX(BoothRes[16]),
      .Carry(Carry[16])
  );
  reg [16:0] SecStageCarry;
  reg [63:0] SecStageBoothRes[17];
  integer p;
  always @(posedge clock) begin
    if (!reset) begin
      SecStageCarry <= Carry;
      for (p = 0; p < 17; p = p + 1) begin
        SecStageBoothRes[p] <= BoothRes[p];
      end
    end else begin
      SecStageCarry <= 0;
      for (p = 0; p < 17; p = p + 1) begin
        SecStageBoothRes[p] <= 0;
      end
    end
  end
  wire [13:0] WallaceInter[65]  /*verilator split_var*/;
  wire [63:0] COut, SOut;
  ysyx_040656_mul_WallaceTreeBase firs (
      .InData({
        SecStageBoothRes[0][0],
        SecStageBoothRes[1][0],
        SecStageBoothRes[2][0],
        SecStageBoothRes[3][0],
        SecStageBoothRes[4][0],
        SecStageBoothRes[5][0],
        SecStageBoothRes[6][0],
        SecStageBoothRes[7][0],
        SecStageBoothRes[8][0],
        SecStageBoothRes[9][0],
        SecStageBoothRes[10][0],
        SecStageBoothRes[11][0],
        SecStageBoothRes[12][0],
        SecStageBoothRes[13][0],
        SecStageBoothRes[14][0],
        SecStageBoothRes[15][0],
        SecStageBoothRes[16][0]
      }),
      .CIn(SecStageCarry[13:0]),
      .COut(WallaceInter[1]),
      .C(COut[0]),
      .S(SOut[0])
  );
  generate
    genvar n;
    for (n = 1; n < 64; n = n + 1) begin : g_wallacefor
      ysyx_040656_mul_WallaceTreeBase bi (
          .InData({
            SecStageBoothRes[0][n],
            SecStageBoothRes[1][n],
            SecStageBoothRes[2][n],
            SecStageBoothRes[3][n],
            SecStageBoothRes[4][n],
            SecStageBoothRes[5][n],
            SecStageBoothRes[6][n],
            SecStageBoothRes[7][n],
            SecStageBoothRes[8][n],
            SecStageBoothRes[9][n],
            SecStageBoothRes[10][n],
            SecStageBoothRes[11][n],
            SecStageBoothRes[12][n],
            SecStageBoothRes[13][n],
            SecStageBoothRes[14][n],
            SecStageBoothRes[15][n],
            SecStageBoothRes[16][n]
          }),
          .CIn(WallaceInter[n]),
          .COut(WallaceInter[n+1]),
          .C(COut[n]),
          .S(SOut[n])
      );
    end
  endgenerate
  assign result = SOut + {COut[62:0], SecStageCarry[14]} + {63'd0, SecStageCarry[15]};
endmodule
module ysyx_040656_div_div (
    input clock,
    input reset,
    input valid,
    input out_ready,
    input sign,
    input [63:0] x,
    input [63:0] y,
    output [63:0] s,
    output [63:0] r,
    output reg ready,
    output reg out_valid
);
  reg  [64:0] UnsignS;
  reg  [64:0] UnsignR;
  reg  [64:0] tmp_r;
  reg  [ 6:0] count;
  wire [64:0] tmp_d;
  wire [64:0] result_r;
  wire [64:0] UnsignX, UnsignY;
  reg        sign_buffer;
  reg        x_63_buffer;
  reg        y_63_buffer;
  wire       real_sign;
  wire       real_x_63;
  wire       real_y_63;
  reg [31:0] st_cur;
  assign UnsignX = {1'b0, (real_sign ? (x[63] ? (~x + 1) : x) : x)};
  assign UnsignY = {1'b0, (real_sign ? (y[63] ? (~y + 1) : y) : y)};
  localparam int IDLE = 0;
  localparam int RUN = 1;
  localparam int COMPLETE = 2;
  wire real_complete = st_cur == COMPLETE;
  assign real_sign = real_complete ? sign_buffer : sign;
  assign real_x_63 = real_complete ? x_63_buffer : x[63];
  assign real_y_63 = real_complete ? y_63_buffer : y[63];
  always @(posedge clock) begin
    if (reset) begin
      st_cur      <= IDLE;
      sign_buffer <= 0;
      x_63_buffer <= 0;
      y_63_buffer <= 0;
      count       <= 7'd64;
      tmp_r       <= 0;
      out_valid   <= 0;
    end else begin
      case (st_cur)
        IDLE: begin
          out_valid <= 0;
          ready     <= 1;
          if (valid) begin
            ready       <= 1'b0;
            sign_buffer <= sign;
            x_63_buffer <= x[63];
            y_63_buffer <= y[63];
            st_cur      <= RUN;
            count       <= 7'd64;
            tmp_r       <= 0;
          end else begin
            ready  <= 1'b1;
            st_cur <= IDLE;
          end
        end
        RUN: begin
          if (count == 7'h7f) begin
            st_cur <= COMPLETE;
            out_valid <= 1;
            UnsignR <= tmp_r;
          end else begin
            ready     <= 1'b0;
            out_valid <= 0;
            count     <= count - 7'd1;
            if (tmp_d[64]) begin
              UnsignS <= {UnsignS[63:0], 1'b0};
              tmp_r   <= result_r;
            end else begin
              UnsignS <= {UnsignS[63:0], 1'b1};
              tmp_r   <= tmp_d;
            end
          end
        end
        COMPLETE: begin
          out_valid <= 0;
          if (out_ready) begin
            st_cur <= IDLE;
          end else ready <= 1'b0;
        end
        default: st_cur <= IDLE;
      endcase
    end
  end
  assign result_r = {tmp_r[63:0], UnsignX[count]};
  assign tmp_d    = result_r - UnsignY;
  wire [64:0] TmpS, TmpR;
  assign TmpS = (real_sign ? ((real_x_63 == real_y_63) ? UnsignS : ~(UnsignS - 1)) : UnsignS);
  assign TmpR = (real_sign ? (real_x_63 ? ~(UnsignR - 1) : UnsignR) : UnsignR);
  assign s = TmpS[63:0];
  assign r = TmpR[63:0];
endmodule
module ysyx_040656_InstructionFetchUnit(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [31:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_inst,
  output [31:0] io_out_bits_pc,
  input         io_redirect_valid,
  input  [31:0] io_redirect_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif
  reg [31:0] pc;
  reg [31:0] lastPC;
  reg [4:0] need2Flush;
  reg [31:0] redirectTarget;
  wire [31:0] if_pc_plus4 = pc + 32'h4;
  wire [31:0] if_pc_next = io_redirect_valid ? io_redirect_target : if_pc_plus4;
  wire  _T = io_imem_req_ready & io_imem_req_valid;
  wire [4:0] _need2Flush_T_1 = need2Flush - 5'h1;
  wire [31:0] _GEN_0 = need2Flush == 5'h1 ? if_pc_next : pc;
  wire [31:0] _GEN_1 = need2Flush == 5'h1 ? pc : lastPC;
  wire [4:0] _GEN_4 = need2Flush != 5'h0 ? _need2Flush_T_1 : need2Flush;
  assign io_imem_req_valid = 1'h1;
  assign io_imem_req_bits_addr = pc;
  assign io_imem_resp_ready = io_out_ready;
  assign io_out_valid = io_imem_resp_valid & need2Flush == 5'h0;
  assign io_out_bits_inst = io_imem_resp_bits_rdata[31:0];
  assign io_out_bits_pc = lastPC;
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h30000000;
    end else if (_T) begin
      if (need2Flush == 5'h3) begin
        pc <= redirectTarget;
      end else if (need2Flush != 5'h0) begin
        pc <= _GEN_0;
      end else begin
        pc <= if_pc_next;
      end
    end
    if (reset) begin
      lastPC <= pc;
    end else if (_T) begin
      if (need2Flush == 5'h3) begin
        lastPC <= pc;
      end else if (need2Flush != 5'h0) begin
        lastPC <= _GEN_1;
      end else begin
        lastPC <= pc;
      end
    end
    if (reset) begin
      need2Flush <= 5'h0;
    end else if (io_redirect_valid) begin
      need2Flush <= 5'h3;
    end else if (_T) begin
      if (need2Flush == 5'h3) begin
        need2Flush <= _need2Flush_T_1;
      end else begin
        need2Flush <= _GEN_4;
      end
    end
    if (reset) begin
      redirectTarget <= 32'h0;
    end else if (io_redirect_valid) begin
      redirectTarget <= io_redirect_target;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  lastPC = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  need2Flush = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  redirectTarget = _RAND_3[31:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_DecodeStage(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_inst,
  input  [31:0] io_in_bits_pc,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_pc,
  output [31:0] io_out_bits_inst,
  output        io_out_bits_valid,
  output        io_out_bits_bubble,
  output [2:0]  io_out_bits_opcode_type,
  output [5:0]  io_out_bits_opcode_func,
  output [3:0]  io_out_bits_br_type,
  output        io_out_bits_rf_en,
  output [4:0]  io_out_bits_wb_addr,
  output [1:0]  io_out_bits_wb_stage,
  output [63:0] io_out_bits_op1_data,
  output [63:0] io_out_bits_op2_data,
  output [63:0] io_out_bits_rs1_data,
  output [63:0] io_out_bits_rs2_data,
  output [4:0]  io_regFile_rs1_addr,
  output [4:0]  io_regFile_rs2_addr,
  input  [63:0] io_regFile_rs1_data,
  input  [63:0] io_regFile_rs2_data,
  input         io_bypass_0_rf_wen,
  input  [4:0]  io_bypass_0_addr,
  input  [63:0] io_bypass_0_data,
  input         io_bypass_1_rf_wen,
  input  [4:0]  io_bypass_1_addr,
  input  [63:0] io_bypass_1_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif
  reg [4:0] last_use_rd;
  reg [31:0] decodeBuffer_inst;
  wire [31:0] _decodeInfo_T = decodeBuffer_inst & 32'h7f;
  wire  _decodeInfo_T_1 = 32'h17 == _decodeInfo_T;
  wire  _decodeInfo_T_3 = 32'h37 == _decodeInfo_T;
  wire [31:0] _decodeInfo_T_4 = decodeBuffer_inst & 32'h707f;
  wire  _decodeInfo_T_5 = 32'h2003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_7 = 32'h1003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_9 = 32'h3 == _decodeInfo_T_4;
  wire  _decodeInfo_T_11 = 32'h3003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_13 = 32'h6003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_15 = 32'h5003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_17 = 32'h4003 == _decodeInfo_T_4;
  wire  _decodeInfo_T_19 = 32'h2023 == _decodeInfo_T_4;
  wire  _decodeInfo_T_21 = 32'h1023 == _decodeInfo_T_4;
  wire  _decodeInfo_T_23 = 32'h23 == _decodeInfo_T_4;
  wire  _decodeInfo_T_25 = 32'h3023 == _decodeInfo_T_4;
  wire  _decodeInfo_T_27 = 32'h13 == _decodeInfo_T_4;
  wire  _decodeInfo_T_29 = 32'h7013 == _decodeInfo_T_4;
  wire  _decodeInfo_T_31 = 32'h6013 == _decodeInfo_T_4;
  wire  _decodeInfo_T_33 = 32'h4013 == _decodeInfo_T_4;
  wire [31:0] _decodeInfo_T_34 = decodeBuffer_inst & 32'hfe00707f;
  wire  _decodeInfo_T_35 = 32'h3033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_37 = 32'h2013 == _decodeInfo_T_4;
  wire  _decodeInfo_T_39 = 32'h3013 == _decodeInfo_T_4;
  wire [31:0] _decodeInfo_T_40 = decodeBuffer_inst & 32'hfc00707f;
  wire  _decodeInfo_T_41 = 32'h1013 == _decodeInfo_T_40;
  wire  _decodeInfo_T_43 = 32'h40005013 == _decodeInfo_T_40;
  wire  _decodeInfo_T_45 = 32'h5013 == _decodeInfo_T_40;
  wire  _decodeInfo_T_47 = 32'h33 == _decodeInfo_T_34;
  wire  _decodeInfo_T_49 = 32'h40000033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_51 = 32'h7033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_53 = 32'h6033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_55 = 32'h4033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_57 = 32'h2033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_59 = 32'h1033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_61 = 32'h40005033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_63 = 32'h5033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_65 = 32'h3b == _decodeInfo_T_34;
  wire  _decodeInfo_T_67 = 32'h4000003b == _decodeInfo_T_34;
  wire  _decodeInfo_T_69 = 32'h103b == _decodeInfo_T_34;
  wire  _decodeInfo_T_71 = 32'h503b == _decodeInfo_T_34;
  wire  _decodeInfo_T_73 = 32'h4000503b == _decodeInfo_T_34;
  wire  _decodeInfo_T_75 = 32'h1b == _decodeInfo_T_4;
  wire  _decodeInfo_T_77 = 32'h101b == _decodeInfo_T_34;
  wire  _decodeInfo_T_79 = 32'h501b == _decodeInfo_T_34;
  wire  _decodeInfo_T_81 = 32'h4000501b == _decodeInfo_T_34;
  wire  _decodeInfo_T_83 = 32'h6f == _decodeInfo_T;
  wire  _decodeInfo_T_85 = 32'h67 == _decodeInfo_T_4;
  wire  _decodeInfo_T_87 = 32'h63 == _decodeInfo_T_4;
  wire  _decodeInfo_T_89 = 32'h1063 == _decodeInfo_T_4;
  wire  _decodeInfo_T_91 = 32'h4063 == _decodeInfo_T_4;
  wire  _decodeInfo_T_93 = 32'h6063 == _decodeInfo_T_4;
  wire  _decodeInfo_T_95 = 32'h5063 == _decodeInfo_T_4;
  wire  _decodeInfo_T_97 = 32'h7063 == _decodeInfo_T_4;
  wire  _decodeInfo_T_99 = 32'h2000033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_101 = 32'h2001033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_103 = 32'h2003033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_105 = 32'h2002033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_107 = 32'h2004033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_109 = 32'h2005033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_111 = 32'h2007033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_113 = 32'h200003b == _decodeInfo_T_34;
  wire  _decodeInfo_T_115 = 32'h200603b == _decodeInfo_T_34;
  wire  _decodeInfo_T_117 = 32'h200703b == _decodeInfo_T_34;
  wire  _decodeInfo_T_119 = 32'h200403b == _decodeInfo_T_34;
  wire  _decodeInfo_T_121 = 32'h200503b == _decodeInfo_T_34;
  wire  _decodeInfo_T_135 = 32'h2006033 == _decodeInfo_T_34;
  wire  _decodeInfo_T_149 = 32'hf == _decodeInfo_T_4;
  wire  _decodeInfo_T_151 = 32'h100f == _decodeInfo_T_4;
  wire [31:0] _decodeInfo_T_152 = decodeBuffer_inst & 32'hfe007fff;
  wire  _decodeInfo_T_153 = 32'h12000073 == _decodeInfo_T_152;
  wire  _decodeInfo_T_155 = 32'h73 == decodeBuffer_inst;
  wire  _decodeInfo_T_157 = 32'h100073 == decodeBuffer_inst;
  wire  _decodeInfo_T_159 = 32'h30200073 == decodeBuffer_inst;
  wire  _decodeInfo_T_161 = 32'h7b200073 == decodeBuffer_inst;
  wire  _decodeInfo_T_163 = 32'h2073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_165 = 32'h1073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_167 = 32'h3073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_169 = 32'h5073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_171 = 32'h6073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_173 = 32'h7073 == _decodeInfo_T_4;
  wire  _decodeInfo_T_438 = _decodeInfo_T_161 ? 1'h0 : _decodeInfo_T_163 | (_decodeInfo_T_165 | (_decodeInfo_T_167 | (
    _decodeInfo_T_169 | (_decodeInfo_T_171 | _decodeInfo_T_173))));
  wire  _decodeInfo_T_439 = _decodeInfo_T_159 ? 1'h0 : _decodeInfo_T_438;
  wire  _decodeInfo_T_440 = _decodeInfo_T_157 ? 1'h0 : _decodeInfo_T_439;
  wire  _decodeInfo_T_441 = _decodeInfo_T_155 ? 1'h0 : _decodeInfo_T_440;
  wire  _decodeInfo_T_442 = _decodeInfo_T_153 ? 1'h0 : _decodeInfo_T_441;
  wire  _decodeInfo_T_443 = _decodeInfo_T_151 ? 1'h0 : _decodeInfo_T_442;
  wire  _decodeInfo_T_444 = _decodeInfo_T_149 ? 1'h0 : _decodeInfo_T_443;
  wire  _decodeInfo_T_474 = _decodeInfo_T_89 | (_decodeInfo_T_91 | (_decodeInfo_T_93 | (_decodeInfo_T_95 | (
    _decodeInfo_T_97 | (_decodeInfo_T_99 | (_decodeInfo_T_101 | (_decodeInfo_T_103 | (_decodeInfo_T_105 | (
    _decodeInfo_T_107 | (_decodeInfo_T_109 | (_decodeInfo_T_111 | (_decodeInfo_T_113 | (_decodeInfo_T_115 | (
    _decodeInfo_T_117 | (_decodeInfo_T_119 | (_decodeInfo_T_121 | (_decodeInfo_T_99 | (_decodeInfo_T_101 | (
    _decodeInfo_T_103 | (_decodeInfo_T_105 | (_decodeInfo_T_107 | (_decodeInfo_T_109 | (_decodeInfo_T_135 | (
    _decodeInfo_T_111 | (_decodeInfo_T_113 | (_decodeInfo_T_115 | (_decodeInfo_T_117 | (_decodeInfo_T_119 | (
    _decodeInfo_T_121 | _decodeInfo_T_444)))))))))))))))))))))))))))));
  wire  _decodeInfo_T_504 = _decodeInfo_T_29 | (_decodeInfo_T_31 | (_decodeInfo_T_33 | (_decodeInfo_T_35 | (
    _decodeInfo_T_37 | (_decodeInfo_T_39 | (_decodeInfo_T_41 | (_decodeInfo_T_43 | (_decodeInfo_T_45 | (_decodeInfo_T_47
     | (_decodeInfo_T_49 | (_decodeInfo_T_51 | (_decodeInfo_T_53 | (_decodeInfo_T_55 | (_decodeInfo_T_57 | (
    _decodeInfo_T_59 | (_decodeInfo_T_61 | (_decodeInfo_T_63 | (_decodeInfo_T_65 | (_decodeInfo_T_67 | (_decodeInfo_T_69
     | (_decodeInfo_T_71 | (_decodeInfo_T_73 | (_decodeInfo_T_75 | (_decodeInfo_T_77 | (_decodeInfo_T_79 | (
    _decodeInfo_T_81 | (_decodeInfo_T_83 | (_decodeInfo_T_85 | (_decodeInfo_T_87 | _decodeInfo_T_474))))))))))))))))))))
    )))))))));
  wire  decodeInfo_3 = _decodeInfo_T_1 | (_decodeInfo_T_3 | (_decodeInfo_T_5 | (_decodeInfo_T_7 | (_decodeInfo_T_9 | (
    _decodeInfo_T_11 | (_decodeInfo_T_13 | (_decodeInfo_T_15 | (_decodeInfo_T_17 | (_decodeInfo_T_19 | (_decodeInfo_T_21
     | (_decodeInfo_T_23 | (_decodeInfo_T_25 | (_decodeInfo_T_27 | _decodeInfo_T_504)))))))))))));
  wire [4:0] dec_rs_addr_0 = decodeBuffer_inst[19:15];
  wire [4:0] _needWait_T_2 = ~decodeInfo_3 ? 5'h0 : dec_rs_addr_0;
  wire  _decodeInfo_T_603 = _decodeInfo_T_3 ? 1'h0 : _decodeInfo_T_5 | (_decodeInfo_T_7 | (_decodeInfo_T_9 | (
    _decodeInfo_T_11 | (_decodeInfo_T_13 | (_decodeInfo_T_15 | (_decodeInfo_T_17 | (_decodeInfo_T_19 | (_decodeInfo_T_21
     | (_decodeInfo_T_23 | (_decodeInfo_T_25 | (_decodeInfo_T_27 | _decodeInfo_T_504)))))))))));
  wire  decodeInfo_4 = _decodeInfo_T_1 | _decodeInfo_T_603;
  wire [4:0] dec_rs_addr_1 = decodeBuffer_inst[24:20];
  wire [4:0] _needWait_T_5 = ~decodeInfo_4 ? 5'h0 : dec_rs_addr_1;
  wire  _needWait_T_6 = _needWait_T_5 == last_use_rd;
  wire  _needWait_T_7 = _needWait_T_2 == last_use_rd | _needWait_T_6;
  wire  needWait = last_use_rd != 5'h0 & _needWait_T_7;
  wire  _io_in_ready_T = ~needWait;
  reg [31:0] decodeBuffer_pc;
  reg  decodeBuffer_bubble;
  wire [2:0] _decodeInfo_T_212 = _decodeInfo_T_97 ? 3'h4 : 3'h0;
  wire [2:0] _decodeInfo_T_213 = _decodeInfo_T_95 ? 3'h3 : _decodeInfo_T_212;
  wire [2:0] _decodeInfo_T_214 = _decodeInfo_T_93 ? 3'h6 : _decodeInfo_T_213;
  wire [2:0] _decodeInfo_T_215 = _decodeInfo_T_91 ? 3'h5 : _decodeInfo_T_214;
  wire [2:0] _decodeInfo_T_216 = _decodeInfo_T_89 ? 3'h1 : _decodeInfo_T_215;
  wire [2:0] _decodeInfo_T_217 = _decodeInfo_T_87 ? 3'h2 : _decodeInfo_T_216;
  wire [3:0] _decodeInfo_T_218 = _decodeInfo_T_85 ? 4'h8 : {{1'd0}, _decodeInfo_T_217};
  wire [3:0] _decodeInfo_T_219 = _decodeInfo_T_83 ? 4'h7 : _decodeInfo_T_218;
  wire [3:0] _decodeInfo_T_220 = _decodeInfo_T_81 ? 4'h0 : _decodeInfo_T_219;
  wire [3:0] _decodeInfo_T_221 = _decodeInfo_T_79 ? 4'h0 : _decodeInfo_T_220;
  wire [3:0] _decodeInfo_T_222 = _decodeInfo_T_77 ? 4'h0 : _decodeInfo_T_221;
  wire [3:0] _decodeInfo_T_223 = _decodeInfo_T_75 ? 4'h0 : _decodeInfo_T_222;
  wire [3:0] _decodeInfo_T_224 = _decodeInfo_T_73 ? 4'h0 : _decodeInfo_T_223;
  wire [3:0] _decodeInfo_T_225 = _decodeInfo_T_71 ? 4'h0 : _decodeInfo_T_224;
  wire [3:0] _decodeInfo_T_226 = _decodeInfo_T_69 ? 4'h0 : _decodeInfo_T_225;
  wire [3:0] _decodeInfo_T_227 = _decodeInfo_T_67 ? 4'h0 : _decodeInfo_T_226;
  wire [3:0] _decodeInfo_T_228 = _decodeInfo_T_65 ? 4'h0 : _decodeInfo_T_227;
  wire [3:0] _decodeInfo_T_229 = _decodeInfo_T_63 ? 4'h0 : _decodeInfo_T_228;
  wire [3:0] _decodeInfo_T_230 = _decodeInfo_T_61 ? 4'h0 : _decodeInfo_T_229;
  wire [3:0] _decodeInfo_T_231 = _decodeInfo_T_59 ? 4'h0 : _decodeInfo_T_230;
  wire [3:0] _decodeInfo_T_232 = _decodeInfo_T_57 ? 4'h0 : _decodeInfo_T_231;
  wire [3:0] _decodeInfo_T_233 = _decodeInfo_T_55 ? 4'h0 : _decodeInfo_T_232;
  wire [3:0] _decodeInfo_T_234 = _decodeInfo_T_53 ? 4'h0 : _decodeInfo_T_233;
  wire [3:0] _decodeInfo_T_235 = _decodeInfo_T_51 ? 4'h0 : _decodeInfo_T_234;
  wire [3:0] _decodeInfo_T_236 = _decodeInfo_T_49 ? 4'h0 : _decodeInfo_T_235;
  wire [3:0] _decodeInfo_T_237 = _decodeInfo_T_47 ? 4'h0 : _decodeInfo_T_236;
  wire [3:0] _decodeInfo_T_238 = _decodeInfo_T_45 ? 4'h0 : _decodeInfo_T_237;
  wire [3:0] _decodeInfo_T_239 = _decodeInfo_T_43 ? 4'h0 : _decodeInfo_T_238;
  wire [3:0] _decodeInfo_T_240 = _decodeInfo_T_41 ? 4'h0 : _decodeInfo_T_239;
  wire [3:0] _decodeInfo_T_241 = _decodeInfo_T_39 ? 4'h0 : _decodeInfo_T_240;
  wire [3:0] _decodeInfo_T_242 = _decodeInfo_T_37 ? 4'h0 : _decodeInfo_T_241;
  wire [3:0] _decodeInfo_T_243 = _decodeInfo_T_35 ? 4'h0 : _decodeInfo_T_242;
  wire [3:0] _decodeInfo_T_244 = _decodeInfo_T_33 ? 4'h0 : _decodeInfo_T_243;
  wire [3:0] _decodeInfo_T_245 = _decodeInfo_T_31 ? 4'h0 : _decodeInfo_T_244;
  wire [3:0] _decodeInfo_T_246 = _decodeInfo_T_29 ? 4'h0 : _decodeInfo_T_245;
  wire [3:0] _decodeInfo_T_247 = _decodeInfo_T_27 ? 4'h0 : _decodeInfo_T_246;
  wire [3:0] _decodeInfo_T_248 = _decodeInfo_T_25 ? 4'h0 : _decodeInfo_T_247;
  wire [3:0] _decodeInfo_T_249 = _decodeInfo_T_23 ? 4'h0 : _decodeInfo_T_248;
  wire [3:0] _decodeInfo_T_250 = _decodeInfo_T_21 ? 4'h0 : _decodeInfo_T_249;
  wire [3:0] _decodeInfo_T_251 = _decodeInfo_T_19 ? 4'h0 : _decodeInfo_T_250;
  wire [3:0] _decodeInfo_T_252 = _decodeInfo_T_17 ? 4'h0 : _decodeInfo_T_251;
  wire [3:0] _decodeInfo_T_253 = _decodeInfo_T_15 ? 4'h0 : _decodeInfo_T_252;
  wire [3:0] _decodeInfo_T_254 = _decodeInfo_T_13 ? 4'h0 : _decodeInfo_T_253;
  wire [3:0] _decodeInfo_T_255 = _decodeInfo_T_11 ? 4'h0 : _decodeInfo_T_254;
  wire [3:0] _decodeInfo_T_256 = _decodeInfo_T_9 ? 4'h0 : _decodeInfo_T_255;
  wire [3:0] _decodeInfo_T_257 = _decodeInfo_T_7 ? 4'h0 : _decodeInfo_T_256;
  wire [3:0] _decodeInfo_T_258 = _decodeInfo_T_5 ? 4'h0 : _decodeInfo_T_257;
  wire [3:0] _decodeInfo_T_259 = _decodeInfo_T_3 ? 4'h0 : _decodeInfo_T_258;
  wire [2:0] _decodeInfo_T_260 = _decodeInfo_T_173 ? 3'h5 : 3'h0;
  wire [2:0] _decodeInfo_T_261 = _decodeInfo_T_171 ? 3'h5 : _decodeInfo_T_260;
  wire [2:0] _decodeInfo_T_262 = _decodeInfo_T_169 ? 3'h5 : _decodeInfo_T_261;
  wire [2:0] _decodeInfo_T_263 = _decodeInfo_T_167 ? 3'h2 : _decodeInfo_T_262;
  wire [2:0] _decodeInfo_T_264 = _decodeInfo_T_165 ? 3'h2 : _decodeInfo_T_263;
  wire [2:0] _decodeInfo_T_265 = _decodeInfo_T_163 ? 3'h2 : _decodeInfo_T_264;
  wire [2:0] _decodeInfo_T_266 = _decodeInfo_T_161 ? 3'h0 : _decodeInfo_T_265;
  wire [2:0] _decodeInfo_T_267 = _decodeInfo_T_159 ? 3'h0 : _decodeInfo_T_266;
  wire [2:0] _decodeInfo_T_268 = _decodeInfo_T_157 ? 3'h0 : _decodeInfo_T_267;
  wire [2:0] _decodeInfo_T_269 = _decodeInfo_T_155 ? 3'h0 : _decodeInfo_T_268;
  wire [2:0] _decodeInfo_T_270 = _decodeInfo_T_153 ? 3'h0 : _decodeInfo_T_269;
  wire [2:0] _decodeInfo_T_271 = _decodeInfo_T_151 ? 3'h0 : _decodeInfo_T_270;
  wire [2:0] _decodeInfo_T_272 = _decodeInfo_T_149 ? 3'h0 : _decodeInfo_T_271;
  wire [2:0] _decodeInfo_T_273 = _decodeInfo_T_121 ? 3'h2 : _decodeInfo_T_272;
  wire [2:0] _decodeInfo_T_274 = _decodeInfo_T_119 ? 3'h2 : _decodeInfo_T_273;
  wire [2:0] _decodeInfo_T_275 = _decodeInfo_T_117 ? 3'h2 : _decodeInfo_T_274;
  wire [2:0] _decodeInfo_T_276 = _decodeInfo_T_115 ? 3'h2 : _decodeInfo_T_275;
  wire [2:0] _decodeInfo_T_277 = _decodeInfo_T_113 ? 3'h2 : _decodeInfo_T_276;
  wire [2:0] _decodeInfo_T_278 = _decodeInfo_T_111 ? 3'h2 : _decodeInfo_T_277;
  wire [2:0] _decodeInfo_T_279 = _decodeInfo_T_135 ? 3'h2 : _decodeInfo_T_278;
  wire [2:0] _decodeInfo_T_280 = _decodeInfo_T_109 ? 3'h2 : _decodeInfo_T_279;
  wire [2:0] _decodeInfo_T_281 = _decodeInfo_T_107 ? 3'h2 : _decodeInfo_T_280;
  wire [2:0] _decodeInfo_T_282 = _decodeInfo_T_105 ? 3'h2 : _decodeInfo_T_281;
  wire [2:0] _decodeInfo_T_283 = _decodeInfo_T_103 ? 3'h2 : _decodeInfo_T_282;
  wire [2:0] _decodeInfo_T_284 = _decodeInfo_T_101 ? 3'h2 : _decodeInfo_T_283;
  wire [2:0] _decodeInfo_T_285 = _decodeInfo_T_99 ? 3'h2 : _decodeInfo_T_284;
  wire [2:0] _decodeInfo_T_286 = _decodeInfo_T_121 ? 3'h2 : _decodeInfo_T_285;
  wire [2:0] _decodeInfo_T_287 = _decodeInfo_T_119 ? 3'h2 : _decodeInfo_T_286;
  wire [2:0] _decodeInfo_T_288 = _decodeInfo_T_117 ? 3'h2 : _decodeInfo_T_287;
  wire [2:0] _decodeInfo_T_289 = _decodeInfo_T_115 ? 3'h2 : _decodeInfo_T_288;
  wire [2:0] _decodeInfo_T_290 = _decodeInfo_T_113 ? 3'h2 : _decodeInfo_T_289;
  wire [2:0] _decodeInfo_T_291 = _decodeInfo_T_111 ? 3'h2 : _decodeInfo_T_290;
  wire [2:0] _decodeInfo_T_292 = _decodeInfo_T_109 ? 3'h2 : _decodeInfo_T_291;
  wire [2:0] _decodeInfo_T_293 = _decodeInfo_T_107 ? 3'h2 : _decodeInfo_T_292;
  wire [2:0] _decodeInfo_T_294 = _decodeInfo_T_105 ? 3'h2 : _decodeInfo_T_293;
  wire [2:0] _decodeInfo_T_295 = _decodeInfo_T_103 ? 3'h2 : _decodeInfo_T_294;
  wire [2:0] _decodeInfo_T_296 = _decodeInfo_T_101 ? 3'h2 : _decodeInfo_T_295;
  wire [2:0] _decodeInfo_T_297 = _decodeInfo_T_99 ? 3'h2 : _decodeInfo_T_296;
  wire [2:0] _decodeInfo_T_298 = _decodeInfo_T_97 ? 3'h7 : _decodeInfo_T_297;
  wire [2:0] _decodeInfo_T_299 = _decodeInfo_T_95 ? 3'h7 : _decodeInfo_T_298;
  wire [2:0] _decodeInfo_T_300 = _decodeInfo_T_93 ? 3'h7 : _decodeInfo_T_299;
  wire [2:0] _decodeInfo_T_301 = _decodeInfo_T_91 ? 3'h7 : _decodeInfo_T_300;
  wire [2:0] _decodeInfo_T_302 = _decodeInfo_T_89 ? 3'h7 : _decodeInfo_T_301;
  wire [2:0] _decodeInfo_T_303 = _decodeInfo_T_87 ? 3'h7 : _decodeInfo_T_302;
  wire [2:0] _decodeInfo_T_304 = _decodeInfo_T_85 ? 3'h2 : _decodeInfo_T_303;
  wire [2:0] _decodeInfo_T_305 = _decodeInfo_T_83 ? 3'h3 : _decodeInfo_T_304;
  wire [2:0] _decodeInfo_T_306 = _decodeInfo_T_81 ? 3'h2 : _decodeInfo_T_305;
  wire [2:0] _decodeInfo_T_307 = _decodeInfo_T_79 ? 3'h2 : _decodeInfo_T_306;
  wire [2:0] _decodeInfo_T_308 = _decodeInfo_T_77 ? 3'h2 : _decodeInfo_T_307;
  wire [2:0] _decodeInfo_T_309 = _decodeInfo_T_75 ? 3'h2 : _decodeInfo_T_308;
  wire [2:0] _decodeInfo_T_310 = _decodeInfo_T_73 ? 3'h2 : _decodeInfo_T_309;
  wire [2:0] _decodeInfo_T_311 = _decodeInfo_T_71 ? 3'h2 : _decodeInfo_T_310;
  wire [2:0] _decodeInfo_T_312 = _decodeInfo_T_69 ? 3'h2 : _decodeInfo_T_311;
  wire [2:0] _decodeInfo_T_313 = _decodeInfo_T_67 ? 3'h2 : _decodeInfo_T_312;
  wire [2:0] _decodeInfo_T_314 = _decodeInfo_T_65 ? 3'h2 : _decodeInfo_T_313;
  wire [2:0] _decodeInfo_T_315 = _decodeInfo_T_63 ? 3'h2 : _decodeInfo_T_314;
  wire [2:0] _decodeInfo_T_316 = _decodeInfo_T_61 ? 3'h2 : _decodeInfo_T_315;
  wire [2:0] _decodeInfo_T_317 = _decodeInfo_T_59 ? 3'h2 : _decodeInfo_T_316;
  wire [2:0] _decodeInfo_T_318 = _decodeInfo_T_57 ? 3'h2 : _decodeInfo_T_317;
  wire [2:0] _decodeInfo_T_319 = _decodeInfo_T_55 ? 3'h2 : _decodeInfo_T_318;
  wire [2:0] _decodeInfo_T_320 = _decodeInfo_T_53 ? 3'h2 : _decodeInfo_T_319;
  wire [2:0] _decodeInfo_T_321 = _decodeInfo_T_51 ? 3'h2 : _decodeInfo_T_320;
  wire [2:0] _decodeInfo_T_322 = _decodeInfo_T_49 ? 3'h2 : _decodeInfo_T_321;
  wire [2:0] _decodeInfo_T_323 = _decodeInfo_T_47 ? 3'h2 : _decodeInfo_T_322;
  wire [2:0] _decodeInfo_T_324 = _decodeInfo_T_45 ? 3'h2 : _decodeInfo_T_323;
  wire [2:0] _decodeInfo_T_325 = _decodeInfo_T_43 ? 3'h2 : _decodeInfo_T_324;
  wire [2:0] _decodeInfo_T_326 = _decodeInfo_T_41 ? 3'h2 : _decodeInfo_T_325;
  wire [2:0] _decodeInfo_T_327 = _decodeInfo_T_39 ? 3'h2 : _decodeInfo_T_326;
  wire [2:0] _decodeInfo_T_328 = _decodeInfo_T_37 ? 3'h2 : _decodeInfo_T_327;
  wire [2:0] _decodeInfo_T_329 = _decodeInfo_T_35 ? 3'h2 : _decodeInfo_T_328;
  wire [2:0] _decodeInfo_T_330 = _decodeInfo_T_33 ? 3'h2 : _decodeInfo_T_329;
  wire [2:0] _decodeInfo_T_331 = _decodeInfo_T_31 ? 3'h2 : _decodeInfo_T_330;
  wire [2:0] _decodeInfo_T_332 = _decodeInfo_T_29 ? 3'h2 : _decodeInfo_T_331;
  wire [2:0] _decodeInfo_T_333 = _decodeInfo_T_27 ? 3'h2 : _decodeInfo_T_332;
  wire [2:0] _decodeInfo_T_334 = _decodeInfo_T_25 ? 3'h2 : _decodeInfo_T_333;
  wire [2:0] _decodeInfo_T_335 = _decodeInfo_T_23 ? 3'h2 : _decodeInfo_T_334;
  wire [2:0] _decodeInfo_T_336 = _decodeInfo_T_21 ? 3'h2 : _decodeInfo_T_335;
  wire [2:0] _decodeInfo_T_337 = _decodeInfo_T_19 ? 3'h2 : _decodeInfo_T_336;
  wire [2:0] _decodeInfo_T_338 = _decodeInfo_T_17 ? 3'h2 : _decodeInfo_T_337;
  wire [2:0] _decodeInfo_T_339 = _decodeInfo_T_15 ? 3'h2 : _decodeInfo_T_338;
  wire [2:0] _decodeInfo_T_340 = _decodeInfo_T_13 ? 3'h2 : _decodeInfo_T_339;
  wire [2:0] _decodeInfo_T_341 = _decodeInfo_T_11 ? 3'h2 : _decodeInfo_T_340;
  wire [2:0] _decodeInfo_T_342 = _decodeInfo_T_9 ? 3'h2 : _decodeInfo_T_341;
  wire [2:0] _decodeInfo_T_343 = _decodeInfo_T_7 ? 3'h2 : _decodeInfo_T_342;
  wire [2:0] _decodeInfo_T_344 = _decodeInfo_T_5 ? 3'h2 : _decodeInfo_T_343;
  wire [2:0] _decodeInfo_T_345 = _decodeInfo_T_3 ? 3'h1 : _decodeInfo_T_344;
  wire [2:0] decodeInfo_1 = _decodeInfo_T_1 ? 3'h1 : _decodeInfo_T_345;
  wire [2:0] _decodeInfo_T_359 = _decodeInfo_T_121 ? 3'h6 : 3'h0;
  wire [2:0] _decodeInfo_T_360 = _decodeInfo_T_119 ? 3'h6 : _decodeInfo_T_359;
  wire [2:0] _decodeInfo_T_361 = _decodeInfo_T_117 ? 3'h6 : _decodeInfo_T_360;
  wire [2:0] _decodeInfo_T_362 = _decodeInfo_T_115 ? 3'h6 : _decodeInfo_T_361;
  wire [2:0] _decodeInfo_T_363 = _decodeInfo_T_113 ? 3'h6 : _decodeInfo_T_362;
  wire [2:0] _decodeInfo_T_364 = _decodeInfo_T_111 ? 3'h6 : _decodeInfo_T_363;
  wire [2:0] _decodeInfo_T_365 = _decodeInfo_T_135 ? 3'h6 : _decodeInfo_T_364;
  wire [2:0] _decodeInfo_T_366 = _decodeInfo_T_109 ? 3'h6 : _decodeInfo_T_365;
  wire [2:0] _decodeInfo_T_367 = _decodeInfo_T_107 ? 3'h6 : _decodeInfo_T_366;
  wire [2:0] _decodeInfo_T_368 = _decodeInfo_T_105 ? 3'h6 : _decodeInfo_T_367;
  wire [2:0] _decodeInfo_T_369 = _decodeInfo_T_103 ? 3'h6 : _decodeInfo_T_368;
  wire [2:0] _decodeInfo_T_370 = _decodeInfo_T_101 ? 3'h6 : _decodeInfo_T_369;
  wire [2:0] _decodeInfo_T_371 = _decodeInfo_T_99 ? 3'h6 : _decodeInfo_T_370;
  wire [2:0] _decodeInfo_T_372 = _decodeInfo_T_121 ? 3'h6 : _decodeInfo_T_371;
  wire [2:0] _decodeInfo_T_373 = _decodeInfo_T_119 ? 3'h6 : _decodeInfo_T_372;
  wire [2:0] _decodeInfo_T_374 = _decodeInfo_T_117 ? 3'h6 : _decodeInfo_T_373;
  wire [2:0] _decodeInfo_T_375 = _decodeInfo_T_115 ? 3'h6 : _decodeInfo_T_374;
  wire [2:0] _decodeInfo_T_376 = _decodeInfo_T_113 ? 3'h6 : _decodeInfo_T_375;
  wire [2:0] _decodeInfo_T_377 = _decodeInfo_T_111 ? 3'h6 : _decodeInfo_T_376;
  wire [2:0] _decodeInfo_T_378 = _decodeInfo_T_109 ? 3'h6 : _decodeInfo_T_377;
  wire [2:0] _decodeInfo_T_379 = _decodeInfo_T_107 ? 3'h6 : _decodeInfo_T_378;
  wire [2:0] _decodeInfo_T_380 = _decodeInfo_T_105 ? 3'h6 : _decodeInfo_T_379;
  wire [2:0] _decodeInfo_T_381 = _decodeInfo_T_103 ? 3'h6 : _decodeInfo_T_380;
  wire [2:0] _decodeInfo_T_382 = _decodeInfo_T_101 ? 3'h6 : _decodeInfo_T_381;
  wire [2:0] _decodeInfo_T_383 = _decodeInfo_T_99 ? 3'h6 : _decodeInfo_T_382;
  wire [3:0] _decodeInfo_T_384 = _decodeInfo_T_97 ? 4'h9 : {{1'd0}, _decodeInfo_T_383};
  wire [3:0] _decodeInfo_T_385 = _decodeInfo_T_95 ? 4'h9 : _decodeInfo_T_384;
  wire [3:0] _decodeInfo_T_386 = _decodeInfo_T_93 ? 4'h9 : _decodeInfo_T_385;
  wire [3:0] _decodeInfo_T_387 = _decodeInfo_T_91 ? 4'h9 : _decodeInfo_T_386;
  wire [3:0] _decodeInfo_T_388 = _decodeInfo_T_89 ? 4'h9 : _decodeInfo_T_387;
  wire [3:0] _decodeInfo_T_389 = _decodeInfo_T_87 ? 4'h9 : _decodeInfo_T_388;
  wire [3:0] _decodeInfo_T_390 = _decodeInfo_T_85 ? 4'h4 : _decodeInfo_T_389;
  wire [3:0] _decodeInfo_T_391 = _decodeInfo_T_83 ? 4'h7 : _decodeInfo_T_390;
  wire [3:0] _decodeInfo_T_392 = _decodeInfo_T_81 ? 4'h4 : _decodeInfo_T_391;
  wire [3:0] _decodeInfo_T_393 = _decodeInfo_T_79 ? 4'h4 : _decodeInfo_T_392;
  wire [3:0] _decodeInfo_T_394 = _decodeInfo_T_77 ? 4'h4 : _decodeInfo_T_393;
  wire [3:0] _decodeInfo_T_395 = _decodeInfo_T_75 ? 4'h4 : _decodeInfo_T_394;
  wire [3:0] _decodeInfo_T_396 = _decodeInfo_T_73 ? 4'h6 : _decodeInfo_T_395;
  wire [3:0] _decodeInfo_T_397 = _decodeInfo_T_71 ? 4'h6 : _decodeInfo_T_396;
  wire [3:0] _decodeInfo_T_398 = _decodeInfo_T_69 ? 4'h6 : _decodeInfo_T_397;
  wire [3:0] _decodeInfo_T_399 = _decodeInfo_T_67 ? 4'h6 : _decodeInfo_T_398;
  wire [3:0] _decodeInfo_T_400 = _decodeInfo_T_65 ? 4'h6 : _decodeInfo_T_399;
  wire [3:0] _decodeInfo_T_401 = _decodeInfo_T_63 ? 4'h6 : _decodeInfo_T_400;
  wire [3:0] _decodeInfo_T_402 = _decodeInfo_T_61 ? 4'h6 : _decodeInfo_T_401;
  wire [3:0] _decodeInfo_T_403 = _decodeInfo_T_59 ? 4'h6 : _decodeInfo_T_402;
  wire [3:0] _decodeInfo_T_404 = _decodeInfo_T_57 ? 4'h6 : _decodeInfo_T_403;
  wire [3:0] _decodeInfo_T_405 = _decodeInfo_T_55 ? 4'h6 : _decodeInfo_T_404;
  wire [3:0] _decodeInfo_T_406 = _decodeInfo_T_53 ? 4'h6 : _decodeInfo_T_405;
  wire [3:0] _decodeInfo_T_407 = _decodeInfo_T_51 ? 4'h6 : _decodeInfo_T_406;
  wire [3:0] _decodeInfo_T_408 = _decodeInfo_T_49 ? 4'h6 : _decodeInfo_T_407;
  wire [3:0] _decodeInfo_T_409 = _decodeInfo_T_47 ? 4'h6 : _decodeInfo_T_408;
  wire [3:0] _decodeInfo_T_410 = _decodeInfo_T_45 ? 4'h4 : _decodeInfo_T_409;
  wire [3:0] _decodeInfo_T_411 = _decodeInfo_T_43 ? 4'h4 : _decodeInfo_T_410;
  wire [3:0] _decodeInfo_T_412 = _decodeInfo_T_41 ? 4'h4 : _decodeInfo_T_411;
  wire [3:0] _decodeInfo_T_413 = _decodeInfo_T_39 ? 4'h4 : _decodeInfo_T_412;
  wire [3:0] _decodeInfo_T_414 = _decodeInfo_T_37 ? 4'h4 : _decodeInfo_T_413;
  wire [3:0] _decodeInfo_T_415 = _decodeInfo_T_35 ? 4'h6 : _decodeInfo_T_414;
  wire [3:0] _decodeInfo_T_416 = _decodeInfo_T_33 ? 4'h4 : _decodeInfo_T_415;
  wire [3:0] _decodeInfo_T_417 = _decodeInfo_T_31 ? 4'h4 : _decodeInfo_T_416;
  wire [3:0] _decodeInfo_T_418 = _decodeInfo_T_29 ? 4'h4 : _decodeInfo_T_417;
  wire [3:0] _decodeInfo_T_419 = _decodeInfo_T_27 ? 4'h4 : _decodeInfo_T_418;
  wire [3:0] _decodeInfo_T_420 = _decodeInfo_T_25 ? 4'h8 : _decodeInfo_T_419;
  wire [3:0] _decodeInfo_T_421 = _decodeInfo_T_23 ? 4'h8 : _decodeInfo_T_420;
  wire [3:0] _decodeInfo_T_422 = _decodeInfo_T_21 ? 4'h8 : _decodeInfo_T_421;
  wire [3:0] _decodeInfo_T_423 = _decodeInfo_T_19 ? 4'h8 : _decodeInfo_T_422;
  wire [3:0] _decodeInfo_T_424 = _decodeInfo_T_17 ? 4'h4 : _decodeInfo_T_423;
  wire [3:0] _decodeInfo_T_425 = _decodeInfo_T_15 ? 4'h4 : _decodeInfo_T_424;
  wire [3:0] _decodeInfo_T_426 = _decodeInfo_T_13 ? 4'h4 : _decodeInfo_T_425;
  wire [3:0] _decodeInfo_T_427 = _decodeInfo_T_11 ? 4'h4 : _decodeInfo_T_426;
  wire [3:0] _decodeInfo_T_428 = _decodeInfo_T_9 ? 4'h4 : _decodeInfo_T_427;
  wire [3:0] _decodeInfo_T_429 = _decodeInfo_T_7 ? 4'h4 : _decodeInfo_T_428;
  wire [3:0] _decodeInfo_T_430 = _decodeInfo_T_5 ? 4'h4 : _decodeInfo_T_429;
  wire [3:0] _decodeInfo_T_431 = _decodeInfo_T_3 ? 4'h0 : _decodeInfo_T_430;
  wire [3:0] decodeInfo_2 = _decodeInfo_T_1 ? 4'h7 : _decodeInfo_T_431;
  wire [1:0] _decodeInfo_T_604 = _decodeInfo_T_173 ? 2'h3 : 2'h0;
  wire [1:0] _decodeInfo_T_605 = _decodeInfo_T_171 ? 2'h3 : _decodeInfo_T_604;
  wire [1:0] _decodeInfo_T_606 = _decodeInfo_T_169 ? 2'h3 : _decodeInfo_T_605;
  wire [1:0] _decodeInfo_T_607 = _decodeInfo_T_167 ? 2'h3 : _decodeInfo_T_606;
  wire [1:0] _decodeInfo_T_608 = _decodeInfo_T_165 ? 2'h3 : _decodeInfo_T_607;
  wire [1:0] _decodeInfo_T_609 = _decodeInfo_T_163 ? 2'h3 : _decodeInfo_T_608;
  wire [1:0] _decodeInfo_T_610 = _decodeInfo_T_161 ? 2'h3 : _decodeInfo_T_609;
  wire [1:0] _decodeInfo_T_611 = _decodeInfo_T_159 ? 2'h3 : _decodeInfo_T_610;
  wire [1:0] _decodeInfo_T_612 = _decodeInfo_T_157 ? 2'h3 : _decodeInfo_T_611;
  wire [1:0] _decodeInfo_T_613 = _decodeInfo_T_155 ? 2'h3 : _decodeInfo_T_612;
  wire [1:0] _decodeInfo_T_614 = _decodeInfo_T_153 ? 2'h3 : _decodeInfo_T_613;
  wire [2:0] _decodeInfo_T_615 = _decodeInfo_T_151 ? 3'h4 : {{1'd0}, _decodeInfo_T_614};
  wire [2:0] _decodeInfo_T_616 = _decodeInfo_T_149 ? 3'h4 : _decodeInfo_T_615;
  wire [2:0] _decodeInfo_T_617 = _decodeInfo_T_121 ? 3'h5 : _decodeInfo_T_616;
  wire [2:0] _decodeInfo_T_618 = _decodeInfo_T_119 ? 3'h5 : _decodeInfo_T_617;
  wire [2:0] _decodeInfo_T_619 = _decodeInfo_T_117 ? 3'h5 : _decodeInfo_T_618;
  wire [2:0] _decodeInfo_T_620 = _decodeInfo_T_115 ? 3'h5 : _decodeInfo_T_619;
  wire [2:0] _decodeInfo_T_621 = _decodeInfo_T_113 ? 3'h5 : _decodeInfo_T_620;
  wire [2:0] _decodeInfo_T_622 = _decodeInfo_T_111 ? 3'h5 : _decodeInfo_T_621;
  wire [2:0] _decodeInfo_T_623 = _decodeInfo_T_135 ? 3'h5 : _decodeInfo_T_622;
  wire [2:0] _decodeInfo_T_624 = _decodeInfo_T_109 ? 3'h5 : _decodeInfo_T_623;
  wire [2:0] _decodeInfo_T_625 = _decodeInfo_T_107 ? 3'h5 : _decodeInfo_T_624;
  wire [2:0] _decodeInfo_T_626 = _decodeInfo_T_105 ? 3'h5 : _decodeInfo_T_625;
  wire [2:0] _decodeInfo_T_627 = _decodeInfo_T_103 ? 3'h5 : _decodeInfo_T_626;
  wire [2:0] _decodeInfo_T_628 = _decodeInfo_T_101 ? 3'h5 : _decodeInfo_T_627;
  wire [2:0] _decodeInfo_T_629 = _decodeInfo_T_99 ? 3'h5 : _decodeInfo_T_628;
  wire [2:0] _decodeInfo_T_630 = _decodeInfo_T_121 ? 3'h5 : _decodeInfo_T_629;
  wire [2:0] _decodeInfo_T_631 = _decodeInfo_T_119 ? 3'h5 : _decodeInfo_T_630;
  wire [2:0] _decodeInfo_T_632 = _decodeInfo_T_117 ? 3'h5 : _decodeInfo_T_631;
  wire [2:0] _decodeInfo_T_633 = _decodeInfo_T_115 ? 3'h5 : _decodeInfo_T_632;
  wire [2:0] _decodeInfo_T_634 = _decodeInfo_T_113 ? 3'h5 : _decodeInfo_T_633;
  wire [2:0] _decodeInfo_T_635 = _decodeInfo_T_111 ? 3'h5 : _decodeInfo_T_634;
  wire [2:0] _decodeInfo_T_636 = _decodeInfo_T_109 ? 3'h5 : _decodeInfo_T_635;
  wire [2:0] _decodeInfo_T_637 = _decodeInfo_T_107 ? 3'h5 : _decodeInfo_T_636;
  wire [2:0] _decodeInfo_T_638 = _decodeInfo_T_105 ? 3'h5 : _decodeInfo_T_637;
  wire [2:0] _decodeInfo_T_639 = _decodeInfo_T_103 ? 3'h5 : _decodeInfo_T_638;
  wire [2:0] _decodeInfo_T_640 = _decodeInfo_T_101 ? 3'h5 : _decodeInfo_T_639;
  wire [2:0] _decodeInfo_T_641 = _decodeInfo_T_99 ? 3'h5 : _decodeInfo_T_640;
  wire [2:0] _decodeInfo_T_642 = _decodeInfo_T_97 ? 3'h6 : _decodeInfo_T_641;
  wire [2:0] _decodeInfo_T_643 = _decodeInfo_T_95 ? 3'h6 : _decodeInfo_T_642;
  wire [2:0] _decodeInfo_T_644 = _decodeInfo_T_93 ? 3'h6 : _decodeInfo_T_643;
  wire [2:0] _decodeInfo_T_645 = _decodeInfo_T_91 ? 3'h6 : _decodeInfo_T_644;
  wire [2:0] _decodeInfo_T_646 = _decodeInfo_T_89 ? 3'h6 : _decodeInfo_T_645;
  wire [2:0] _decodeInfo_T_647 = _decodeInfo_T_87 ? 3'h6 : _decodeInfo_T_646;
  wire [2:0] _decodeInfo_T_648 = _decodeInfo_T_85 ? 3'h6 : _decodeInfo_T_647;
  wire [2:0] _decodeInfo_T_649 = _decodeInfo_T_83 ? 3'h6 : _decodeInfo_T_648;
  wire [2:0] _decodeInfo_T_650 = _decodeInfo_T_81 ? 3'h1 : _decodeInfo_T_649;
  wire [2:0] _decodeInfo_T_651 = _decodeInfo_T_79 ? 3'h1 : _decodeInfo_T_650;
  wire [2:0] _decodeInfo_T_652 = _decodeInfo_T_77 ? 3'h1 : _decodeInfo_T_651;
  wire [2:0] _decodeInfo_T_653 = _decodeInfo_T_75 ? 3'h1 : _decodeInfo_T_652;
  wire [2:0] _decodeInfo_T_654 = _decodeInfo_T_73 ? 3'h1 : _decodeInfo_T_653;
  wire [2:0] _decodeInfo_T_655 = _decodeInfo_T_71 ? 3'h1 : _decodeInfo_T_654;
  wire [2:0] _decodeInfo_T_656 = _decodeInfo_T_69 ? 3'h1 : _decodeInfo_T_655;
  wire [2:0] _decodeInfo_T_657 = _decodeInfo_T_67 ? 3'h1 : _decodeInfo_T_656;
  wire [2:0] _decodeInfo_T_658 = _decodeInfo_T_65 ? 3'h1 : _decodeInfo_T_657;
  wire [2:0] _decodeInfo_T_659 = _decodeInfo_T_63 ? 3'h1 : _decodeInfo_T_658;
  wire [2:0] _decodeInfo_T_660 = _decodeInfo_T_61 ? 3'h1 : _decodeInfo_T_659;
  wire [2:0] _decodeInfo_T_661 = _decodeInfo_T_59 ? 3'h1 : _decodeInfo_T_660;
  wire [2:0] _decodeInfo_T_662 = _decodeInfo_T_57 ? 3'h1 : _decodeInfo_T_661;
  wire [2:0] _decodeInfo_T_663 = _decodeInfo_T_55 ? 3'h1 : _decodeInfo_T_662;
  wire [2:0] _decodeInfo_T_664 = _decodeInfo_T_53 ? 3'h1 : _decodeInfo_T_663;
  wire [2:0] _decodeInfo_T_665 = _decodeInfo_T_51 ? 3'h1 : _decodeInfo_T_664;
  wire [2:0] _decodeInfo_T_666 = _decodeInfo_T_49 ? 3'h1 : _decodeInfo_T_665;
  wire [2:0] _decodeInfo_T_667 = _decodeInfo_T_47 ? 3'h1 : _decodeInfo_T_666;
  wire [2:0] _decodeInfo_T_668 = _decodeInfo_T_45 ? 3'h1 : _decodeInfo_T_667;
  wire [2:0] _decodeInfo_T_669 = _decodeInfo_T_43 ? 3'h1 : _decodeInfo_T_668;
  wire [2:0] _decodeInfo_T_670 = _decodeInfo_T_41 ? 3'h1 : _decodeInfo_T_669;
  wire [2:0] _decodeInfo_T_671 = _decodeInfo_T_39 ? 3'h1 : _decodeInfo_T_670;
  wire [2:0] _decodeInfo_T_672 = _decodeInfo_T_37 ? 3'h1 : _decodeInfo_T_671;
  wire [2:0] _decodeInfo_T_673 = _decodeInfo_T_35 ? 3'h1 : _decodeInfo_T_672;
  wire [2:0] _decodeInfo_T_674 = _decodeInfo_T_33 ? 3'h1 : _decodeInfo_T_673;
  wire [2:0] _decodeInfo_T_675 = _decodeInfo_T_31 ? 3'h1 : _decodeInfo_T_674;
  wire [2:0] _decodeInfo_T_676 = _decodeInfo_T_29 ? 3'h1 : _decodeInfo_T_675;
  wire [2:0] _decodeInfo_T_677 = _decodeInfo_T_27 ? 3'h1 : _decodeInfo_T_676;
  wire [2:0] _decodeInfo_T_678 = _decodeInfo_T_25 ? 3'h2 : _decodeInfo_T_677;
  wire [2:0] _decodeInfo_T_679 = _decodeInfo_T_23 ? 3'h2 : _decodeInfo_T_678;
  wire [2:0] _decodeInfo_T_680 = _decodeInfo_T_21 ? 3'h2 : _decodeInfo_T_679;
  wire [2:0] _decodeInfo_T_681 = _decodeInfo_T_19 ? 3'h2 : _decodeInfo_T_680;
  wire [2:0] _decodeInfo_T_682 = _decodeInfo_T_17 ? 3'h2 : _decodeInfo_T_681;
  wire [2:0] _decodeInfo_T_683 = _decodeInfo_T_15 ? 3'h2 : _decodeInfo_T_682;
  wire [2:0] _decodeInfo_T_684 = _decodeInfo_T_13 ? 3'h2 : _decodeInfo_T_683;
  wire [2:0] _decodeInfo_T_685 = _decodeInfo_T_11 ? 3'h2 : _decodeInfo_T_684;
  wire [2:0] _decodeInfo_T_686 = _decodeInfo_T_9 ? 3'h2 : _decodeInfo_T_685;
  wire [2:0] _decodeInfo_T_687 = _decodeInfo_T_7 ? 3'h2 : _decodeInfo_T_686;
  wire [2:0] _decodeInfo_T_688 = _decodeInfo_T_5 ? 3'h2 : _decodeInfo_T_687;
  wire [2:0] _decodeInfo_T_689 = _decodeInfo_T_3 ? 3'h1 : _decodeInfo_T_688;
  wire [2:0] decodeInfo_5 = _decodeInfo_T_1 ? 3'h1 : _decodeInfo_T_689;
  wire [5:0] _decodeInfo_T_690 = _decodeInfo_T_173 ? 6'h30 : 6'h0;
  wire [5:0] _decodeInfo_T_691 = _decodeInfo_T_171 ? 6'h2f : _decodeInfo_T_690;
  wire [5:0] _decodeInfo_T_692 = _decodeInfo_T_169 ? 6'h2e : _decodeInfo_T_691;
  wire [5:0] _decodeInfo_T_693 = _decodeInfo_T_167 ? 6'h30 : _decodeInfo_T_692;
  wire [5:0] _decodeInfo_T_694 = _decodeInfo_T_165 ? 6'h2e : _decodeInfo_T_693;
  wire [5:0] _decodeInfo_T_695 = _decodeInfo_T_163 ? 6'h2f : _decodeInfo_T_694;
  wire [5:0] _decodeInfo_T_696 = _decodeInfo_T_161 ? 6'h31 : _decodeInfo_T_695;
  wire [5:0] _decodeInfo_T_697 = _decodeInfo_T_159 ? 6'h31 : _decodeInfo_T_696;
  wire [5:0] _decodeInfo_T_698 = _decodeInfo_T_157 ? 6'h31 : _decodeInfo_T_697;
  wire [5:0] _decodeInfo_T_699 = _decodeInfo_T_155 ? 6'h31 : _decodeInfo_T_698;
  wire [5:0] _decodeInfo_T_700 = _decodeInfo_T_153 ? 6'h2c : _decodeInfo_T_699;
  wire [5:0] _decodeInfo_T_701 = _decodeInfo_T_151 ? 6'h2b : _decodeInfo_T_700;
  wire [5:0] _decodeInfo_T_702 = _decodeInfo_T_149 ? 6'h2a : _decodeInfo_T_701;
  wire [5:0] _decodeInfo_T_703 = _decodeInfo_T_121 ? 6'h27 : _decodeInfo_T_702;
  wire [5:0] _decodeInfo_T_704 = _decodeInfo_T_119 ? 6'h26 : _decodeInfo_T_703;
  wire [5:0] _decodeInfo_T_705 = _decodeInfo_T_117 ? 6'h29 : _decodeInfo_T_704;
  wire [5:0] _decodeInfo_T_706 = _decodeInfo_T_115 ? 6'h28 : _decodeInfo_T_705;
  wire [5:0] _decodeInfo_T_707 = _decodeInfo_T_113 ? 6'h25 : _decodeInfo_T_706;
  wire [5:0] _decodeInfo_T_708 = _decodeInfo_T_111 ? 6'h24 : _decodeInfo_T_707;
  wire [5:0] _decodeInfo_T_709 = _decodeInfo_T_135 ? 6'h23 : _decodeInfo_T_708;
  wire [5:0] _decodeInfo_T_710 = _decodeInfo_T_109 ? 6'h22 : _decodeInfo_T_709;
  wire [5:0] _decodeInfo_T_711 = _decodeInfo_T_107 ? 6'h21 : _decodeInfo_T_710;
  wire [5:0] _decodeInfo_T_712 = _decodeInfo_T_105 ? 6'h1f : _decodeInfo_T_711;
  wire [5:0] _decodeInfo_T_713 = _decodeInfo_T_103 ? 6'h20 : _decodeInfo_T_712;
  wire [5:0] _decodeInfo_T_714 = _decodeInfo_T_101 ? 6'h1e : _decodeInfo_T_713;
  wire [5:0] _decodeInfo_T_715 = _decodeInfo_T_99 ? 6'h1d : _decodeInfo_T_714;
  wire [5:0] _decodeInfo_T_716 = _decodeInfo_T_121 ? 6'h27 : _decodeInfo_T_715;
  wire [5:0] _decodeInfo_T_717 = _decodeInfo_T_119 ? 6'h26 : _decodeInfo_T_716;
  wire [5:0] _decodeInfo_T_718 = _decodeInfo_T_117 ? 6'h29 : _decodeInfo_T_717;
  wire [5:0] _decodeInfo_T_719 = _decodeInfo_T_115 ? 6'h28 : _decodeInfo_T_718;
  wire [5:0] _decodeInfo_T_720 = _decodeInfo_T_113 ? 6'h25 : _decodeInfo_T_719;
  wire [5:0] _decodeInfo_T_721 = _decodeInfo_T_111 ? 6'h24 : _decodeInfo_T_720;
  wire [5:0] _decodeInfo_T_722 = _decodeInfo_T_109 ? 6'h22 : _decodeInfo_T_721;
  wire [5:0] _decodeInfo_T_723 = _decodeInfo_T_107 ? 6'h21 : _decodeInfo_T_722;
  wire [5:0] _decodeInfo_T_724 = _decodeInfo_T_105 ? 6'h1f : _decodeInfo_T_723;
  wire [5:0] _decodeInfo_T_725 = _decodeInfo_T_103 ? 6'h20 : _decodeInfo_T_724;
  wire [5:0] _decodeInfo_T_726 = _decodeInfo_T_101 ? 6'h1e : _decodeInfo_T_725;
  wire [5:0] _decodeInfo_T_727 = _decodeInfo_T_99 ? 6'h1d : _decodeInfo_T_726;
  wire [5:0] _decodeInfo_T_728 = _decodeInfo_T_97 ? 6'h0 : _decodeInfo_T_727;
  wire [5:0] _decodeInfo_T_729 = _decodeInfo_T_95 ? 6'h0 : _decodeInfo_T_728;
  wire [5:0] _decodeInfo_T_730 = _decodeInfo_T_93 ? 6'h0 : _decodeInfo_T_729;
  wire [5:0] _decodeInfo_T_731 = _decodeInfo_T_91 ? 6'h0 : _decodeInfo_T_730;
  wire [5:0] _decodeInfo_T_732 = _decodeInfo_T_89 ? 6'h0 : _decodeInfo_T_731;
  wire [5:0] _decodeInfo_T_733 = _decodeInfo_T_87 ? 6'h0 : _decodeInfo_T_732;
  wire [5:0] _decodeInfo_T_734 = _decodeInfo_T_85 ? 6'h0 : _decodeInfo_T_733;
  wire [5:0] _decodeInfo_T_735 = _decodeInfo_T_83 ? 6'h0 : _decodeInfo_T_734;
  wire [5:0] _decodeInfo_T_736 = _decodeInfo_T_81 ? 6'h10 : _decodeInfo_T_735;
  wire [5:0] _decodeInfo_T_737 = _decodeInfo_T_79 ? 6'hf : _decodeInfo_T_736;
  wire [5:0] _decodeInfo_T_738 = _decodeInfo_T_77 ? 6'he : _decodeInfo_T_737;
  wire [5:0] _decodeInfo_T_739 = _decodeInfo_T_75 ? 6'hc : _decodeInfo_T_738;
  wire [5:0] _decodeInfo_T_740 = _decodeInfo_T_73 ? 6'h10 : _decodeInfo_T_739;
  wire [5:0] _decodeInfo_T_741 = _decodeInfo_T_71 ? 6'hf : _decodeInfo_T_740;
  wire [5:0] _decodeInfo_T_742 = _decodeInfo_T_69 ? 6'he : _decodeInfo_T_741;
  wire [5:0] _decodeInfo_T_743 = _decodeInfo_T_67 ? 6'hd : _decodeInfo_T_742;
  wire [5:0] _decodeInfo_T_744 = _decodeInfo_T_65 ? 6'hc : _decodeInfo_T_743;
  wire [5:0] _decodeInfo_T_745 = _decodeInfo_T_63 ? 6'h5 : _decodeInfo_T_744;
  wire [5:0] _decodeInfo_T_746 = _decodeInfo_T_61 ? 6'h6 : _decodeInfo_T_745;
  wire [5:0] _decodeInfo_T_747 = _decodeInfo_T_59 ? 6'h4 : _decodeInfo_T_746;
  wire [5:0] _decodeInfo_T_748 = _decodeInfo_T_57 ? 6'ha : _decodeInfo_T_747;
  wire [5:0] _decodeInfo_T_749 = _decodeInfo_T_55 ? 6'h9 : _decodeInfo_T_748;
  wire [5:0] _decodeInfo_T_750 = _decodeInfo_T_53 ? 6'h8 : _decodeInfo_T_749;
  wire [5:0] _decodeInfo_T_751 = _decodeInfo_T_51 ? 6'h7 : _decodeInfo_T_750;
  wire [5:0] _decodeInfo_T_752 = _decodeInfo_T_49 ? 6'h3 : _decodeInfo_T_751;
  wire [5:0] _decodeInfo_T_753 = _decodeInfo_T_47 ? 6'h2 : _decodeInfo_T_752;
  wire [5:0] _decodeInfo_T_754 = _decodeInfo_T_45 ? 6'h5 : _decodeInfo_T_753;
  wire [5:0] _decodeInfo_T_755 = _decodeInfo_T_43 ? 6'h6 : _decodeInfo_T_754;
  wire [5:0] _decodeInfo_T_756 = _decodeInfo_T_41 ? 6'h4 : _decodeInfo_T_755;
  wire [5:0] _decodeInfo_T_757 = _decodeInfo_T_39 ? 6'hb : _decodeInfo_T_756;
  wire [5:0] _decodeInfo_T_758 = _decodeInfo_T_37 ? 6'ha : _decodeInfo_T_757;
  wire [5:0] _decodeInfo_T_759 = _decodeInfo_T_35 ? 6'hb : _decodeInfo_T_758;
  wire [5:0] _decodeInfo_T_760 = _decodeInfo_T_33 ? 6'h9 : _decodeInfo_T_759;
  wire [5:0] _decodeInfo_T_761 = _decodeInfo_T_31 ? 6'h8 : _decodeInfo_T_760;
  wire [5:0] _decodeInfo_T_762 = _decodeInfo_T_29 ? 6'h7 : _decodeInfo_T_761;
  wire [5:0] _decodeInfo_T_763 = _decodeInfo_T_27 ? 6'h2 : _decodeInfo_T_762;
  wire [5:0] _decodeInfo_T_764 = _decodeInfo_T_25 ? 6'h1c : _decodeInfo_T_763;
  wire [5:0] _decodeInfo_T_765 = _decodeInfo_T_23 ? 6'h19 : _decodeInfo_T_764;
  wire [5:0] _decodeInfo_T_766 = _decodeInfo_T_21 ? 6'h1a : _decodeInfo_T_765;
  wire [5:0] _decodeInfo_T_767 = _decodeInfo_T_19 ? 6'h1b : _decodeInfo_T_766;
  wire [5:0] _decodeInfo_T_768 = _decodeInfo_T_17 ? 6'h16 : _decodeInfo_T_767;
  wire [5:0] _decodeInfo_T_769 = _decodeInfo_T_15 ? 6'h17 : _decodeInfo_T_768;
  wire [5:0] _decodeInfo_T_770 = _decodeInfo_T_13 ? 6'h18 : _decodeInfo_T_769;
  wire [5:0] _decodeInfo_T_771 = _decodeInfo_T_11 ? 6'h15 : _decodeInfo_T_770;
  wire [5:0] _decodeInfo_T_772 = _decodeInfo_T_9 ? 6'h12 : _decodeInfo_T_771;
  wire [5:0] _decodeInfo_T_773 = _decodeInfo_T_7 ? 6'h13 : _decodeInfo_T_772;
  wire [5:0] _decodeInfo_T_774 = _decodeInfo_T_5 ? 6'h14 : _decodeInfo_T_773;
  wire [5:0] _decodeInfo_T_775 = _decodeInfo_T_3 ? 6'h11 : _decodeInfo_T_774;
  wire [5:0] decodeInfo_6 = _decodeInfo_T_1 ? 6'h2 : _decodeInfo_T_775;
  wire  _decodeInfo_T_814 = _decodeInfo_T_97 ? 1'h0 : _decodeInfo_T_99 | (_decodeInfo_T_101 | (_decodeInfo_T_103 | (
    _decodeInfo_T_105 | (_decodeInfo_T_107 | (_decodeInfo_T_109 | (_decodeInfo_T_111 | (_decodeInfo_T_113 | (
    _decodeInfo_T_115 | (_decodeInfo_T_117 | (_decodeInfo_T_119 | (_decodeInfo_T_121 | (_decodeInfo_T_99 | (
    _decodeInfo_T_101 | (_decodeInfo_T_103 | (_decodeInfo_T_105 | (_decodeInfo_T_107 | (_decodeInfo_T_109 | (
    _decodeInfo_T_135 | (_decodeInfo_T_111 | (_decodeInfo_T_113 | (_decodeInfo_T_115 | (_decodeInfo_T_117 | (
    _decodeInfo_T_119 | (_decodeInfo_T_121 | _decodeInfo_T_444))))))))))))))))))))))));
  wire  _decodeInfo_T_815 = _decodeInfo_T_95 ? 1'h0 : _decodeInfo_T_814;
  wire  _decodeInfo_T_816 = _decodeInfo_T_93 ? 1'h0 : _decodeInfo_T_815;
  wire  _decodeInfo_T_817 = _decodeInfo_T_91 ? 1'h0 : _decodeInfo_T_816;
  wire  _decodeInfo_T_818 = _decodeInfo_T_89 ? 1'h0 : _decodeInfo_T_817;
  wire  _decodeInfo_T_819 = _decodeInfo_T_87 ? 1'h0 : _decodeInfo_T_818;
  wire [1:0] _decodeInfo_T_820 = _decodeInfo_T_85 ? 2'h2 : {{1'd0}, _decodeInfo_T_819};
  wire [1:0] _decodeInfo_T_821 = _decodeInfo_T_83 ? 2'h2 : _decodeInfo_T_820;
  wire [1:0] _decodeInfo_T_822 = _decodeInfo_T_81 ? 2'h1 : _decodeInfo_T_821;
  wire [1:0] _decodeInfo_T_823 = _decodeInfo_T_79 ? 2'h1 : _decodeInfo_T_822;
  wire [1:0] _decodeInfo_T_824 = _decodeInfo_T_77 ? 2'h1 : _decodeInfo_T_823;
  wire [1:0] _decodeInfo_T_825 = _decodeInfo_T_75 ? 2'h1 : _decodeInfo_T_824;
  wire [1:0] _decodeInfo_T_826 = _decodeInfo_T_73 ? 2'h1 : _decodeInfo_T_825;
  wire [1:0] _decodeInfo_T_827 = _decodeInfo_T_71 ? 2'h1 : _decodeInfo_T_826;
  wire [1:0] _decodeInfo_T_828 = _decodeInfo_T_69 ? 2'h1 : _decodeInfo_T_827;
  wire [1:0] _decodeInfo_T_829 = _decodeInfo_T_67 ? 2'h1 : _decodeInfo_T_828;
  wire [1:0] _decodeInfo_T_830 = _decodeInfo_T_65 ? 2'h1 : _decodeInfo_T_829;
  wire [1:0] _decodeInfo_T_831 = _decodeInfo_T_63 ? 2'h1 : _decodeInfo_T_830;
  wire [1:0] _decodeInfo_T_832 = _decodeInfo_T_61 ? 2'h1 : _decodeInfo_T_831;
  wire [1:0] _decodeInfo_T_833 = _decodeInfo_T_59 ? 2'h1 : _decodeInfo_T_832;
  wire [1:0] _decodeInfo_T_834 = _decodeInfo_T_57 ? 2'h1 : _decodeInfo_T_833;
  wire [1:0] _decodeInfo_T_835 = _decodeInfo_T_55 ? 2'h1 : _decodeInfo_T_834;
  wire [1:0] _decodeInfo_T_836 = _decodeInfo_T_53 ? 2'h1 : _decodeInfo_T_835;
  wire [1:0] _decodeInfo_T_837 = _decodeInfo_T_51 ? 2'h1 : _decodeInfo_T_836;
  wire [1:0] _decodeInfo_T_838 = _decodeInfo_T_49 ? 2'h1 : _decodeInfo_T_837;
  wire [1:0] _decodeInfo_T_839 = _decodeInfo_T_47 ? 2'h1 : _decodeInfo_T_838;
  wire [1:0] _decodeInfo_T_840 = _decodeInfo_T_45 ? 2'h1 : _decodeInfo_T_839;
  wire [1:0] _decodeInfo_T_841 = _decodeInfo_T_43 ? 2'h1 : _decodeInfo_T_840;
  wire [1:0] _decodeInfo_T_842 = _decodeInfo_T_41 ? 2'h1 : _decodeInfo_T_841;
  wire [1:0] _decodeInfo_T_843 = _decodeInfo_T_39 ? 2'h1 : _decodeInfo_T_842;
  wire [1:0] _decodeInfo_T_844 = _decodeInfo_T_37 ? 2'h1 : _decodeInfo_T_843;
  wire [1:0] _decodeInfo_T_845 = _decodeInfo_T_35 ? 2'h1 : _decodeInfo_T_844;
  wire [1:0] _decodeInfo_T_846 = _decodeInfo_T_33 ? 2'h1 : _decodeInfo_T_845;
  wire [1:0] _decodeInfo_T_847 = _decodeInfo_T_31 ? 2'h1 : _decodeInfo_T_846;
  wire [1:0] _decodeInfo_T_848 = _decodeInfo_T_29 ? 2'h1 : _decodeInfo_T_847;
  wire [1:0] _decodeInfo_T_849 = _decodeInfo_T_27 ? 2'h1 : _decodeInfo_T_848;
  wire [1:0] _decodeInfo_T_850 = _decodeInfo_T_25 ? 2'h0 : _decodeInfo_T_849;
  wire [1:0] _decodeInfo_T_851 = _decodeInfo_T_23 ? 2'h0 : _decodeInfo_T_850;
  wire [1:0] _decodeInfo_T_852 = _decodeInfo_T_21 ? 2'h0 : _decodeInfo_T_851;
  wire [1:0] _decodeInfo_T_853 = _decodeInfo_T_19 ? 2'h0 : _decodeInfo_T_852;
  wire [1:0] _decodeInfo_T_854 = _decodeInfo_T_17 ? 2'h1 : _decodeInfo_T_853;
  wire [1:0] _decodeInfo_T_855 = _decodeInfo_T_15 ? 2'h1 : _decodeInfo_T_854;
  wire [1:0] _decodeInfo_T_856 = _decodeInfo_T_13 ? 2'h1 : _decodeInfo_T_855;
  wire [1:0] _decodeInfo_T_857 = _decodeInfo_T_11 ? 2'h1 : _decodeInfo_T_856;
  wire [1:0] _decodeInfo_T_858 = _decodeInfo_T_9 ? 2'h1 : _decodeInfo_T_857;
  wire [1:0] _decodeInfo_T_859 = _decodeInfo_T_7 ? 2'h1 : _decodeInfo_T_858;
  wire [1:0] _decodeInfo_T_860 = _decodeInfo_T_5 ? 2'h1 : _decodeInfo_T_859;
  wire [1:0] _decodeInfo_T_861 = _decodeInfo_T_3 ? 2'h1 : _decodeInfo_T_860;
  wire [1:0] decodeInfo_7 = _decodeInfo_T_1 ? 2'h1 : _decodeInfo_T_861;
  wire  _decodeInfo_T_892 = _decodeInfo_T_113 | (_decodeInfo_T_115 | (_decodeInfo_T_117 | (_decodeInfo_T_119 | (
    _decodeInfo_T_121 | (_decodeInfo_T_99 | (_decodeInfo_T_101 | (_decodeInfo_T_103 | (_decodeInfo_T_105 | (
    _decodeInfo_T_107 | (_decodeInfo_T_109 | (_decodeInfo_T_135 | (_decodeInfo_T_111 | (_decodeInfo_T_113 | (
    _decodeInfo_T_115 | (_decodeInfo_T_117 | (_decodeInfo_T_119 | (_decodeInfo_T_121 | (_decodeInfo_T_149 | (
    _decodeInfo_T_151 | (_decodeInfo_T_153 | (_decodeInfo_T_155 | (_decodeInfo_T_157 | (_decodeInfo_T_159 | (
    _decodeInfo_T_161 | (_decodeInfo_T_163 | (_decodeInfo_T_165 | (_decodeInfo_T_167 | (_decodeInfo_T_169 | (
    _decodeInfo_T_171 | _decodeInfo_T_173)))))))))))))))))))))))))))));
  wire  _decodeInfo_T_900 = _decodeInfo_T_97 ? 1'h0 : _decodeInfo_T_99 | (_decodeInfo_T_101 | (_decodeInfo_T_103 | (
    _decodeInfo_T_105 | (_decodeInfo_T_107 | (_decodeInfo_T_109 | (_decodeInfo_T_111 | _decodeInfo_T_892))))));
  wire  _decodeInfo_T_901 = _decodeInfo_T_95 ? 1'h0 : _decodeInfo_T_900;
  wire  _decodeInfo_T_902 = _decodeInfo_T_93 ? 1'h0 : _decodeInfo_T_901;
  wire  _decodeInfo_T_903 = _decodeInfo_T_91 ? 1'h0 : _decodeInfo_T_902;
  wire  _decodeInfo_T_904 = _decodeInfo_T_89 ? 1'h0 : _decodeInfo_T_903;
  wire  _decodeInfo_T_905 = _decodeInfo_T_87 ? 1'h0 : _decodeInfo_T_904;
  wire  _decodeInfo_T_935 = _decodeInfo_T_27 | (_decodeInfo_T_29 | (_decodeInfo_T_31 | (_decodeInfo_T_33 | (
    _decodeInfo_T_35 | (_decodeInfo_T_37 | (_decodeInfo_T_39 | (_decodeInfo_T_41 | (_decodeInfo_T_43 | (_decodeInfo_T_45
     | (_decodeInfo_T_47 | (_decodeInfo_T_49 | (_decodeInfo_T_51 | (_decodeInfo_T_53 | (_decodeInfo_T_55 | (
    _decodeInfo_T_57 | (_decodeInfo_T_59 | (_decodeInfo_T_61 | (_decodeInfo_T_63 | (_decodeInfo_T_65 | (_decodeInfo_T_67
     | (_decodeInfo_T_69 | (_decodeInfo_T_71 | (_decodeInfo_T_73 | (_decodeInfo_T_75 | (_decodeInfo_T_77 | (
    _decodeInfo_T_79 | (_decodeInfo_T_81 | (_decodeInfo_T_83 | (_decodeInfo_T_85 | _decodeInfo_T_905))))))))))))))))))))
    )))))))));
  wire  _decodeInfo_T_936 = _decodeInfo_T_25 ? 1'h0 : _decodeInfo_T_935;
  wire  _decodeInfo_T_937 = _decodeInfo_T_23 ? 1'h0 : _decodeInfo_T_936;
  wire  _decodeInfo_T_938 = _decodeInfo_T_21 ? 1'h0 : _decodeInfo_T_937;
  wire  _decodeInfo_T_939 = _decodeInfo_T_19 ? 1'h0 : _decodeInfo_T_938;
  wire  decodeInfo_8 = _decodeInfo_T_1 | (_decodeInfo_T_3 | (_decodeInfo_T_5 | (_decodeInfo_T_7 | (_decodeInfo_T_9 | (
    _decodeInfo_T_11 | (_decodeInfo_T_13 | (_decodeInfo_T_15 | (_decodeInfo_T_17 | _decodeInfo_T_939))))))));
  wire [11:0] imm_i = decodeBuffer_inst[31:20];
  wire [19:0] imm_u = decodeBuffer_inst[31:12];
  wire [63:0] imm_z = {59'h0,dec_rs_addr_0};
  wire [51:0] _imm_i_sext_T_2 = imm_i[11] ? 52'hfffffffffffff : 52'h0;
  wire [63:0] imm_i_sext = {_imm_i_sext_T_2,imm_i};
  wire [51:0] _imm_s_sext_T_2 = decodeBuffer_inst[31] ? 52'hfffffffffffff : 52'h0;
  wire [63:0] imm_s_sext = {_imm_s_sext_T_2,decodeBuffer_inst[31:25],decodeBuffer_inst[11:7]};
  wire [50:0] _imm_b_sext_T_2 = decodeBuffer_inst[31] ? 51'h7ffffffffffff : 51'h0;
  wire [63:0] imm_b_sext = {_imm_b_sext_T_2,decodeBuffer_inst[31],decodeBuffer_inst[7],decodeBuffer_inst[30:25],
    decodeBuffer_inst[11:8],1'h0};
  wire [31:0] _imm_u_sext_T_2 = imm_u[19] ? 32'hffffffff : 32'h0;
  wire [63:0] imm_u_sext = {_imm_u_sext_T_2,imm_u,12'h0};
  wire [42:0] _imm_j_sext_T_2 = decodeBuffer_inst[31] ? 43'h7ffffffffff : 43'h0;
  wire [63:0] imm_j_sext = {_imm_j_sext_T_2,decodeBuffer_inst[31],decodeBuffer_inst[19:12],decodeBuffer_inst[20],
    decodeBuffer_inst[30:21],1'h0};
  wire [31:0] _GEN_1 = io_flush ? 32'h13 : decodeBuffer_inst;
  wire [31:0] _GEN_2 = io_flush ? 32'h0 : decodeBuffer_pc;
  wire  _GEN_3 = io_flush | decodeBuffer_bubble;
  wire  _T = io_out_ready & io_out_valid;
  wire  _T_1 = io_in_ready & io_in_valid;
  wire  _T_4 = ~io_flush;
  wire  _GEN_8 = ~_T_1 & _T | io_flush | _GEN_3;
  wire  _GEN_12 = _T_1 & _T & ~io_flush ? 1'h0 : _GEN_8;
  wire  _GEN_18 = needWait ? _GEN_3 : _GEN_12;
  wire  _rs1_data_T_1 = dec_rs_addr_0 != 5'h0;
  wire  _rs1_data_T_3 = io_bypass_0_addr == dec_rs_addr_0 & dec_rs_addr_0 != 5'h0 & io_bypass_0_rf_wen;
  wire  _rs1_data_T_7 = io_bypass_1_addr == dec_rs_addr_0 & _rs1_data_T_1 & io_bypass_1_rf_wen;
  wire [63:0] _rs1_data_T_8 = _rs1_data_T_7 ? io_bypass_1_data : io_regFile_rs1_data;
  wire [63:0] rs1_data = _rs1_data_T_3 ? io_bypass_0_data : _rs1_data_T_8;
  wire  _rs2_data_T_1 = dec_rs_addr_1 != 5'h0;
  wire  _rs2_data_T_3 = io_bypass_0_addr == dec_rs_addr_1 & dec_rs_addr_1 != 5'h0 & io_bypass_0_rf_wen;
  wire  _rs2_data_T_7 = io_bypass_1_addr == dec_rs_addr_1 & _rs2_data_T_1 & io_bypass_1_rf_wen;
  wire [63:0] _rs2_data_T_8 = _rs2_data_T_7 ? io_bypass_1_data : io_regFile_rs2_data;
  wire [63:0] rs2_data = _rs2_data_T_3 ? io_bypass_0_data : _rs2_data_T_8;
  wire [63:0] _dec_op1_data_T_2 = 3'h1 == decodeInfo_1 ? imm_u_sext : 64'hdeadc0de;
  wire [63:0] _dec_op1_data_T_4 = 3'h2 == decodeInfo_1 ? rs1_data : _dec_op1_data_T_2;
  wire [63:0] _dec_op1_data_T_6 = 3'h3 == decodeInfo_1 ? imm_j_sext : _dec_op1_data_T_4;
  wire [63:0] _dec_op1_data_T_8 = 3'h4 == decodeInfo_1 ? imm_i_sext : _dec_op1_data_T_6;
  wire [63:0] _dec_op1_data_T_10 = 3'h5 == decodeInfo_1 ? imm_z : _dec_op1_data_T_8;
  wire [63:0] _dec_op1_data_T_12 = 3'h6 == decodeInfo_1 ? rs2_data : _dec_op1_data_T_10;
  wire [63:0] _dec_op1_data_T_14 = 3'h7 == decodeInfo_1 ? {{32'd0}, decodeBuffer_pc} : _dec_op1_data_T_12;
  wire [3:0] _GEN_19 = {{1'd0}, decodeInfo_1};
  wire [63:0] _dec_op1_data_T_16 = 4'h8 == _GEN_19 ? imm_s_sext : _dec_op1_data_T_14;
  wire [63:0] dec_op1_data = 4'h9 == _GEN_19 ? imm_b_sext : _dec_op1_data_T_16;
  wire [63:0] _dec_op2_data_T_2 = 4'h1 == decodeInfo_2 ? imm_u_sext : 64'hdeadc0de;
  wire [63:0] _dec_op2_data_T_4 = 4'h2 == decodeInfo_2 ? rs1_data : _dec_op2_data_T_2;
  wire [63:0] _dec_op2_data_T_6 = 4'h3 == decodeInfo_2 ? imm_j_sext : _dec_op2_data_T_4;
  wire [63:0] _dec_op2_data_T_8 = 4'h4 == decodeInfo_2 ? imm_i_sext : _dec_op2_data_T_6;
  wire [63:0] _dec_op2_data_T_10 = 4'h5 == decodeInfo_2 ? imm_z : _dec_op2_data_T_8;
  wire [63:0] _dec_op2_data_T_12 = 4'h6 == decodeInfo_2 ? rs2_data : _dec_op2_data_T_10;
  wire [63:0] _dec_op2_data_T_14 = 4'h7 == decodeInfo_2 ? {{32'd0}, decodeBuffer_pc} : _dec_op2_data_T_12;
  wire [63:0] _dec_op2_data_T_16 = 4'h8 == decodeInfo_2 ? imm_s_sext : _dec_op2_data_T_14;
  wire [63:0] dec_op2_data = 4'h9 == decodeInfo_2 ? imm_b_sext : _dec_op2_data_T_16;
  wire  isCSR = decodeInfo_5 == 3'h3;
  wire  csr_en = isCSR & (decodeInfo_6 == 6'h2f | decodeInfo_6 == 6'h30) & (decodeInfo_3 & dec_rs_addr_0 == 5'h0);
  wire [5:0] opcode_func = csr_en ? 6'h32 : decodeInfo_6;
  assign io_in_ready = io_out_ready & ~needWait;
  assign io_out_valid = 1'h1;
  assign io_out_bits_pc = needWait ? 32'h0 : decodeBuffer_pc;
  assign io_out_bits_inst = needWait ? 32'h13 : decodeBuffer_inst;
  assign io_out_bits_valid = _io_in_ready_T & _T_4;
  assign io_out_bits_bubble = decodeBuffer_bubble;
  assign io_out_bits_opcode_type = needWait ? 3'h1 : decodeInfo_5;
  assign io_out_bits_opcode_func = needWait ? 6'h2 : opcode_func;
  assign io_out_bits_br_type = _decodeInfo_T_1 ? 4'h0 : _decodeInfo_T_259;
  assign io_out_bits_rf_en = needWait ? 1'h0 : decodeInfo_8;
  assign io_out_bits_wb_addr = needWait ? 5'h0 : decodeBuffer_inst[11:7];
  assign io_out_bits_wb_stage = needWait ? 2'h0 : decodeInfo_7;
  assign io_out_bits_op1_data = needWait ? 64'h0 : dec_op1_data;
  assign io_out_bits_op2_data = needWait ? 64'h0 : dec_op2_data;
  assign io_out_bits_rs1_data = needWait ? 64'h0 : rs1_data;
  assign io_out_bits_rs2_data = needWait ? 64'h0 : rs2_data;
  assign io_regFile_rs1_addr = decodeBuffer_inst[19:15];
  assign io_regFile_rs2_addr = decodeBuffer_inst[24:20];
  always @(posedge clock) begin
    if (reset) begin
      last_use_rd <= 5'h0;
    end else if (needWait) begin
      if (_T) begin
        last_use_rd <= 5'h0;
      end
    end else if (_T_1 & _T & ~io_flush) begin
      if (~decodeInfo_8) begin
        last_use_rd <= 5'h0;
      end else begin
        last_use_rd <= decodeBuffer_inst[11:7];
      end
    end
    if (reset) begin
      decodeBuffer_inst <= 32'h13;
    end else if (needWait) begin
      decodeBuffer_inst <= _GEN_1;
    end else if (_T_1 & _T & ~io_flush) begin
      decodeBuffer_inst <= io_in_bits_inst;
    end else if (~_T_1 & _T | io_flush) begin
      decodeBuffer_inst <= 32'h13;
    end else begin
      decodeBuffer_inst <= _GEN_1;
    end
    if (reset) begin
      decodeBuffer_pc <= 32'h0;
    end else if (needWait) begin
      decodeBuffer_pc <= _GEN_2;
    end else if (_T_1 & _T & ~io_flush) begin
      decodeBuffer_pc <= io_in_bits_pc;
    end else if (~_T_1 & _T | io_flush) begin
      decodeBuffer_pc <= 32'h0;
    end else begin
      decodeBuffer_pc <= _GEN_2;
    end
    decodeBuffer_bubble <= reset | _GEN_18;
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_use_rd = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  decodeBuffer_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  decodeBuffer_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  decodeBuffer_bubble = _RAND_3[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Alu(
  input  [63:0] io_in_bits_op1_data,
  input  [63:0] io_in_bits_op2_data,
  input  [5:0]  io_in_bits_func,
  output [63:0] io_out_bits
);
  wire [5:0] alu_shamt = io_in_bits_op2_data[5:0];
  wire [63:0] _alu_out_T_3 = io_in_bits_op1_data + io_in_bits_op2_data;
  wire [63:0] _alu_out_T_9 = io_in_bits_op1_data - io_in_bits_op2_data;
  wire [63:0] _alu_out_T_14 = io_in_bits_op1_data & io_in_bits_op2_data;
  wire [63:0] _alu_out_T_16 = io_in_bits_op1_data | io_in_bits_op2_data;
  wire [63:0] _alu_out_T_18 = io_in_bits_op1_data ^ io_in_bits_op2_data;
  wire  _alu_out_T_22 = $signed(io_in_bits_op1_data) < $signed(io_in_bits_op2_data);
  wire  _alu_out_T_24 = io_in_bits_op1_data < io_in_bits_op2_data;
  wire [126:0] _GEN_0 = {{63'd0}, io_in_bits_op1_data};
  wire [126:0] _alu_out_T_26 = _GEN_0 << alu_shamt;
  wire [62:0] _GEN_1 = {{31'd0}, io_in_bits_op1_data[31:0]};
  wire [62:0] _alu_out_T_30 = _GEN_1 << alu_shamt[4:0];
  wire [63:0] _alu_out_T_34 = $signed(io_in_bits_op1_data) >>> alu_shamt;
  wire [31:0] _alu_out_T_37 = io_in_bits_op1_data[31:0];
  wire [31:0] _alu_out_T_40 = $signed(_alu_out_T_37) >>> alu_shamt[4:0];
  wire [63:0] _alu_out_T_42 = io_in_bits_op1_data >> alu_shamt;
  wire [31:0] _alu_out_T_46 = io_in_bits_op1_data[31:0] >> alu_shamt[4:0];
  wire [63:0] _alu_out_T_49 = 6'h2 == io_in_bits_func ? _alu_out_T_3 : 64'h0;
  wire [63:0] _alu_out_T_51 = 6'hc == io_in_bits_func ? _alu_out_T_3 : _alu_out_T_49;
  wire [63:0] _alu_out_T_53 = 6'h3 == io_in_bits_func ? _alu_out_T_9 : _alu_out_T_51;
  wire [63:0] _alu_out_T_55 = 6'hd == io_in_bits_func ? _alu_out_T_9 : _alu_out_T_53;
  wire [63:0] _alu_out_T_57 = 6'h7 == io_in_bits_func ? _alu_out_T_14 : _alu_out_T_55;
  wire [63:0] _alu_out_T_59 = 6'h8 == io_in_bits_func ? _alu_out_T_16 : _alu_out_T_57;
  wire [63:0] _alu_out_T_61 = 6'h9 == io_in_bits_func ? _alu_out_T_18 : _alu_out_T_59;
  wire [63:0] _alu_out_T_63 = 6'ha == io_in_bits_func ? {{63'd0}, _alu_out_T_22} : _alu_out_T_61;
  wire [63:0] _alu_out_T_65 = 6'hb == io_in_bits_func ? {{63'd0}, _alu_out_T_24} : _alu_out_T_63;
  wire [126:0] _alu_out_T_67 = 6'h4 == io_in_bits_func ? _alu_out_T_26 : {{63'd0}, _alu_out_T_65};
  wire [126:0] _alu_out_T_69 = 6'he == io_in_bits_func ? {{64'd0}, _alu_out_T_30} : _alu_out_T_67;
  wire [126:0] _alu_out_T_71 = 6'h6 == io_in_bits_func ? {{63'd0}, _alu_out_T_34} : _alu_out_T_69;
  wire [126:0] _alu_out_T_73 = 6'h10 == io_in_bits_func ? {{95'd0}, _alu_out_T_40} : _alu_out_T_71;
  wire [126:0] _alu_out_T_75 = 6'h5 == io_in_bits_func ? {{63'd0}, _alu_out_T_42} : _alu_out_T_73;
  wire [126:0] _alu_out_T_77 = 6'hf == io_in_bits_func ? {{95'd0}, _alu_out_T_46} : _alu_out_T_75;
  wire [126:0] _alu_out_T_79 = 6'h11 == io_in_bits_func ? {{63'd0}, io_in_bits_op1_data} : _alu_out_T_77;
  wire [63:0] alu_out = _alu_out_T_79[63:0];
  wire [31:0] _io_out_bits_T_4 = alu_out[31] ? 32'hffffffff : 32'h0;
  wire [63:0] _io_out_bits_T_6 = {_io_out_bits_T_4,alu_out[31:0]};
  wire [63:0] _io_out_bits_T_32 = 6'hc == io_in_bits_func ? _io_out_bits_T_6 : alu_out;
  wire [63:0] _io_out_bits_T_34 = 6'hd == io_in_bits_func ? _io_out_bits_T_6 : _io_out_bits_T_32;
  wire [63:0] _io_out_bits_T_36 = 6'he == io_in_bits_func ? _io_out_bits_T_6 : _io_out_bits_T_34;
  wire [63:0] _io_out_bits_T_38 = 6'h10 == io_in_bits_func ? _io_out_bits_T_6 : _io_out_bits_T_36;
  assign io_out_bits = 6'hf == io_in_bits_func ? _io_out_bits_T_6 : _io_out_bits_T_38;
endmodule
module ysyx_040656_Jmp(
  input         io_in_valid,
  input  [63:0] io_in_bits_op1_data,
  input  [63:0] io_in_bits_op2_data,
  input  [63:0] io_in_bits_rs1_data,
  input  [63:0] io_in_bits_rs2_data,
  input  [3:0]  io_in_bits_br_type,
  input  [31:0] io_in_bits_pc,
  output        io_out_bits_redirect_valid,
  output [31:0] io_out_bits_redirect_target
);
  wire  br_eq = io_in_bits_rs2_data == io_in_bits_rs1_data;
  wire  br_lt = $signed(io_in_bits_rs2_data) < $signed(io_in_bits_rs1_data);
  wire  br_ltu = io_in_bits_rs2_data < io_in_bits_rs1_data;
  wire [1:0] _exe_ctrl_pc_sel_T_4 = ~br_eq ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_6 = br_eq ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_9 = ~br_lt ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_12 = ~br_ltu ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_14 = br_lt ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_16 = br_ltu ? 2'h0 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_24 = 4'h1 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_4 : 2'h3;
  wire [1:0] _exe_ctrl_pc_sel_T_26 = 4'h2 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_6 : _exe_ctrl_pc_sel_T_24;
  wire [1:0] _exe_ctrl_pc_sel_T_28 = 4'h3 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_9 : _exe_ctrl_pc_sel_T_26;
  wire [1:0] _exe_ctrl_pc_sel_T_30 = 4'h4 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_12 : _exe_ctrl_pc_sel_T_28;
  wire [1:0] _exe_ctrl_pc_sel_T_32 = 4'h5 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_14 : _exe_ctrl_pc_sel_T_30;
  wire [1:0] _exe_ctrl_pc_sel_T_34 = 4'h6 == io_in_bits_br_type ? _exe_ctrl_pc_sel_T_16 : _exe_ctrl_pc_sel_T_32;
  wire [1:0] _exe_ctrl_pc_sel_T_36 = 4'h7 == io_in_bits_br_type ? 2'h1 : _exe_ctrl_pc_sel_T_34;
  wire [1:0] _exe_ctrl_pc_sel_T_38 = 4'h8 == io_in_bits_br_type ? 2'h2 : _exe_ctrl_pc_sel_T_36;
  wire [1:0] _exe_ctrl_pc_sel_T_40 = 4'h9 == io_in_bits_br_type ? 2'h1 : _exe_ctrl_pc_sel_T_38;
  wire [1:0] exe_ctrl_pc_sel = 4'ha == io_in_bits_br_type ? 2'h2 : _exe_ctrl_pc_sel_T_40;
  wire [31:0] _io_out_bits_redirect_target_T_2 = io_in_bits_pc + 32'h4;
  wire [63:0] _io_out_bits_redirect_target_T_4 = io_in_bits_op1_data + io_in_bits_op2_data;
  wire [63:0] _io_out_bits_redirect_target_T_5 = exe_ctrl_pc_sel == 2'h3 ? {{32'd0}, _io_out_bits_redirect_target_T_2}
     : _io_out_bits_redirect_target_T_4;
  assign io_out_bits_redirect_valid = io_in_valid & io_out_bits_redirect_target != _io_out_bits_redirect_target_T_2;
  assign io_out_bits_redirect_target = _io_out_bits_redirect_target_T_5[31:0];
endmodule
module ysyx_040656_ExternalMul(
  input          clock,
  input          reset,
  input          io_in_valid,
  input  [63:0]  io_in_bits_op1,
  input  [63:0]  io_in_bits_op2,
  input  [5:0]   io_in_bits_func,
  output         io_out_valid,
  output [127:0] io_out_bits_dataout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
`endif
  wire  mul1_clock;
  wire  mul1_reset;
  wire  mul1_sign;
  wire [31:0] mul1_x;
  wire [31:0] mul1_y;
  wire [63:0] mul1_result;
  wire  mul2_clock;
  wire  mul2_reset;
  wire  mul2_sign;
  wire [31:0] mul2_x;
  wire [31:0] mul2_y;
  wire [63:0] mul2_result;
  wire  mul3_clock;
  wire  mul3_reset;
  wire  mul3_sign;
  wire [31:0] mul3_x;
  wire [31:0] mul3_y;
  wire [63:0] mul3_result;
  wire  mul4_clock;
  wire  mul4_reset;
  wire  mul4_sign;
  wire [31:0] mul4_x;
  wire [31:0] mul4_y;
  wire [63:0] mul4_result;
  wire  xIsNegative = io_in_bits_op1[63];
  wire  yIsNegative = io_in_bits_op2[63];
  reg [1:0] state;
  reg  valid;
  reg [127:0] dataout;
  wire  _T = io_in_bits_func == 6'h1e;
  wire  _T_1 = xIsNegative ^ yIsNegative;
  wire [63:0] _x_T_4 = 64'sh0 - $signed(io_in_bits_op1);
  wire [63:0] _GEN_0 = xIsNegative ? _x_T_4 : io_in_bits_op1;
  wire [63:0] _GEN_2 = xIsNegative & yIsNegative ? _x_T_4 : io_in_bits_op1;
  wire [63:0] _GEN_4 = xIsNegative ^ yIsNegative ? _GEN_0 : _GEN_2;
  wire  _T_3 = io_in_bits_func == 6'h1f;
  wire [63:0] _GEN_8 = io_in_bits_func == 6'h1f ? _GEN_0 : io_in_bits_op1;
  wire [63:0] x = io_in_bits_func == 6'h1e ? _GEN_4 : _GEN_8;
  wire [63:0] _y_T_4 = 64'sh0 - $signed(io_in_bits_op2);
  wire [63:0] _GEN_1 = xIsNegative ? io_in_bits_op2 : _y_T_4;
  wire [63:0] _GEN_3 = xIsNegative & yIsNegative ? _y_T_4 : io_in_bits_op2;
  wire [63:0] _GEN_5 = xIsNegative ^ yIsNegative ? _GEN_1 : _GEN_3;
  wire [63:0] y = io_in_bits_func == 6'h1e ? _GEN_5 : io_in_bits_op2;
  wire [127:0] _result_T = {64'h0,mul1_result};
  wire [127:0] _result_T_2 = {64'h0,mul2_result};
  wire [159:0] _result_T_3 = {_result_T_2, 32'h0};
  wire [127:0] _result_T_6 = _result_T + _result_T_3[127:0];
  wire [127:0] _result_T_7 = {64'h0,mul3_result};
  wire [159:0] _result_T_8 = {_result_T_7, 32'h0};
  wire [127:0] _result_T_11 = _result_T_6 + _result_T_8[127:0];
  wire [127:0] _result_T_12 = {64'h0,mul4_result};
  wire [191:0] _result_T_13 = {_result_T_12, 64'h0};
  wire [127:0] result = _result_T_11 + _result_T_13[127:0];
  wire [127:0] _dataout_T = _result_T_11 + _result_T_13[127:0];
  wire [127:0] _dataout_T_4 = 128'sh0 - $signed(_dataout_T);
  wire [127:0] _GEN_14 = _T_1 ? _dataout_T_4 : result;
  wire  dataout_signBit = result[31];
  wire [95:0] _dataout_T_7 = dataout_signBit ? 96'hffffffffffffffffffffffff : 96'h0;
  wire [127:0] _dataout_T_8 = {_dataout_T_7,result[31:0]};
  wire [127:0] _GEN_15 = xIsNegative ? _dataout_T_4 : result;
  wire [127:0] _GEN_16 = _T_3 ? _GEN_15 : result;
  wire [127:0] _GEN_17 = io_in_bits_func == 6'h25 ? _dataout_T_8 : _GEN_16;
  wire [127:0] _GEN_18 = _T ? _GEN_14 : _GEN_17;
  wire [1:0] _GEN_22 = 2'h3 == state ? 2'h0 : state;
  wire  _GEN_24 = 2'h3 == state ? 1'h0 : valid;
  wire  _GEN_27 = 2'h2 == state | _GEN_24;
  ysyx_040656_mul_mul mul1 (
    .clock(mul1_clock),
    .reset(mul1_reset),
    .sign(mul1_sign),
    .x(mul1_x),
    .y(mul1_y),
    .result(mul1_result)
  );
  ysyx_040656_mul_mul mul2 (
    .clock(mul2_clock),
    .reset(mul2_reset),
    .sign(mul2_sign),
    .x(mul2_x),
    .y(mul2_y),
    .result(mul2_result)
  );
  ysyx_040656_mul_mul mul3 (
    .clock(mul3_clock),
    .reset(mul3_reset),
    .sign(mul3_sign),
    .x(mul3_x),
    .y(mul3_y),
    .result(mul3_result)
  );
  ysyx_040656_mul_mul mul4 (
    .clock(mul4_clock),
    .reset(mul4_reset),
    .sign(mul4_sign),
    .x(mul4_x),
    .y(mul4_y),
    .result(mul4_result)
  );
  assign io_out_valid = valid;
  assign io_out_bits_dataout = dataout;
  assign mul1_clock = clock;
  assign mul1_reset = reset;
  assign mul1_sign = 1'h0;
  assign mul1_x = x[31:0];
  assign mul1_y = y[31:0];
  assign mul2_clock = clock;
  assign mul2_reset = reset;
  assign mul2_sign = 1'h0;
  assign mul2_x = x[31:0];
  assign mul2_y = y[63:32];
  assign mul3_clock = clock;
  assign mul3_reset = reset;
  assign mul3_sign = 1'h0;
  assign mul3_x = x[63:32];
  assign mul3_y = y[31:0];
  assign mul4_clock = clock;
  assign mul4_reset = reset;
  assign mul4_sign = 1'h0;
  assign mul4_x = x[63:32];
  assign mul4_y = y[63:32];
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (2'h0 == state) begin
      if (io_in_valid) begin
        state <= 2'h1;
      end
    end else if (2'h1 == state) begin
      state <= 2'h2;
    end else if (2'h2 == state) begin
      state <= 2'h3;
    end else begin
      state <= _GEN_22;
    end
    if (reset) begin
      valid <= 1'h0;
    end else if (2'h0 == state) begin
      valid <= 1'h0;
    end else if (!(2'h1 == state)) begin
      valid <= _GEN_27;
    end
    if (reset) begin
      dataout <= 128'h0;
    end else if (2'h0 == state) begin
      dataout <= 128'h0;
    end else if (!(2'h1 == state)) begin
      if (2'h2 == state) begin
        dataout <= _GEN_18;
      end
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  valid = _RAND_1[0:0];
  _RAND_2 = {4{`RANDOM}};
  dataout = _RAND_2[127:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_ExternalDiv(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_sign,
  input  [63:0] io_in_bits_x,
  input  [63:0] io_in_bits_y,
  input  [5:0]  io_in_bits_func,
  output        io_out_valid,
  output [63:0] io_out_bits_s,
  output [63:0] io_out_bits_r
);
  wire  div_clock;
  wire  div_reset;
  wire  div_valid;
  wire  div_sign;
  wire [63:0] div_x;
  wire [63:0] div_y;
  wire [63:0] div_s;
  wire [63:0] div_r;
  wire  div_ready;
  wire  div_out_valid;
  wire  div_out_ready;
  wire  _div_io_x_T = io_in_bits_y == 64'h0;
  wire [63:0] _div_io_x_T_1 = io_in_bits_y == 64'h0 ? 64'hfadefade : io_in_bits_x;
  wire [63:0] _div_io_y_T_1 = _div_io_x_T ? 64'hfadefade : io_in_bits_y;
  wire [63:0] _io_out_bits_s_T_2 = _div_io_x_T ? 64'hffffffffffffffff : div_s;
  wire [63:0] _io_out_bits_r_T_5 = io_in_bits_x - 64'h2;
  wire [63:0] _io_out_bits_r_T_9 = 6'h29 == io_in_bits_func ? io_in_bits_x : 64'h0;
  wire [63:0] _io_out_bits_r_T_11 = 6'h28 == io_in_bits_func ? _io_out_bits_r_T_5 : _io_out_bits_r_T_9;
  wire [63:0] _io_out_bits_r_T_13 = 6'h23 == io_in_bits_func ? io_in_bits_x : _io_out_bits_r_T_11;
  wire [63:0] _io_out_bits_r_T_15 = 6'h24 == io_in_bits_func ? io_in_bits_x : _io_out_bits_r_T_13;
  wire [63:0] _io_out_bits_r_T_16 = _div_io_x_T ? _io_out_bits_r_T_15 : div_r;
  ysyx_040656_div_div div (
    .clock(div_clock),
    .reset(div_reset),
    .valid(div_valid),
    .sign(div_sign),
    .x(div_x),
    .y(div_y),
    .s(div_s),
    .r(div_r),
    .ready(div_ready),
    .out_valid(div_out_valid),
    .out_ready(div_out_ready)
  );
  assign io_out_valid = div_out_valid;
  assign io_out_bits_s = io_in_valid ? _io_out_bits_s_T_2 : 64'h0;
  assign io_out_bits_r = io_in_valid ? _io_out_bits_r_T_16 : 64'h0;
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_valid = io_in_valid;
  assign div_sign = io_in_valid & io_in_bits_sign;
  assign div_x = io_in_valid ? _div_io_x_T_1 : 64'h0;
  assign div_y = io_in_valid ? _div_io_y_T_1 : 64'h1;
  assign div_out_ready = 1'h1;
endmodule
module ysyx_040656_FastDivShift(
  input  [63:0] io_in_op1_data,
  input  [63:0] io_in_op2_data,
  output [63:0] io_out_r,
  output [63:0] io_out_s
);
  wire [31:0] io_out_s_hi = io_in_op2_data[63:32];
  wire [31:0] io_out_s_lo = io_in_op2_data[31:0];
  wire  io_out_s_useHi = |io_out_s_hi;
  wire [15:0] io_out_s_hi_1 = io_out_s_hi[31:16];
  wire [15:0] io_out_s_lo_1 = io_out_s_hi[15:0];
  wire  io_out_s_useHi_1 = |io_out_s_hi_1;
  wire [7:0] io_out_s_hi_2 = io_out_s_hi_1[15:8];
  wire [7:0] io_out_s_lo_2 = io_out_s_hi_1[7:0];
  wire  io_out_s_useHi_2 = |io_out_s_hi_2;
  wire [3:0] io_out_s_hi_3 = io_out_s_hi_2[7:4];
  wire [3:0] io_out_s_lo_3 = io_out_s_hi_2[3:0];
  wire  io_out_s_useHi_3 = |io_out_s_hi_3;
  wire [1:0] _io_out_s_T_3 = io_out_s_hi_3[2] ? 2'h2 : {{1'd0}, io_out_s_hi_3[1]};
  wire [1:0] _io_out_s_T_4 = io_out_s_hi_3[3] ? 2'h3 : _io_out_s_T_3;
  wire [1:0] _io_out_s_T_8 = io_out_s_lo_3[2] ? 2'h2 : {{1'd0}, io_out_s_lo_3[1]};
  wire [1:0] _io_out_s_T_9 = io_out_s_lo_3[3] ? 2'h3 : _io_out_s_T_8;
  wire [1:0] _io_out_s_T_10 = io_out_s_useHi_3 ? _io_out_s_T_4 : _io_out_s_T_9;
  wire [2:0] _io_out_s_T_11 = {io_out_s_useHi_3,_io_out_s_T_10};
  wire [3:0] io_out_s_hi_4 = io_out_s_lo_2[7:4];
  wire [3:0] io_out_s_lo_4 = io_out_s_lo_2[3:0];
  wire  io_out_s_useHi_4 = |io_out_s_hi_4;
  wire [1:0] _io_out_s_T_15 = io_out_s_hi_4[2] ? 2'h2 : {{1'd0}, io_out_s_hi_4[1]};
  wire [1:0] _io_out_s_T_16 = io_out_s_hi_4[3] ? 2'h3 : _io_out_s_T_15;
  wire [1:0] _io_out_s_T_20 = io_out_s_lo_4[2] ? 2'h2 : {{1'd0}, io_out_s_lo_4[1]};
  wire [1:0] _io_out_s_T_21 = io_out_s_lo_4[3] ? 2'h3 : _io_out_s_T_20;
  wire [1:0] _io_out_s_T_22 = io_out_s_useHi_4 ? _io_out_s_T_16 : _io_out_s_T_21;
  wire [2:0] _io_out_s_T_23 = {io_out_s_useHi_4,_io_out_s_T_22};
  wire [2:0] _io_out_s_T_24 = io_out_s_useHi_2 ? _io_out_s_T_11 : _io_out_s_T_23;
  wire [3:0] _io_out_s_T_25 = {io_out_s_useHi_2,_io_out_s_T_24};
  wire [7:0] io_out_s_hi_5 = io_out_s_lo_1[15:8];
  wire [7:0] io_out_s_lo_5 = io_out_s_lo_1[7:0];
  wire  io_out_s_useHi_5 = |io_out_s_hi_5;
  wire [3:0] io_out_s_hi_6 = io_out_s_hi_5[7:4];
  wire [3:0] io_out_s_lo_6 = io_out_s_hi_5[3:0];
  wire  io_out_s_useHi_6 = |io_out_s_hi_6;
  wire [1:0] _io_out_s_T_29 = io_out_s_hi_6[2] ? 2'h2 : {{1'd0}, io_out_s_hi_6[1]};
  wire [1:0] _io_out_s_T_30 = io_out_s_hi_6[3] ? 2'h3 : _io_out_s_T_29;
  wire [1:0] _io_out_s_T_34 = io_out_s_lo_6[2] ? 2'h2 : {{1'd0}, io_out_s_lo_6[1]};
  wire [1:0] _io_out_s_T_35 = io_out_s_lo_6[3] ? 2'h3 : _io_out_s_T_34;
  wire [1:0] _io_out_s_T_36 = io_out_s_useHi_6 ? _io_out_s_T_30 : _io_out_s_T_35;
  wire [2:0] _io_out_s_T_37 = {io_out_s_useHi_6,_io_out_s_T_36};
  wire [3:0] io_out_s_hi_7 = io_out_s_lo_5[7:4];
  wire [3:0] io_out_s_lo_7 = io_out_s_lo_5[3:0];
  wire  io_out_s_useHi_7 = |io_out_s_hi_7;
  wire [1:0] _io_out_s_T_41 = io_out_s_hi_7[2] ? 2'h2 : {{1'd0}, io_out_s_hi_7[1]};
  wire [1:0] _io_out_s_T_42 = io_out_s_hi_7[3] ? 2'h3 : _io_out_s_T_41;
  wire [1:0] _io_out_s_T_46 = io_out_s_lo_7[2] ? 2'h2 : {{1'd0}, io_out_s_lo_7[1]};
  wire [1:0] _io_out_s_T_47 = io_out_s_lo_7[3] ? 2'h3 : _io_out_s_T_46;
  wire [1:0] _io_out_s_T_48 = io_out_s_useHi_7 ? _io_out_s_T_42 : _io_out_s_T_47;
  wire [2:0] _io_out_s_T_49 = {io_out_s_useHi_7,_io_out_s_T_48};
  wire [2:0] _io_out_s_T_50 = io_out_s_useHi_5 ? _io_out_s_T_37 : _io_out_s_T_49;
  wire [3:0] _io_out_s_T_51 = {io_out_s_useHi_5,_io_out_s_T_50};
  wire [3:0] _io_out_s_T_52 = io_out_s_useHi_1 ? _io_out_s_T_25 : _io_out_s_T_51;
  wire [4:0] _io_out_s_T_53 = {io_out_s_useHi_1,_io_out_s_T_52};
  wire [15:0] io_out_s_hi_8 = io_out_s_lo[31:16];
  wire [15:0] io_out_s_lo_8 = io_out_s_lo[15:0];
  wire  io_out_s_useHi_8 = |io_out_s_hi_8;
  wire [7:0] io_out_s_hi_9 = io_out_s_hi_8[15:8];
  wire [7:0] io_out_s_lo_9 = io_out_s_hi_8[7:0];
  wire  io_out_s_useHi_9 = |io_out_s_hi_9;
  wire [3:0] io_out_s_hi_10 = io_out_s_hi_9[7:4];
  wire [3:0] io_out_s_lo_10 = io_out_s_hi_9[3:0];
  wire  io_out_s_useHi_10 = |io_out_s_hi_10;
  wire [1:0] _io_out_s_T_57 = io_out_s_hi_10[2] ? 2'h2 : {{1'd0}, io_out_s_hi_10[1]};
  wire [1:0] _io_out_s_T_58 = io_out_s_hi_10[3] ? 2'h3 : _io_out_s_T_57;
  wire [1:0] _io_out_s_T_62 = io_out_s_lo_10[2] ? 2'h2 : {{1'd0}, io_out_s_lo_10[1]};
  wire [1:0] _io_out_s_T_63 = io_out_s_lo_10[3] ? 2'h3 : _io_out_s_T_62;
  wire [1:0] _io_out_s_T_64 = io_out_s_useHi_10 ? _io_out_s_T_58 : _io_out_s_T_63;
  wire [2:0] _io_out_s_T_65 = {io_out_s_useHi_10,_io_out_s_T_64};
  wire [3:0] io_out_s_hi_11 = io_out_s_lo_9[7:4];
  wire [3:0] io_out_s_lo_11 = io_out_s_lo_9[3:0];
  wire  io_out_s_useHi_11 = |io_out_s_hi_11;
  wire [1:0] _io_out_s_T_69 = io_out_s_hi_11[2] ? 2'h2 : {{1'd0}, io_out_s_hi_11[1]};
  wire [1:0] _io_out_s_T_70 = io_out_s_hi_11[3] ? 2'h3 : _io_out_s_T_69;
  wire [1:0] _io_out_s_T_74 = io_out_s_lo_11[2] ? 2'h2 : {{1'd0}, io_out_s_lo_11[1]};
  wire [1:0] _io_out_s_T_75 = io_out_s_lo_11[3] ? 2'h3 : _io_out_s_T_74;
  wire [1:0] _io_out_s_T_76 = io_out_s_useHi_11 ? _io_out_s_T_70 : _io_out_s_T_75;
  wire [2:0] _io_out_s_T_77 = {io_out_s_useHi_11,_io_out_s_T_76};
  wire [2:0] _io_out_s_T_78 = io_out_s_useHi_9 ? _io_out_s_T_65 : _io_out_s_T_77;
  wire [3:0] _io_out_s_T_79 = {io_out_s_useHi_9,_io_out_s_T_78};
  wire [7:0] io_out_s_hi_12 = io_out_s_lo_8[15:8];
  wire [7:0] io_out_s_lo_12 = io_out_s_lo_8[7:0];
  wire  io_out_s_useHi_12 = |io_out_s_hi_12;
  wire [3:0] io_out_s_hi_13 = io_out_s_hi_12[7:4];
  wire [3:0] io_out_s_lo_13 = io_out_s_hi_12[3:0];
  wire  io_out_s_useHi_13 = |io_out_s_hi_13;
  wire [1:0] _io_out_s_T_83 = io_out_s_hi_13[2] ? 2'h2 : {{1'd0}, io_out_s_hi_13[1]};
  wire [1:0] _io_out_s_T_84 = io_out_s_hi_13[3] ? 2'h3 : _io_out_s_T_83;
  wire [1:0] _io_out_s_T_88 = io_out_s_lo_13[2] ? 2'h2 : {{1'd0}, io_out_s_lo_13[1]};
  wire [1:0] _io_out_s_T_89 = io_out_s_lo_13[3] ? 2'h3 : _io_out_s_T_88;
  wire [1:0] _io_out_s_T_90 = io_out_s_useHi_13 ? _io_out_s_T_84 : _io_out_s_T_89;
  wire [2:0] _io_out_s_T_91 = {io_out_s_useHi_13,_io_out_s_T_90};
  wire [3:0] io_out_s_hi_14 = io_out_s_lo_12[7:4];
  wire [3:0] io_out_s_lo_14 = io_out_s_lo_12[3:0];
  wire  io_out_s_useHi_14 = |io_out_s_hi_14;
  wire [1:0] _io_out_s_T_95 = io_out_s_hi_14[2] ? 2'h2 : {{1'd0}, io_out_s_hi_14[1]};
  wire [1:0] _io_out_s_T_96 = io_out_s_hi_14[3] ? 2'h3 : _io_out_s_T_95;
  wire [1:0] _io_out_s_T_100 = io_out_s_lo_14[2] ? 2'h2 : {{1'd0}, io_out_s_lo_14[1]};
  wire [1:0] _io_out_s_T_101 = io_out_s_lo_14[3] ? 2'h3 : _io_out_s_T_100;
  wire [1:0] _io_out_s_T_102 = io_out_s_useHi_14 ? _io_out_s_T_96 : _io_out_s_T_101;
  wire [2:0] _io_out_s_T_103 = {io_out_s_useHi_14,_io_out_s_T_102};
  wire [2:0] _io_out_s_T_104 = io_out_s_useHi_12 ? _io_out_s_T_91 : _io_out_s_T_103;
  wire [3:0] _io_out_s_T_105 = {io_out_s_useHi_12,_io_out_s_T_104};
  wire [3:0] _io_out_s_T_106 = io_out_s_useHi_8 ? _io_out_s_T_79 : _io_out_s_T_105;
  wire [4:0] _io_out_s_T_107 = {io_out_s_useHi_8,_io_out_s_T_106};
  wire [4:0] _io_out_s_T_108 = io_out_s_useHi ? _io_out_s_T_53 : _io_out_s_T_107;
  wire [5:0] _io_out_s_T_109 = {io_out_s_useHi,_io_out_s_T_108};
  wire [63:0] _io_out_r_T_1 = io_in_op2_data - 64'h1;
  assign io_out_r = io_in_op1_data & _io_out_r_T_1;
  assign io_out_s = io_in_op1_data >> _io_out_s_T_109;
endmodule
module ysyx_040656_FastDiv(
  input  [63:0] io_in_op1_data,
  input  [63:0] io_in_op2_data,
  input         io_in_valid,
  input         io_in_isPow,
  output [63:0] io_out_r,
  output [63:0] io_out_s,
  output        io_out_valid
);
  wire [63:0] fastDivShift_io_in_op1_data;
  wire [63:0] fastDivShift_io_in_op2_data;
  wire [63:0] fastDivShift_io_out_r;
  wire [63:0] fastDivShift_io_out_s;
  wire [13:0] index = {io_in_op1_data[6:0],io_in_op2_data[6:0]};
  wire [13:0] _GEN_129 = 14'h81 == index ? 14'h80 : 14'h0;
  wire [13:0] _GEN_130 = 14'h82 == index ? 14'h1 : _GEN_129;
  wire [13:0] _GEN_131 = 14'h83 == index ? 14'h1 : _GEN_130;
  wire [13:0] _GEN_132 = 14'h84 == index ? 14'h1 : _GEN_131;
  wire [13:0] _GEN_133 = 14'h85 == index ? 14'h1 : _GEN_132;
  wire [13:0] _GEN_134 = 14'h86 == index ? 14'h1 : _GEN_133;
  wire [13:0] _GEN_135 = 14'h87 == index ? 14'h1 : _GEN_134;
  wire [13:0] _GEN_136 = 14'h88 == index ? 14'h1 : _GEN_135;
  wire [13:0] _GEN_137 = 14'h89 == index ? 14'h1 : _GEN_136;
  wire [13:0] _GEN_138 = 14'h8a == index ? 14'h1 : _GEN_137;
  wire [13:0] _GEN_139 = 14'h8b == index ? 14'h1 : _GEN_138;
  wire [13:0] _GEN_140 = 14'h8c == index ? 14'h1 : _GEN_139;
  wire [13:0] _GEN_141 = 14'h8d == index ? 14'h1 : _GEN_140;
  wire [13:0] _GEN_142 = 14'h8e == index ? 14'h1 : _GEN_141;
  wire [13:0] _GEN_143 = 14'h8f == index ? 14'h1 : _GEN_142;
  wire [13:0] _GEN_144 = 14'h90 == index ? 14'h1 : _GEN_143;
  wire [13:0] _GEN_145 = 14'h91 == index ? 14'h1 : _GEN_144;
  wire [13:0] _GEN_146 = 14'h92 == index ? 14'h1 : _GEN_145;
  wire [13:0] _GEN_147 = 14'h93 == index ? 14'h1 : _GEN_146;
  wire [13:0] _GEN_148 = 14'h94 == index ? 14'h1 : _GEN_147;
  wire [13:0] _GEN_149 = 14'h95 == index ? 14'h1 : _GEN_148;
  wire [13:0] _GEN_150 = 14'h96 == index ? 14'h1 : _GEN_149;
  wire [13:0] _GEN_151 = 14'h97 == index ? 14'h1 : _GEN_150;
  wire [13:0] _GEN_152 = 14'h98 == index ? 14'h1 : _GEN_151;
  wire [13:0] _GEN_153 = 14'h99 == index ? 14'h1 : _GEN_152;
  wire [13:0] _GEN_154 = 14'h9a == index ? 14'h1 : _GEN_153;
  wire [13:0] _GEN_155 = 14'h9b == index ? 14'h1 : _GEN_154;
  wire [13:0] _GEN_156 = 14'h9c == index ? 14'h1 : _GEN_155;
  wire [13:0] _GEN_157 = 14'h9d == index ? 14'h1 : _GEN_156;
  wire [13:0] _GEN_158 = 14'h9e == index ? 14'h1 : _GEN_157;
  wire [13:0] _GEN_159 = 14'h9f == index ? 14'h1 : _GEN_158;
  wire [13:0] _GEN_160 = 14'ha0 == index ? 14'h1 : _GEN_159;
  wire [13:0] _GEN_161 = 14'ha1 == index ? 14'h1 : _GEN_160;
  wire [13:0] _GEN_162 = 14'ha2 == index ? 14'h1 : _GEN_161;
  wire [13:0] _GEN_163 = 14'ha3 == index ? 14'h1 : _GEN_162;
  wire [13:0] _GEN_164 = 14'ha4 == index ? 14'h1 : _GEN_163;
  wire [13:0] _GEN_165 = 14'ha5 == index ? 14'h1 : _GEN_164;
  wire [13:0] _GEN_166 = 14'ha6 == index ? 14'h1 : _GEN_165;
  wire [13:0] _GEN_167 = 14'ha7 == index ? 14'h1 : _GEN_166;
  wire [13:0] _GEN_168 = 14'ha8 == index ? 14'h1 : _GEN_167;
  wire [13:0] _GEN_169 = 14'ha9 == index ? 14'h1 : _GEN_168;
  wire [13:0] _GEN_170 = 14'haa == index ? 14'h1 : _GEN_169;
  wire [13:0] _GEN_171 = 14'hab == index ? 14'h1 : _GEN_170;
  wire [13:0] _GEN_172 = 14'hac == index ? 14'h1 : _GEN_171;
  wire [13:0] _GEN_173 = 14'had == index ? 14'h1 : _GEN_172;
  wire [13:0] _GEN_174 = 14'hae == index ? 14'h1 : _GEN_173;
  wire [13:0] _GEN_175 = 14'haf == index ? 14'h1 : _GEN_174;
  wire [13:0] _GEN_176 = 14'hb0 == index ? 14'h1 : _GEN_175;
  wire [13:0] _GEN_177 = 14'hb1 == index ? 14'h1 : _GEN_176;
  wire [13:0] _GEN_178 = 14'hb2 == index ? 14'h1 : _GEN_177;
  wire [13:0] _GEN_179 = 14'hb3 == index ? 14'h1 : _GEN_178;
  wire [13:0] _GEN_180 = 14'hb4 == index ? 14'h1 : _GEN_179;
  wire [13:0] _GEN_181 = 14'hb5 == index ? 14'h1 : _GEN_180;
  wire [13:0] _GEN_182 = 14'hb6 == index ? 14'h1 : _GEN_181;
  wire [13:0] _GEN_183 = 14'hb7 == index ? 14'h1 : _GEN_182;
  wire [13:0] _GEN_184 = 14'hb8 == index ? 14'h1 : _GEN_183;
  wire [13:0] _GEN_185 = 14'hb9 == index ? 14'h1 : _GEN_184;
  wire [13:0] _GEN_186 = 14'hba == index ? 14'h1 : _GEN_185;
  wire [13:0] _GEN_187 = 14'hbb == index ? 14'h1 : _GEN_186;
  wire [13:0] _GEN_188 = 14'hbc == index ? 14'h1 : _GEN_187;
  wire [13:0] _GEN_189 = 14'hbd == index ? 14'h1 : _GEN_188;
  wire [13:0] _GEN_190 = 14'hbe == index ? 14'h1 : _GEN_189;
  wire [13:0] _GEN_191 = 14'hbf == index ? 14'h1 : _GEN_190;
  wire [13:0] _GEN_192 = 14'hc0 == index ? 14'h1 : _GEN_191;
  wire [13:0] _GEN_193 = 14'hc1 == index ? 14'h1 : _GEN_192;
  wire [13:0] _GEN_194 = 14'hc2 == index ? 14'h1 : _GEN_193;
  wire [13:0] _GEN_195 = 14'hc3 == index ? 14'h1 : _GEN_194;
  wire [13:0] _GEN_196 = 14'hc4 == index ? 14'h1 : _GEN_195;
  wire [13:0] _GEN_197 = 14'hc5 == index ? 14'h1 : _GEN_196;
  wire [13:0] _GEN_198 = 14'hc6 == index ? 14'h1 : _GEN_197;
  wire [13:0] _GEN_199 = 14'hc7 == index ? 14'h1 : _GEN_198;
  wire [13:0] _GEN_200 = 14'hc8 == index ? 14'h1 : _GEN_199;
  wire [13:0] _GEN_201 = 14'hc9 == index ? 14'h1 : _GEN_200;
  wire [13:0] _GEN_202 = 14'hca == index ? 14'h1 : _GEN_201;
  wire [13:0] _GEN_203 = 14'hcb == index ? 14'h1 : _GEN_202;
  wire [13:0] _GEN_204 = 14'hcc == index ? 14'h1 : _GEN_203;
  wire [13:0] _GEN_205 = 14'hcd == index ? 14'h1 : _GEN_204;
  wire [13:0] _GEN_206 = 14'hce == index ? 14'h1 : _GEN_205;
  wire [13:0] _GEN_207 = 14'hcf == index ? 14'h1 : _GEN_206;
  wire [13:0] _GEN_208 = 14'hd0 == index ? 14'h1 : _GEN_207;
  wire [13:0] _GEN_209 = 14'hd1 == index ? 14'h1 : _GEN_208;
  wire [13:0] _GEN_210 = 14'hd2 == index ? 14'h1 : _GEN_209;
  wire [13:0] _GEN_211 = 14'hd3 == index ? 14'h1 : _GEN_210;
  wire [13:0] _GEN_212 = 14'hd4 == index ? 14'h1 : _GEN_211;
  wire [13:0] _GEN_213 = 14'hd5 == index ? 14'h1 : _GEN_212;
  wire [13:0] _GEN_214 = 14'hd6 == index ? 14'h1 : _GEN_213;
  wire [13:0] _GEN_215 = 14'hd7 == index ? 14'h1 : _GEN_214;
  wire [13:0] _GEN_216 = 14'hd8 == index ? 14'h1 : _GEN_215;
  wire [13:0] _GEN_217 = 14'hd9 == index ? 14'h1 : _GEN_216;
  wire [13:0] _GEN_218 = 14'hda == index ? 14'h1 : _GEN_217;
  wire [13:0] _GEN_219 = 14'hdb == index ? 14'h1 : _GEN_218;
  wire [13:0] _GEN_220 = 14'hdc == index ? 14'h1 : _GEN_219;
  wire [13:0] _GEN_221 = 14'hdd == index ? 14'h1 : _GEN_220;
  wire [13:0] _GEN_222 = 14'hde == index ? 14'h1 : _GEN_221;
  wire [13:0] _GEN_223 = 14'hdf == index ? 14'h1 : _GEN_222;
  wire [13:0] _GEN_224 = 14'he0 == index ? 14'h1 : _GEN_223;
  wire [13:0] _GEN_225 = 14'he1 == index ? 14'h1 : _GEN_224;
  wire [13:0] _GEN_226 = 14'he2 == index ? 14'h1 : _GEN_225;
  wire [13:0] _GEN_227 = 14'he3 == index ? 14'h1 : _GEN_226;
  wire [13:0] _GEN_228 = 14'he4 == index ? 14'h1 : _GEN_227;
  wire [13:0] _GEN_229 = 14'he5 == index ? 14'h1 : _GEN_228;
  wire [13:0] _GEN_230 = 14'he6 == index ? 14'h1 : _GEN_229;
  wire [13:0] _GEN_231 = 14'he7 == index ? 14'h1 : _GEN_230;
  wire [13:0] _GEN_232 = 14'he8 == index ? 14'h1 : _GEN_231;
  wire [13:0] _GEN_233 = 14'he9 == index ? 14'h1 : _GEN_232;
  wire [13:0] _GEN_234 = 14'hea == index ? 14'h1 : _GEN_233;
  wire [13:0] _GEN_235 = 14'heb == index ? 14'h1 : _GEN_234;
  wire [13:0] _GEN_236 = 14'hec == index ? 14'h1 : _GEN_235;
  wire [13:0] _GEN_237 = 14'hed == index ? 14'h1 : _GEN_236;
  wire [13:0] _GEN_238 = 14'hee == index ? 14'h1 : _GEN_237;
  wire [13:0] _GEN_239 = 14'hef == index ? 14'h1 : _GEN_238;
  wire [13:0] _GEN_240 = 14'hf0 == index ? 14'h1 : _GEN_239;
  wire [13:0] _GEN_241 = 14'hf1 == index ? 14'h1 : _GEN_240;
  wire [13:0] _GEN_242 = 14'hf2 == index ? 14'h1 : _GEN_241;
  wire [13:0] _GEN_243 = 14'hf3 == index ? 14'h1 : _GEN_242;
  wire [13:0] _GEN_244 = 14'hf4 == index ? 14'h1 : _GEN_243;
  wire [13:0] _GEN_245 = 14'hf5 == index ? 14'h1 : _GEN_244;
  wire [13:0] _GEN_246 = 14'hf6 == index ? 14'h1 : _GEN_245;
  wire [13:0] _GEN_247 = 14'hf7 == index ? 14'h1 : _GEN_246;
  wire [13:0] _GEN_248 = 14'hf8 == index ? 14'h1 : _GEN_247;
  wire [13:0] _GEN_249 = 14'hf9 == index ? 14'h1 : _GEN_248;
  wire [13:0] _GEN_250 = 14'hfa == index ? 14'h1 : _GEN_249;
  wire [13:0] _GEN_251 = 14'hfb == index ? 14'h1 : _GEN_250;
  wire [13:0] _GEN_252 = 14'hfc == index ? 14'h1 : _GEN_251;
  wire [13:0] _GEN_253 = 14'hfd == index ? 14'h1 : _GEN_252;
  wire [13:0] _GEN_254 = 14'hfe == index ? 14'h1 : _GEN_253;
  wire [13:0] _GEN_255 = 14'hff == index ? 14'h1 : _GEN_254;
  wire [13:0] _GEN_256 = 14'h100 == index ? 14'h0 : _GEN_255;
  wire [13:0] _GEN_257 = 14'h101 == index ? 14'h100 : _GEN_256;
  wire [13:0] _GEN_258 = 14'h102 == index ? 14'h80 : _GEN_257;
  wire [13:0] _GEN_259 = 14'h103 == index ? 14'h2 : _GEN_258;
  wire [13:0] _GEN_260 = 14'h104 == index ? 14'h2 : _GEN_259;
  wire [13:0] _GEN_261 = 14'h105 == index ? 14'h2 : _GEN_260;
  wire [13:0] _GEN_262 = 14'h106 == index ? 14'h2 : _GEN_261;
  wire [13:0] _GEN_263 = 14'h107 == index ? 14'h2 : _GEN_262;
  wire [13:0] _GEN_264 = 14'h108 == index ? 14'h2 : _GEN_263;
  wire [13:0] _GEN_265 = 14'h109 == index ? 14'h2 : _GEN_264;
  wire [13:0] _GEN_266 = 14'h10a == index ? 14'h2 : _GEN_265;
  wire [13:0] _GEN_267 = 14'h10b == index ? 14'h2 : _GEN_266;
  wire [13:0] _GEN_268 = 14'h10c == index ? 14'h2 : _GEN_267;
  wire [13:0] _GEN_269 = 14'h10d == index ? 14'h2 : _GEN_268;
  wire [13:0] _GEN_270 = 14'h10e == index ? 14'h2 : _GEN_269;
  wire [13:0] _GEN_271 = 14'h10f == index ? 14'h2 : _GEN_270;
  wire [13:0] _GEN_272 = 14'h110 == index ? 14'h2 : _GEN_271;
  wire [13:0] _GEN_273 = 14'h111 == index ? 14'h2 : _GEN_272;
  wire [13:0] _GEN_274 = 14'h112 == index ? 14'h2 : _GEN_273;
  wire [13:0] _GEN_275 = 14'h113 == index ? 14'h2 : _GEN_274;
  wire [13:0] _GEN_276 = 14'h114 == index ? 14'h2 : _GEN_275;
  wire [13:0] _GEN_277 = 14'h115 == index ? 14'h2 : _GEN_276;
  wire [13:0] _GEN_278 = 14'h116 == index ? 14'h2 : _GEN_277;
  wire [13:0] _GEN_279 = 14'h117 == index ? 14'h2 : _GEN_278;
  wire [13:0] _GEN_280 = 14'h118 == index ? 14'h2 : _GEN_279;
  wire [13:0] _GEN_281 = 14'h119 == index ? 14'h2 : _GEN_280;
  wire [13:0] _GEN_282 = 14'h11a == index ? 14'h2 : _GEN_281;
  wire [13:0] _GEN_283 = 14'h11b == index ? 14'h2 : _GEN_282;
  wire [13:0] _GEN_284 = 14'h11c == index ? 14'h2 : _GEN_283;
  wire [13:0] _GEN_285 = 14'h11d == index ? 14'h2 : _GEN_284;
  wire [13:0] _GEN_286 = 14'h11e == index ? 14'h2 : _GEN_285;
  wire [13:0] _GEN_287 = 14'h11f == index ? 14'h2 : _GEN_286;
  wire [13:0] _GEN_288 = 14'h120 == index ? 14'h2 : _GEN_287;
  wire [13:0] _GEN_289 = 14'h121 == index ? 14'h2 : _GEN_288;
  wire [13:0] _GEN_290 = 14'h122 == index ? 14'h2 : _GEN_289;
  wire [13:0] _GEN_291 = 14'h123 == index ? 14'h2 : _GEN_290;
  wire [13:0] _GEN_292 = 14'h124 == index ? 14'h2 : _GEN_291;
  wire [13:0] _GEN_293 = 14'h125 == index ? 14'h2 : _GEN_292;
  wire [13:0] _GEN_294 = 14'h126 == index ? 14'h2 : _GEN_293;
  wire [13:0] _GEN_295 = 14'h127 == index ? 14'h2 : _GEN_294;
  wire [13:0] _GEN_296 = 14'h128 == index ? 14'h2 : _GEN_295;
  wire [13:0] _GEN_297 = 14'h129 == index ? 14'h2 : _GEN_296;
  wire [13:0] _GEN_298 = 14'h12a == index ? 14'h2 : _GEN_297;
  wire [13:0] _GEN_299 = 14'h12b == index ? 14'h2 : _GEN_298;
  wire [13:0] _GEN_300 = 14'h12c == index ? 14'h2 : _GEN_299;
  wire [13:0] _GEN_301 = 14'h12d == index ? 14'h2 : _GEN_300;
  wire [13:0] _GEN_302 = 14'h12e == index ? 14'h2 : _GEN_301;
  wire [13:0] _GEN_303 = 14'h12f == index ? 14'h2 : _GEN_302;
  wire [13:0] _GEN_304 = 14'h130 == index ? 14'h2 : _GEN_303;
  wire [13:0] _GEN_305 = 14'h131 == index ? 14'h2 : _GEN_304;
  wire [13:0] _GEN_306 = 14'h132 == index ? 14'h2 : _GEN_305;
  wire [13:0] _GEN_307 = 14'h133 == index ? 14'h2 : _GEN_306;
  wire [13:0] _GEN_308 = 14'h134 == index ? 14'h2 : _GEN_307;
  wire [13:0] _GEN_309 = 14'h135 == index ? 14'h2 : _GEN_308;
  wire [13:0] _GEN_310 = 14'h136 == index ? 14'h2 : _GEN_309;
  wire [13:0] _GEN_311 = 14'h137 == index ? 14'h2 : _GEN_310;
  wire [13:0] _GEN_312 = 14'h138 == index ? 14'h2 : _GEN_311;
  wire [13:0] _GEN_313 = 14'h139 == index ? 14'h2 : _GEN_312;
  wire [13:0] _GEN_314 = 14'h13a == index ? 14'h2 : _GEN_313;
  wire [13:0] _GEN_315 = 14'h13b == index ? 14'h2 : _GEN_314;
  wire [13:0] _GEN_316 = 14'h13c == index ? 14'h2 : _GEN_315;
  wire [13:0] _GEN_317 = 14'h13d == index ? 14'h2 : _GEN_316;
  wire [13:0] _GEN_318 = 14'h13e == index ? 14'h2 : _GEN_317;
  wire [13:0] _GEN_319 = 14'h13f == index ? 14'h2 : _GEN_318;
  wire [13:0] _GEN_320 = 14'h140 == index ? 14'h2 : _GEN_319;
  wire [13:0] _GEN_321 = 14'h141 == index ? 14'h2 : _GEN_320;
  wire [13:0] _GEN_322 = 14'h142 == index ? 14'h2 : _GEN_321;
  wire [13:0] _GEN_323 = 14'h143 == index ? 14'h2 : _GEN_322;
  wire [13:0] _GEN_324 = 14'h144 == index ? 14'h2 : _GEN_323;
  wire [13:0] _GEN_325 = 14'h145 == index ? 14'h2 : _GEN_324;
  wire [13:0] _GEN_326 = 14'h146 == index ? 14'h2 : _GEN_325;
  wire [13:0] _GEN_327 = 14'h147 == index ? 14'h2 : _GEN_326;
  wire [13:0] _GEN_328 = 14'h148 == index ? 14'h2 : _GEN_327;
  wire [13:0] _GEN_329 = 14'h149 == index ? 14'h2 : _GEN_328;
  wire [13:0] _GEN_330 = 14'h14a == index ? 14'h2 : _GEN_329;
  wire [13:0] _GEN_331 = 14'h14b == index ? 14'h2 : _GEN_330;
  wire [13:0] _GEN_332 = 14'h14c == index ? 14'h2 : _GEN_331;
  wire [13:0] _GEN_333 = 14'h14d == index ? 14'h2 : _GEN_332;
  wire [13:0] _GEN_334 = 14'h14e == index ? 14'h2 : _GEN_333;
  wire [13:0] _GEN_335 = 14'h14f == index ? 14'h2 : _GEN_334;
  wire [13:0] _GEN_336 = 14'h150 == index ? 14'h2 : _GEN_335;
  wire [13:0] _GEN_337 = 14'h151 == index ? 14'h2 : _GEN_336;
  wire [13:0] _GEN_338 = 14'h152 == index ? 14'h2 : _GEN_337;
  wire [13:0] _GEN_339 = 14'h153 == index ? 14'h2 : _GEN_338;
  wire [13:0] _GEN_340 = 14'h154 == index ? 14'h2 : _GEN_339;
  wire [13:0] _GEN_341 = 14'h155 == index ? 14'h2 : _GEN_340;
  wire [13:0] _GEN_342 = 14'h156 == index ? 14'h2 : _GEN_341;
  wire [13:0] _GEN_343 = 14'h157 == index ? 14'h2 : _GEN_342;
  wire [13:0] _GEN_344 = 14'h158 == index ? 14'h2 : _GEN_343;
  wire [13:0] _GEN_345 = 14'h159 == index ? 14'h2 : _GEN_344;
  wire [13:0] _GEN_346 = 14'h15a == index ? 14'h2 : _GEN_345;
  wire [13:0] _GEN_347 = 14'h15b == index ? 14'h2 : _GEN_346;
  wire [13:0] _GEN_348 = 14'h15c == index ? 14'h2 : _GEN_347;
  wire [13:0] _GEN_349 = 14'h15d == index ? 14'h2 : _GEN_348;
  wire [13:0] _GEN_350 = 14'h15e == index ? 14'h2 : _GEN_349;
  wire [13:0] _GEN_351 = 14'h15f == index ? 14'h2 : _GEN_350;
  wire [13:0] _GEN_352 = 14'h160 == index ? 14'h2 : _GEN_351;
  wire [13:0] _GEN_353 = 14'h161 == index ? 14'h2 : _GEN_352;
  wire [13:0] _GEN_354 = 14'h162 == index ? 14'h2 : _GEN_353;
  wire [13:0] _GEN_355 = 14'h163 == index ? 14'h2 : _GEN_354;
  wire [13:0] _GEN_356 = 14'h164 == index ? 14'h2 : _GEN_355;
  wire [13:0] _GEN_357 = 14'h165 == index ? 14'h2 : _GEN_356;
  wire [13:0] _GEN_358 = 14'h166 == index ? 14'h2 : _GEN_357;
  wire [13:0] _GEN_359 = 14'h167 == index ? 14'h2 : _GEN_358;
  wire [13:0] _GEN_360 = 14'h168 == index ? 14'h2 : _GEN_359;
  wire [13:0] _GEN_361 = 14'h169 == index ? 14'h2 : _GEN_360;
  wire [13:0] _GEN_362 = 14'h16a == index ? 14'h2 : _GEN_361;
  wire [13:0] _GEN_363 = 14'h16b == index ? 14'h2 : _GEN_362;
  wire [13:0] _GEN_364 = 14'h16c == index ? 14'h2 : _GEN_363;
  wire [13:0] _GEN_365 = 14'h16d == index ? 14'h2 : _GEN_364;
  wire [13:0] _GEN_366 = 14'h16e == index ? 14'h2 : _GEN_365;
  wire [13:0] _GEN_367 = 14'h16f == index ? 14'h2 : _GEN_366;
  wire [13:0] _GEN_368 = 14'h170 == index ? 14'h2 : _GEN_367;
  wire [13:0] _GEN_369 = 14'h171 == index ? 14'h2 : _GEN_368;
  wire [13:0] _GEN_370 = 14'h172 == index ? 14'h2 : _GEN_369;
  wire [13:0] _GEN_371 = 14'h173 == index ? 14'h2 : _GEN_370;
  wire [13:0] _GEN_372 = 14'h174 == index ? 14'h2 : _GEN_371;
  wire [13:0] _GEN_373 = 14'h175 == index ? 14'h2 : _GEN_372;
  wire [13:0] _GEN_374 = 14'h176 == index ? 14'h2 : _GEN_373;
  wire [13:0] _GEN_375 = 14'h177 == index ? 14'h2 : _GEN_374;
  wire [13:0] _GEN_376 = 14'h178 == index ? 14'h2 : _GEN_375;
  wire [13:0] _GEN_377 = 14'h179 == index ? 14'h2 : _GEN_376;
  wire [13:0] _GEN_378 = 14'h17a == index ? 14'h2 : _GEN_377;
  wire [13:0] _GEN_379 = 14'h17b == index ? 14'h2 : _GEN_378;
  wire [13:0] _GEN_380 = 14'h17c == index ? 14'h2 : _GEN_379;
  wire [13:0] _GEN_381 = 14'h17d == index ? 14'h2 : _GEN_380;
  wire [13:0] _GEN_382 = 14'h17e == index ? 14'h2 : _GEN_381;
  wire [13:0] _GEN_383 = 14'h17f == index ? 14'h2 : _GEN_382;
  wire [13:0] _GEN_384 = 14'h180 == index ? 14'h0 : _GEN_383;
  wire [13:0] _GEN_385 = 14'h181 == index ? 14'h180 : _GEN_384;
  wire [13:0] _GEN_386 = 14'h182 == index ? 14'h81 : _GEN_385;
  wire [13:0] _GEN_387 = 14'h183 == index ? 14'h80 : _GEN_386;
  wire [13:0] _GEN_388 = 14'h184 == index ? 14'h3 : _GEN_387;
  wire [13:0] _GEN_389 = 14'h185 == index ? 14'h3 : _GEN_388;
  wire [13:0] _GEN_390 = 14'h186 == index ? 14'h3 : _GEN_389;
  wire [13:0] _GEN_391 = 14'h187 == index ? 14'h3 : _GEN_390;
  wire [13:0] _GEN_392 = 14'h188 == index ? 14'h3 : _GEN_391;
  wire [13:0] _GEN_393 = 14'h189 == index ? 14'h3 : _GEN_392;
  wire [13:0] _GEN_394 = 14'h18a == index ? 14'h3 : _GEN_393;
  wire [13:0] _GEN_395 = 14'h18b == index ? 14'h3 : _GEN_394;
  wire [13:0] _GEN_396 = 14'h18c == index ? 14'h3 : _GEN_395;
  wire [13:0] _GEN_397 = 14'h18d == index ? 14'h3 : _GEN_396;
  wire [13:0] _GEN_398 = 14'h18e == index ? 14'h3 : _GEN_397;
  wire [13:0] _GEN_399 = 14'h18f == index ? 14'h3 : _GEN_398;
  wire [13:0] _GEN_400 = 14'h190 == index ? 14'h3 : _GEN_399;
  wire [13:0] _GEN_401 = 14'h191 == index ? 14'h3 : _GEN_400;
  wire [13:0] _GEN_402 = 14'h192 == index ? 14'h3 : _GEN_401;
  wire [13:0] _GEN_403 = 14'h193 == index ? 14'h3 : _GEN_402;
  wire [13:0] _GEN_404 = 14'h194 == index ? 14'h3 : _GEN_403;
  wire [13:0] _GEN_405 = 14'h195 == index ? 14'h3 : _GEN_404;
  wire [13:0] _GEN_406 = 14'h196 == index ? 14'h3 : _GEN_405;
  wire [13:0] _GEN_407 = 14'h197 == index ? 14'h3 : _GEN_406;
  wire [13:0] _GEN_408 = 14'h198 == index ? 14'h3 : _GEN_407;
  wire [13:0] _GEN_409 = 14'h199 == index ? 14'h3 : _GEN_408;
  wire [13:0] _GEN_410 = 14'h19a == index ? 14'h3 : _GEN_409;
  wire [13:0] _GEN_411 = 14'h19b == index ? 14'h3 : _GEN_410;
  wire [13:0] _GEN_412 = 14'h19c == index ? 14'h3 : _GEN_411;
  wire [13:0] _GEN_413 = 14'h19d == index ? 14'h3 : _GEN_412;
  wire [13:0] _GEN_414 = 14'h19e == index ? 14'h3 : _GEN_413;
  wire [13:0] _GEN_415 = 14'h19f == index ? 14'h3 : _GEN_414;
  wire [13:0] _GEN_416 = 14'h1a0 == index ? 14'h3 : _GEN_415;
  wire [13:0] _GEN_417 = 14'h1a1 == index ? 14'h3 : _GEN_416;
  wire [13:0] _GEN_418 = 14'h1a2 == index ? 14'h3 : _GEN_417;
  wire [13:0] _GEN_419 = 14'h1a3 == index ? 14'h3 : _GEN_418;
  wire [13:0] _GEN_420 = 14'h1a4 == index ? 14'h3 : _GEN_419;
  wire [13:0] _GEN_421 = 14'h1a5 == index ? 14'h3 : _GEN_420;
  wire [13:0] _GEN_422 = 14'h1a6 == index ? 14'h3 : _GEN_421;
  wire [13:0] _GEN_423 = 14'h1a7 == index ? 14'h3 : _GEN_422;
  wire [13:0] _GEN_424 = 14'h1a8 == index ? 14'h3 : _GEN_423;
  wire [13:0] _GEN_425 = 14'h1a9 == index ? 14'h3 : _GEN_424;
  wire [13:0] _GEN_426 = 14'h1aa == index ? 14'h3 : _GEN_425;
  wire [13:0] _GEN_427 = 14'h1ab == index ? 14'h3 : _GEN_426;
  wire [13:0] _GEN_428 = 14'h1ac == index ? 14'h3 : _GEN_427;
  wire [13:0] _GEN_429 = 14'h1ad == index ? 14'h3 : _GEN_428;
  wire [13:0] _GEN_430 = 14'h1ae == index ? 14'h3 : _GEN_429;
  wire [13:0] _GEN_431 = 14'h1af == index ? 14'h3 : _GEN_430;
  wire [13:0] _GEN_432 = 14'h1b0 == index ? 14'h3 : _GEN_431;
  wire [13:0] _GEN_433 = 14'h1b1 == index ? 14'h3 : _GEN_432;
  wire [13:0] _GEN_434 = 14'h1b2 == index ? 14'h3 : _GEN_433;
  wire [13:0] _GEN_435 = 14'h1b3 == index ? 14'h3 : _GEN_434;
  wire [13:0] _GEN_436 = 14'h1b4 == index ? 14'h3 : _GEN_435;
  wire [13:0] _GEN_437 = 14'h1b5 == index ? 14'h3 : _GEN_436;
  wire [13:0] _GEN_438 = 14'h1b6 == index ? 14'h3 : _GEN_437;
  wire [13:0] _GEN_439 = 14'h1b7 == index ? 14'h3 : _GEN_438;
  wire [13:0] _GEN_440 = 14'h1b8 == index ? 14'h3 : _GEN_439;
  wire [13:0] _GEN_441 = 14'h1b9 == index ? 14'h3 : _GEN_440;
  wire [13:0] _GEN_442 = 14'h1ba == index ? 14'h3 : _GEN_441;
  wire [13:0] _GEN_443 = 14'h1bb == index ? 14'h3 : _GEN_442;
  wire [13:0] _GEN_444 = 14'h1bc == index ? 14'h3 : _GEN_443;
  wire [13:0] _GEN_445 = 14'h1bd == index ? 14'h3 : _GEN_444;
  wire [13:0] _GEN_446 = 14'h1be == index ? 14'h3 : _GEN_445;
  wire [13:0] _GEN_447 = 14'h1bf == index ? 14'h3 : _GEN_446;
  wire [13:0] _GEN_448 = 14'h1c0 == index ? 14'h3 : _GEN_447;
  wire [13:0] _GEN_449 = 14'h1c1 == index ? 14'h3 : _GEN_448;
  wire [13:0] _GEN_450 = 14'h1c2 == index ? 14'h3 : _GEN_449;
  wire [13:0] _GEN_451 = 14'h1c3 == index ? 14'h3 : _GEN_450;
  wire [13:0] _GEN_452 = 14'h1c4 == index ? 14'h3 : _GEN_451;
  wire [13:0] _GEN_453 = 14'h1c5 == index ? 14'h3 : _GEN_452;
  wire [13:0] _GEN_454 = 14'h1c6 == index ? 14'h3 : _GEN_453;
  wire [13:0] _GEN_455 = 14'h1c7 == index ? 14'h3 : _GEN_454;
  wire [13:0] _GEN_456 = 14'h1c8 == index ? 14'h3 : _GEN_455;
  wire [13:0] _GEN_457 = 14'h1c9 == index ? 14'h3 : _GEN_456;
  wire [13:0] _GEN_458 = 14'h1ca == index ? 14'h3 : _GEN_457;
  wire [13:0] _GEN_459 = 14'h1cb == index ? 14'h3 : _GEN_458;
  wire [13:0] _GEN_460 = 14'h1cc == index ? 14'h3 : _GEN_459;
  wire [13:0] _GEN_461 = 14'h1cd == index ? 14'h3 : _GEN_460;
  wire [13:0] _GEN_462 = 14'h1ce == index ? 14'h3 : _GEN_461;
  wire [13:0] _GEN_463 = 14'h1cf == index ? 14'h3 : _GEN_462;
  wire [13:0] _GEN_464 = 14'h1d0 == index ? 14'h3 : _GEN_463;
  wire [13:0] _GEN_465 = 14'h1d1 == index ? 14'h3 : _GEN_464;
  wire [13:0] _GEN_466 = 14'h1d2 == index ? 14'h3 : _GEN_465;
  wire [13:0] _GEN_467 = 14'h1d3 == index ? 14'h3 : _GEN_466;
  wire [13:0] _GEN_468 = 14'h1d4 == index ? 14'h3 : _GEN_467;
  wire [13:0] _GEN_469 = 14'h1d5 == index ? 14'h3 : _GEN_468;
  wire [13:0] _GEN_470 = 14'h1d6 == index ? 14'h3 : _GEN_469;
  wire [13:0] _GEN_471 = 14'h1d7 == index ? 14'h3 : _GEN_470;
  wire [13:0] _GEN_472 = 14'h1d8 == index ? 14'h3 : _GEN_471;
  wire [13:0] _GEN_473 = 14'h1d9 == index ? 14'h3 : _GEN_472;
  wire [13:0] _GEN_474 = 14'h1da == index ? 14'h3 : _GEN_473;
  wire [13:0] _GEN_475 = 14'h1db == index ? 14'h3 : _GEN_474;
  wire [13:0] _GEN_476 = 14'h1dc == index ? 14'h3 : _GEN_475;
  wire [13:0] _GEN_477 = 14'h1dd == index ? 14'h3 : _GEN_476;
  wire [13:0] _GEN_478 = 14'h1de == index ? 14'h3 : _GEN_477;
  wire [13:0] _GEN_479 = 14'h1df == index ? 14'h3 : _GEN_478;
  wire [13:0] _GEN_480 = 14'h1e0 == index ? 14'h3 : _GEN_479;
  wire [13:0] _GEN_481 = 14'h1e1 == index ? 14'h3 : _GEN_480;
  wire [13:0] _GEN_482 = 14'h1e2 == index ? 14'h3 : _GEN_481;
  wire [13:0] _GEN_483 = 14'h1e3 == index ? 14'h3 : _GEN_482;
  wire [13:0] _GEN_484 = 14'h1e4 == index ? 14'h3 : _GEN_483;
  wire [13:0] _GEN_485 = 14'h1e5 == index ? 14'h3 : _GEN_484;
  wire [13:0] _GEN_486 = 14'h1e6 == index ? 14'h3 : _GEN_485;
  wire [13:0] _GEN_487 = 14'h1e7 == index ? 14'h3 : _GEN_486;
  wire [13:0] _GEN_488 = 14'h1e8 == index ? 14'h3 : _GEN_487;
  wire [13:0] _GEN_489 = 14'h1e9 == index ? 14'h3 : _GEN_488;
  wire [13:0] _GEN_490 = 14'h1ea == index ? 14'h3 : _GEN_489;
  wire [13:0] _GEN_491 = 14'h1eb == index ? 14'h3 : _GEN_490;
  wire [13:0] _GEN_492 = 14'h1ec == index ? 14'h3 : _GEN_491;
  wire [13:0] _GEN_493 = 14'h1ed == index ? 14'h3 : _GEN_492;
  wire [13:0] _GEN_494 = 14'h1ee == index ? 14'h3 : _GEN_493;
  wire [13:0] _GEN_495 = 14'h1ef == index ? 14'h3 : _GEN_494;
  wire [13:0] _GEN_496 = 14'h1f0 == index ? 14'h3 : _GEN_495;
  wire [13:0] _GEN_497 = 14'h1f1 == index ? 14'h3 : _GEN_496;
  wire [13:0] _GEN_498 = 14'h1f2 == index ? 14'h3 : _GEN_497;
  wire [13:0] _GEN_499 = 14'h1f3 == index ? 14'h3 : _GEN_498;
  wire [13:0] _GEN_500 = 14'h1f4 == index ? 14'h3 : _GEN_499;
  wire [13:0] _GEN_501 = 14'h1f5 == index ? 14'h3 : _GEN_500;
  wire [13:0] _GEN_502 = 14'h1f6 == index ? 14'h3 : _GEN_501;
  wire [13:0] _GEN_503 = 14'h1f7 == index ? 14'h3 : _GEN_502;
  wire [13:0] _GEN_504 = 14'h1f8 == index ? 14'h3 : _GEN_503;
  wire [13:0] _GEN_505 = 14'h1f9 == index ? 14'h3 : _GEN_504;
  wire [13:0] _GEN_506 = 14'h1fa == index ? 14'h3 : _GEN_505;
  wire [13:0] _GEN_507 = 14'h1fb == index ? 14'h3 : _GEN_506;
  wire [13:0] _GEN_508 = 14'h1fc == index ? 14'h3 : _GEN_507;
  wire [13:0] _GEN_509 = 14'h1fd == index ? 14'h3 : _GEN_508;
  wire [13:0] _GEN_510 = 14'h1fe == index ? 14'h3 : _GEN_509;
  wire [13:0] _GEN_511 = 14'h1ff == index ? 14'h3 : _GEN_510;
  wire [13:0] _GEN_512 = 14'h200 == index ? 14'h0 : _GEN_511;
  wire [13:0] _GEN_513 = 14'h201 == index ? 14'h200 : _GEN_512;
  wire [13:0] _GEN_514 = 14'h202 == index ? 14'h100 : _GEN_513;
  wire [13:0] _GEN_515 = 14'h203 == index ? 14'h81 : _GEN_514;
  wire [13:0] _GEN_516 = 14'h204 == index ? 14'h80 : _GEN_515;
  wire [13:0] _GEN_517 = 14'h205 == index ? 14'h4 : _GEN_516;
  wire [13:0] _GEN_518 = 14'h206 == index ? 14'h4 : _GEN_517;
  wire [13:0] _GEN_519 = 14'h207 == index ? 14'h4 : _GEN_518;
  wire [13:0] _GEN_520 = 14'h208 == index ? 14'h4 : _GEN_519;
  wire [13:0] _GEN_521 = 14'h209 == index ? 14'h4 : _GEN_520;
  wire [13:0] _GEN_522 = 14'h20a == index ? 14'h4 : _GEN_521;
  wire [13:0] _GEN_523 = 14'h20b == index ? 14'h4 : _GEN_522;
  wire [13:0] _GEN_524 = 14'h20c == index ? 14'h4 : _GEN_523;
  wire [13:0] _GEN_525 = 14'h20d == index ? 14'h4 : _GEN_524;
  wire [13:0] _GEN_526 = 14'h20e == index ? 14'h4 : _GEN_525;
  wire [13:0] _GEN_527 = 14'h20f == index ? 14'h4 : _GEN_526;
  wire [13:0] _GEN_528 = 14'h210 == index ? 14'h4 : _GEN_527;
  wire [13:0] _GEN_529 = 14'h211 == index ? 14'h4 : _GEN_528;
  wire [13:0] _GEN_530 = 14'h212 == index ? 14'h4 : _GEN_529;
  wire [13:0] _GEN_531 = 14'h213 == index ? 14'h4 : _GEN_530;
  wire [13:0] _GEN_532 = 14'h214 == index ? 14'h4 : _GEN_531;
  wire [13:0] _GEN_533 = 14'h215 == index ? 14'h4 : _GEN_532;
  wire [13:0] _GEN_534 = 14'h216 == index ? 14'h4 : _GEN_533;
  wire [13:0] _GEN_535 = 14'h217 == index ? 14'h4 : _GEN_534;
  wire [13:0] _GEN_536 = 14'h218 == index ? 14'h4 : _GEN_535;
  wire [13:0] _GEN_537 = 14'h219 == index ? 14'h4 : _GEN_536;
  wire [13:0] _GEN_538 = 14'h21a == index ? 14'h4 : _GEN_537;
  wire [13:0] _GEN_539 = 14'h21b == index ? 14'h4 : _GEN_538;
  wire [13:0] _GEN_540 = 14'h21c == index ? 14'h4 : _GEN_539;
  wire [13:0] _GEN_541 = 14'h21d == index ? 14'h4 : _GEN_540;
  wire [13:0] _GEN_542 = 14'h21e == index ? 14'h4 : _GEN_541;
  wire [13:0] _GEN_543 = 14'h21f == index ? 14'h4 : _GEN_542;
  wire [13:0] _GEN_544 = 14'h220 == index ? 14'h4 : _GEN_543;
  wire [13:0] _GEN_545 = 14'h221 == index ? 14'h4 : _GEN_544;
  wire [13:0] _GEN_546 = 14'h222 == index ? 14'h4 : _GEN_545;
  wire [13:0] _GEN_547 = 14'h223 == index ? 14'h4 : _GEN_546;
  wire [13:0] _GEN_548 = 14'h224 == index ? 14'h4 : _GEN_547;
  wire [13:0] _GEN_549 = 14'h225 == index ? 14'h4 : _GEN_548;
  wire [13:0] _GEN_550 = 14'h226 == index ? 14'h4 : _GEN_549;
  wire [13:0] _GEN_551 = 14'h227 == index ? 14'h4 : _GEN_550;
  wire [13:0] _GEN_552 = 14'h228 == index ? 14'h4 : _GEN_551;
  wire [13:0] _GEN_553 = 14'h229 == index ? 14'h4 : _GEN_552;
  wire [13:0] _GEN_554 = 14'h22a == index ? 14'h4 : _GEN_553;
  wire [13:0] _GEN_555 = 14'h22b == index ? 14'h4 : _GEN_554;
  wire [13:0] _GEN_556 = 14'h22c == index ? 14'h4 : _GEN_555;
  wire [13:0] _GEN_557 = 14'h22d == index ? 14'h4 : _GEN_556;
  wire [13:0] _GEN_558 = 14'h22e == index ? 14'h4 : _GEN_557;
  wire [13:0] _GEN_559 = 14'h22f == index ? 14'h4 : _GEN_558;
  wire [13:0] _GEN_560 = 14'h230 == index ? 14'h4 : _GEN_559;
  wire [13:0] _GEN_561 = 14'h231 == index ? 14'h4 : _GEN_560;
  wire [13:0] _GEN_562 = 14'h232 == index ? 14'h4 : _GEN_561;
  wire [13:0] _GEN_563 = 14'h233 == index ? 14'h4 : _GEN_562;
  wire [13:0] _GEN_564 = 14'h234 == index ? 14'h4 : _GEN_563;
  wire [13:0] _GEN_565 = 14'h235 == index ? 14'h4 : _GEN_564;
  wire [13:0] _GEN_566 = 14'h236 == index ? 14'h4 : _GEN_565;
  wire [13:0] _GEN_567 = 14'h237 == index ? 14'h4 : _GEN_566;
  wire [13:0] _GEN_568 = 14'h238 == index ? 14'h4 : _GEN_567;
  wire [13:0] _GEN_569 = 14'h239 == index ? 14'h4 : _GEN_568;
  wire [13:0] _GEN_570 = 14'h23a == index ? 14'h4 : _GEN_569;
  wire [13:0] _GEN_571 = 14'h23b == index ? 14'h4 : _GEN_570;
  wire [13:0] _GEN_572 = 14'h23c == index ? 14'h4 : _GEN_571;
  wire [13:0] _GEN_573 = 14'h23d == index ? 14'h4 : _GEN_572;
  wire [13:0] _GEN_574 = 14'h23e == index ? 14'h4 : _GEN_573;
  wire [13:0] _GEN_575 = 14'h23f == index ? 14'h4 : _GEN_574;
  wire [13:0] _GEN_576 = 14'h240 == index ? 14'h4 : _GEN_575;
  wire [13:0] _GEN_577 = 14'h241 == index ? 14'h4 : _GEN_576;
  wire [13:0] _GEN_578 = 14'h242 == index ? 14'h4 : _GEN_577;
  wire [13:0] _GEN_579 = 14'h243 == index ? 14'h4 : _GEN_578;
  wire [13:0] _GEN_580 = 14'h244 == index ? 14'h4 : _GEN_579;
  wire [13:0] _GEN_581 = 14'h245 == index ? 14'h4 : _GEN_580;
  wire [13:0] _GEN_582 = 14'h246 == index ? 14'h4 : _GEN_581;
  wire [13:0] _GEN_583 = 14'h247 == index ? 14'h4 : _GEN_582;
  wire [13:0] _GEN_584 = 14'h248 == index ? 14'h4 : _GEN_583;
  wire [13:0] _GEN_585 = 14'h249 == index ? 14'h4 : _GEN_584;
  wire [13:0] _GEN_586 = 14'h24a == index ? 14'h4 : _GEN_585;
  wire [13:0] _GEN_587 = 14'h24b == index ? 14'h4 : _GEN_586;
  wire [13:0] _GEN_588 = 14'h24c == index ? 14'h4 : _GEN_587;
  wire [13:0] _GEN_589 = 14'h24d == index ? 14'h4 : _GEN_588;
  wire [13:0] _GEN_590 = 14'h24e == index ? 14'h4 : _GEN_589;
  wire [13:0] _GEN_591 = 14'h24f == index ? 14'h4 : _GEN_590;
  wire [13:0] _GEN_592 = 14'h250 == index ? 14'h4 : _GEN_591;
  wire [13:0] _GEN_593 = 14'h251 == index ? 14'h4 : _GEN_592;
  wire [13:0] _GEN_594 = 14'h252 == index ? 14'h4 : _GEN_593;
  wire [13:0] _GEN_595 = 14'h253 == index ? 14'h4 : _GEN_594;
  wire [13:0] _GEN_596 = 14'h254 == index ? 14'h4 : _GEN_595;
  wire [13:0] _GEN_597 = 14'h255 == index ? 14'h4 : _GEN_596;
  wire [13:0] _GEN_598 = 14'h256 == index ? 14'h4 : _GEN_597;
  wire [13:0] _GEN_599 = 14'h257 == index ? 14'h4 : _GEN_598;
  wire [13:0] _GEN_600 = 14'h258 == index ? 14'h4 : _GEN_599;
  wire [13:0] _GEN_601 = 14'h259 == index ? 14'h4 : _GEN_600;
  wire [13:0] _GEN_602 = 14'h25a == index ? 14'h4 : _GEN_601;
  wire [13:0] _GEN_603 = 14'h25b == index ? 14'h4 : _GEN_602;
  wire [13:0] _GEN_604 = 14'h25c == index ? 14'h4 : _GEN_603;
  wire [13:0] _GEN_605 = 14'h25d == index ? 14'h4 : _GEN_604;
  wire [13:0] _GEN_606 = 14'h25e == index ? 14'h4 : _GEN_605;
  wire [13:0] _GEN_607 = 14'h25f == index ? 14'h4 : _GEN_606;
  wire [13:0] _GEN_608 = 14'h260 == index ? 14'h4 : _GEN_607;
  wire [13:0] _GEN_609 = 14'h261 == index ? 14'h4 : _GEN_608;
  wire [13:0] _GEN_610 = 14'h262 == index ? 14'h4 : _GEN_609;
  wire [13:0] _GEN_611 = 14'h263 == index ? 14'h4 : _GEN_610;
  wire [13:0] _GEN_612 = 14'h264 == index ? 14'h4 : _GEN_611;
  wire [13:0] _GEN_613 = 14'h265 == index ? 14'h4 : _GEN_612;
  wire [13:0] _GEN_614 = 14'h266 == index ? 14'h4 : _GEN_613;
  wire [13:0] _GEN_615 = 14'h267 == index ? 14'h4 : _GEN_614;
  wire [13:0] _GEN_616 = 14'h268 == index ? 14'h4 : _GEN_615;
  wire [13:0] _GEN_617 = 14'h269 == index ? 14'h4 : _GEN_616;
  wire [13:0] _GEN_618 = 14'h26a == index ? 14'h4 : _GEN_617;
  wire [13:0] _GEN_619 = 14'h26b == index ? 14'h4 : _GEN_618;
  wire [13:0] _GEN_620 = 14'h26c == index ? 14'h4 : _GEN_619;
  wire [13:0] _GEN_621 = 14'h26d == index ? 14'h4 : _GEN_620;
  wire [13:0] _GEN_622 = 14'h26e == index ? 14'h4 : _GEN_621;
  wire [13:0] _GEN_623 = 14'h26f == index ? 14'h4 : _GEN_622;
  wire [13:0] _GEN_624 = 14'h270 == index ? 14'h4 : _GEN_623;
  wire [13:0] _GEN_625 = 14'h271 == index ? 14'h4 : _GEN_624;
  wire [13:0] _GEN_626 = 14'h272 == index ? 14'h4 : _GEN_625;
  wire [13:0] _GEN_627 = 14'h273 == index ? 14'h4 : _GEN_626;
  wire [13:0] _GEN_628 = 14'h274 == index ? 14'h4 : _GEN_627;
  wire [13:0] _GEN_629 = 14'h275 == index ? 14'h4 : _GEN_628;
  wire [13:0] _GEN_630 = 14'h276 == index ? 14'h4 : _GEN_629;
  wire [13:0] _GEN_631 = 14'h277 == index ? 14'h4 : _GEN_630;
  wire [13:0] _GEN_632 = 14'h278 == index ? 14'h4 : _GEN_631;
  wire [13:0] _GEN_633 = 14'h279 == index ? 14'h4 : _GEN_632;
  wire [13:0] _GEN_634 = 14'h27a == index ? 14'h4 : _GEN_633;
  wire [13:0] _GEN_635 = 14'h27b == index ? 14'h4 : _GEN_634;
  wire [13:0] _GEN_636 = 14'h27c == index ? 14'h4 : _GEN_635;
  wire [13:0] _GEN_637 = 14'h27d == index ? 14'h4 : _GEN_636;
  wire [13:0] _GEN_638 = 14'h27e == index ? 14'h4 : _GEN_637;
  wire [13:0] _GEN_639 = 14'h27f == index ? 14'h4 : _GEN_638;
  wire [13:0] _GEN_640 = 14'h280 == index ? 14'h0 : _GEN_639;
  wire [13:0] _GEN_641 = 14'h281 == index ? 14'h280 : _GEN_640;
  wire [13:0] _GEN_642 = 14'h282 == index ? 14'h101 : _GEN_641;
  wire [13:0] _GEN_643 = 14'h283 == index ? 14'h82 : _GEN_642;
  wire [13:0] _GEN_644 = 14'h284 == index ? 14'h81 : _GEN_643;
  wire [13:0] _GEN_645 = 14'h285 == index ? 14'h80 : _GEN_644;
  wire [13:0] _GEN_646 = 14'h286 == index ? 14'h5 : _GEN_645;
  wire [13:0] _GEN_647 = 14'h287 == index ? 14'h5 : _GEN_646;
  wire [13:0] _GEN_648 = 14'h288 == index ? 14'h5 : _GEN_647;
  wire [13:0] _GEN_649 = 14'h289 == index ? 14'h5 : _GEN_648;
  wire [13:0] _GEN_650 = 14'h28a == index ? 14'h5 : _GEN_649;
  wire [13:0] _GEN_651 = 14'h28b == index ? 14'h5 : _GEN_650;
  wire [13:0] _GEN_652 = 14'h28c == index ? 14'h5 : _GEN_651;
  wire [13:0] _GEN_653 = 14'h28d == index ? 14'h5 : _GEN_652;
  wire [13:0] _GEN_654 = 14'h28e == index ? 14'h5 : _GEN_653;
  wire [13:0] _GEN_655 = 14'h28f == index ? 14'h5 : _GEN_654;
  wire [13:0] _GEN_656 = 14'h290 == index ? 14'h5 : _GEN_655;
  wire [13:0] _GEN_657 = 14'h291 == index ? 14'h5 : _GEN_656;
  wire [13:0] _GEN_658 = 14'h292 == index ? 14'h5 : _GEN_657;
  wire [13:0] _GEN_659 = 14'h293 == index ? 14'h5 : _GEN_658;
  wire [13:0] _GEN_660 = 14'h294 == index ? 14'h5 : _GEN_659;
  wire [13:0] _GEN_661 = 14'h295 == index ? 14'h5 : _GEN_660;
  wire [13:0] _GEN_662 = 14'h296 == index ? 14'h5 : _GEN_661;
  wire [13:0] _GEN_663 = 14'h297 == index ? 14'h5 : _GEN_662;
  wire [13:0] _GEN_664 = 14'h298 == index ? 14'h5 : _GEN_663;
  wire [13:0] _GEN_665 = 14'h299 == index ? 14'h5 : _GEN_664;
  wire [13:0] _GEN_666 = 14'h29a == index ? 14'h5 : _GEN_665;
  wire [13:0] _GEN_667 = 14'h29b == index ? 14'h5 : _GEN_666;
  wire [13:0] _GEN_668 = 14'h29c == index ? 14'h5 : _GEN_667;
  wire [13:0] _GEN_669 = 14'h29d == index ? 14'h5 : _GEN_668;
  wire [13:0] _GEN_670 = 14'h29e == index ? 14'h5 : _GEN_669;
  wire [13:0] _GEN_671 = 14'h29f == index ? 14'h5 : _GEN_670;
  wire [13:0] _GEN_672 = 14'h2a0 == index ? 14'h5 : _GEN_671;
  wire [13:0] _GEN_673 = 14'h2a1 == index ? 14'h5 : _GEN_672;
  wire [13:0] _GEN_674 = 14'h2a2 == index ? 14'h5 : _GEN_673;
  wire [13:0] _GEN_675 = 14'h2a3 == index ? 14'h5 : _GEN_674;
  wire [13:0] _GEN_676 = 14'h2a4 == index ? 14'h5 : _GEN_675;
  wire [13:0] _GEN_677 = 14'h2a5 == index ? 14'h5 : _GEN_676;
  wire [13:0] _GEN_678 = 14'h2a6 == index ? 14'h5 : _GEN_677;
  wire [13:0] _GEN_679 = 14'h2a7 == index ? 14'h5 : _GEN_678;
  wire [13:0] _GEN_680 = 14'h2a8 == index ? 14'h5 : _GEN_679;
  wire [13:0] _GEN_681 = 14'h2a9 == index ? 14'h5 : _GEN_680;
  wire [13:0] _GEN_682 = 14'h2aa == index ? 14'h5 : _GEN_681;
  wire [13:0] _GEN_683 = 14'h2ab == index ? 14'h5 : _GEN_682;
  wire [13:0] _GEN_684 = 14'h2ac == index ? 14'h5 : _GEN_683;
  wire [13:0] _GEN_685 = 14'h2ad == index ? 14'h5 : _GEN_684;
  wire [13:0] _GEN_686 = 14'h2ae == index ? 14'h5 : _GEN_685;
  wire [13:0] _GEN_687 = 14'h2af == index ? 14'h5 : _GEN_686;
  wire [13:0] _GEN_688 = 14'h2b0 == index ? 14'h5 : _GEN_687;
  wire [13:0] _GEN_689 = 14'h2b1 == index ? 14'h5 : _GEN_688;
  wire [13:0] _GEN_690 = 14'h2b2 == index ? 14'h5 : _GEN_689;
  wire [13:0] _GEN_691 = 14'h2b3 == index ? 14'h5 : _GEN_690;
  wire [13:0] _GEN_692 = 14'h2b4 == index ? 14'h5 : _GEN_691;
  wire [13:0] _GEN_693 = 14'h2b5 == index ? 14'h5 : _GEN_692;
  wire [13:0] _GEN_694 = 14'h2b6 == index ? 14'h5 : _GEN_693;
  wire [13:0] _GEN_695 = 14'h2b7 == index ? 14'h5 : _GEN_694;
  wire [13:0] _GEN_696 = 14'h2b8 == index ? 14'h5 : _GEN_695;
  wire [13:0] _GEN_697 = 14'h2b9 == index ? 14'h5 : _GEN_696;
  wire [13:0] _GEN_698 = 14'h2ba == index ? 14'h5 : _GEN_697;
  wire [13:0] _GEN_699 = 14'h2bb == index ? 14'h5 : _GEN_698;
  wire [13:0] _GEN_700 = 14'h2bc == index ? 14'h5 : _GEN_699;
  wire [13:0] _GEN_701 = 14'h2bd == index ? 14'h5 : _GEN_700;
  wire [13:0] _GEN_702 = 14'h2be == index ? 14'h5 : _GEN_701;
  wire [13:0] _GEN_703 = 14'h2bf == index ? 14'h5 : _GEN_702;
  wire [13:0] _GEN_704 = 14'h2c0 == index ? 14'h5 : _GEN_703;
  wire [13:0] _GEN_705 = 14'h2c1 == index ? 14'h5 : _GEN_704;
  wire [13:0] _GEN_706 = 14'h2c2 == index ? 14'h5 : _GEN_705;
  wire [13:0] _GEN_707 = 14'h2c3 == index ? 14'h5 : _GEN_706;
  wire [13:0] _GEN_708 = 14'h2c4 == index ? 14'h5 : _GEN_707;
  wire [13:0] _GEN_709 = 14'h2c5 == index ? 14'h5 : _GEN_708;
  wire [13:0] _GEN_710 = 14'h2c6 == index ? 14'h5 : _GEN_709;
  wire [13:0] _GEN_711 = 14'h2c7 == index ? 14'h5 : _GEN_710;
  wire [13:0] _GEN_712 = 14'h2c8 == index ? 14'h5 : _GEN_711;
  wire [13:0] _GEN_713 = 14'h2c9 == index ? 14'h5 : _GEN_712;
  wire [13:0] _GEN_714 = 14'h2ca == index ? 14'h5 : _GEN_713;
  wire [13:0] _GEN_715 = 14'h2cb == index ? 14'h5 : _GEN_714;
  wire [13:0] _GEN_716 = 14'h2cc == index ? 14'h5 : _GEN_715;
  wire [13:0] _GEN_717 = 14'h2cd == index ? 14'h5 : _GEN_716;
  wire [13:0] _GEN_718 = 14'h2ce == index ? 14'h5 : _GEN_717;
  wire [13:0] _GEN_719 = 14'h2cf == index ? 14'h5 : _GEN_718;
  wire [13:0] _GEN_720 = 14'h2d0 == index ? 14'h5 : _GEN_719;
  wire [13:0] _GEN_721 = 14'h2d1 == index ? 14'h5 : _GEN_720;
  wire [13:0] _GEN_722 = 14'h2d2 == index ? 14'h5 : _GEN_721;
  wire [13:0] _GEN_723 = 14'h2d3 == index ? 14'h5 : _GEN_722;
  wire [13:0] _GEN_724 = 14'h2d4 == index ? 14'h5 : _GEN_723;
  wire [13:0] _GEN_725 = 14'h2d5 == index ? 14'h5 : _GEN_724;
  wire [13:0] _GEN_726 = 14'h2d6 == index ? 14'h5 : _GEN_725;
  wire [13:0] _GEN_727 = 14'h2d7 == index ? 14'h5 : _GEN_726;
  wire [13:0] _GEN_728 = 14'h2d8 == index ? 14'h5 : _GEN_727;
  wire [13:0] _GEN_729 = 14'h2d9 == index ? 14'h5 : _GEN_728;
  wire [13:0] _GEN_730 = 14'h2da == index ? 14'h5 : _GEN_729;
  wire [13:0] _GEN_731 = 14'h2db == index ? 14'h5 : _GEN_730;
  wire [13:0] _GEN_732 = 14'h2dc == index ? 14'h5 : _GEN_731;
  wire [13:0] _GEN_733 = 14'h2dd == index ? 14'h5 : _GEN_732;
  wire [13:0] _GEN_734 = 14'h2de == index ? 14'h5 : _GEN_733;
  wire [13:0] _GEN_735 = 14'h2df == index ? 14'h5 : _GEN_734;
  wire [13:0] _GEN_736 = 14'h2e0 == index ? 14'h5 : _GEN_735;
  wire [13:0] _GEN_737 = 14'h2e1 == index ? 14'h5 : _GEN_736;
  wire [13:0] _GEN_738 = 14'h2e2 == index ? 14'h5 : _GEN_737;
  wire [13:0] _GEN_739 = 14'h2e3 == index ? 14'h5 : _GEN_738;
  wire [13:0] _GEN_740 = 14'h2e4 == index ? 14'h5 : _GEN_739;
  wire [13:0] _GEN_741 = 14'h2e5 == index ? 14'h5 : _GEN_740;
  wire [13:0] _GEN_742 = 14'h2e6 == index ? 14'h5 : _GEN_741;
  wire [13:0] _GEN_743 = 14'h2e7 == index ? 14'h5 : _GEN_742;
  wire [13:0] _GEN_744 = 14'h2e8 == index ? 14'h5 : _GEN_743;
  wire [13:0] _GEN_745 = 14'h2e9 == index ? 14'h5 : _GEN_744;
  wire [13:0] _GEN_746 = 14'h2ea == index ? 14'h5 : _GEN_745;
  wire [13:0] _GEN_747 = 14'h2eb == index ? 14'h5 : _GEN_746;
  wire [13:0] _GEN_748 = 14'h2ec == index ? 14'h5 : _GEN_747;
  wire [13:0] _GEN_749 = 14'h2ed == index ? 14'h5 : _GEN_748;
  wire [13:0] _GEN_750 = 14'h2ee == index ? 14'h5 : _GEN_749;
  wire [13:0] _GEN_751 = 14'h2ef == index ? 14'h5 : _GEN_750;
  wire [13:0] _GEN_752 = 14'h2f0 == index ? 14'h5 : _GEN_751;
  wire [13:0] _GEN_753 = 14'h2f1 == index ? 14'h5 : _GEN_752;
  wire [13:0] _GEN_754 = 14'h2f2 == index ? 14'h5 : _GEN_753;
  wire [13:0] _GEN_755 = 14'h2f3 == index ? 14'h5 : _GEN_754;
  wire [13:0] _GEN_756 = 14'h2f4 == index ? 14'h5 : _GEN_755;
  wire [13:0] _GEN_757 = 14'h2f5 == index ? 14'h5 : _GEN_756;
  wire [13:0] _GEN_758 = 14'h2f6 == index ? 14'h5 : _GEN_757;
  wire [13:0] _GEN_759 = 14'h2f7 == index ? 14'h5 : _GEN_758;
  wire [13:0] _GEN_760 = 14'h2f8 == index ? 14'h5 : _GEN_759;
  wire [13:0] _GEN_761 = 14'h2f9 == index ? 14'h5 : _GEN_760;
  wire [13:0] _GEN_762 = 14'h2fa == index ? 14'h5 : _GEN_761;
  wire [13:0] _GEN_763 = 14'h2fb == index ? 14'h5 : _GEN_762;
  wire [13:0] _GEN_764 = 14'h2fc == index ? 14'h5 : _GEN_763;
  wire [13:0] _GEN_765 = 14'h2fd == index ? 14'h5 : _GEN_764;
  wire [13:0] _GEN_766 = 14'h2fe == index ? 14'h5 : _GEN_765;
  wire [13:0] _GEN_767 = 14'h2ff == index ? 14'h5 : _GEN_766;
  wire [13:0] _GEN_768 = 14'h300 == index ? 14'h0 : _GEN_767;
  wire [13:0] _GEN_769 = 14'h301 == index ? 14'h300 : _GEN_768;
  wire [13:0] _GEN_770 = 14'h302 == index ? 14'h180 : _GEN_769;
  wire [13:0] _GEN_771 = 14'h303 == index ? 14'h100 : _GEN_770;
  wire [13:0] _GEN_772 = 14'h304 == index ? 14'h82 : _GEN_771;
  wire [13:0] _GEN_773 = 14'h305 == index ? 14'h81 : _GEN_772;
  wire [13:0] _GEN_774 = 14'h306 == index ? 14'h80 : _GEN_773;
  wire [13:0] _GEN_775 = 14'h307 == index ? 14'h6 : _GEN_774;
  wire [13:0] _GEN_776 = 14'h308 == index ? 14'h6 : _GEN_775;
  wire [13:0] _GEN_777 = 14'h309 == index ? 14'h6 : _GEN_776;
  wire [13:0] _GEN_778 = 14'h30a == index ? 14'h6 : _GEN_777;
  wire [13:0] _GEN_779 = 14'h30b == index ? 14'h6 : _GEN_778;
  wire [13:0] _GEN_780 = 14'h30c == index ? 14'h6 : _GEN_779;
  wire [13:0] _GEN_781 = 14'h30d == index ? 14'h6 : _GEN_780;
  wire [13:0] _GEN_782 = 14'h30e == index ? 14'h6 : _GEN_781;
  wire [13:0] _GEN_783 = 14'h30f == index ? 14'h6 : _GEN_782;
  wire [13:0] _GEN_784 = 14'h310 == index ? 14'h6 : _GEN_783;
  wire [13:0] _GEN_785 = 14'h311 == index ? 14'h6 : _GEN_784;
  wire [13:0] _GEN_786 = 14'h312 == index ? 14'h6 : _GEN_785;
  wire [13:0] _GEN_787 = 14'h313 == index ? 14'h6 : _GEN_786;
  wire [13:0] _GEN_788 = 14'h314 == index ? 14'h6 : _GEN_787;
  wire [13:0] _GEN_789 = 14'h315 == index ? 14'h6 : _GEN_788;
  wire [13:0] _GEN_790 = 14'h316 == index ? 14'h6 : _GEN_789;
  wire [13:0] _GEN_791 = 14'h317 == index ? 14'h6 : _GEN_790;
  wire [13:0] _GEN_792 = 14'h318 == index ? 14'h6 : _GEN_791;
  wire [13:0] _GEN_793 = 14'h319 == index ? 14'h6 : _GEN_792;
  wire [13:0] _GEN_794 = 14'h31a == index ? 14'h6 : _GEN_793;
  wire [13:0] _GEN_795 = 14'h31b == index ? 14'h6 : _GEN_794;
  wire [13:0] _GEN_796 = 14'h31c == index ? 14'h6 : _GEN_795;
  wire [13:0] _GEN_797 = 14'h31d == index ? 14'h6 : _GEN_796;
  wire [13:0] _GEN_798 = 14'h31e == index ? 14'h6 : _GEN_797;
  wire [13:0] _GEN_799 = 14'h31f == index ? 14'h6 : _GEN_798;
  wire [13:0] _GEN_800 = 14'h320 == index ? 14'h6 : _GEN_799;
  wire [13:0] _GEN_801 = 14'h321 == index ? 14'h6 : _GEN_800;
  wire [13:0] _GEN_802 = 14'h322 == index ? 14'h6 : _GEN_801;
  wire [13:0] _GEN_803 = 14'h323 == index ? 14'h6 : _GEN_802;
  wire [13:0] _GEN_804 = 14'h324 == index ? 14'h6 : _GEN_803;
  wire [13:0] _GEN_805 = 14'h325 == index ? 14'h6 : _GEN_804;
  wire [13:0] _GEN_806 = 14'h326 == index ? 14'h6 : _GEN_805;
  wire [13:0] _GEN_807 = 14'h327 == index ? 14'h6 : _GEN_806;
  wire [13:0] _GEN_808 = 14'h328 == index ? 14'h6 : _GEN_807;
  wire [13:0] _GEN_809 = 14'h329 == index ? 14'h6 : _GEN_808;
  wire [13:0] _GEN_810 = 14'h32a == index ? 14'h6 : _GEN_809;
  wire [13:0] _GEN_811 = 14'h32b == index ? 14'h6 : _GEN_810;
  wire [13:0] _GEN_812 = 14'h32c == index ? 14'h6 : _GEN_811;
  wire [13:0] _GEN_813 = 14'h32d == index ? 14'h6 : _GEN_812;
  wire [13:0] _GEN_814 = 14'h32e == index ? 14'h6 : _GEN_813;
  wire [13:0] _GEN_815 = 14'h32f == index ? 14'h6 : _GEN_814;
  wire [13:0] _GEN_816 = 14'h330 == index ? 14'h6 : _GEN_815;
  wire [13:0] _GEN_817 = 14'h331 == index ? 14'h6 : _GEN_816;
  wire [13:0] _GEN_818 = 14'h332 == index ? 14'h6 : _GEN_817;
  wire [13:0] _GEN_819 = 14'h333 == index ? 14'h6 : _GEN_818;
  wire [13:0] _GEN_820 = 14'h334 == index ? 14'h6 : _GEN_819;
  wire [13:0] _GEN_821 = 14'h335 == index ? 14'h6 : _GEN_820;
  wire [13:0] _GEN_822 = 14'h336 == index ? 14'h6 : _GEN_821;
  wire [13:0] _GEN_823 = 14'h337 == index ? 14'h6 : _GEN_822;
  wire [13:0] _GEN_824 = 14'h338 == index ? 14'h6 : _GEN_823;
  wire [13:0] _GEN_825 = 14'h339 == index ? 14'h6 : _GEN_824;
  wire [13:0] _GEN_826 = 14'h33a == index ? 14'h6 : _GEN_825;
  wire [13:0] _GEN_827 = 14'h33b == index ? 14'h6 : _GEN_826;
  wire [13:0] _GEN_828 = 14'h33c == index ? 14'h6 : _GEN_827;
  wire [13:0] _GEN_829 = 14'h33d == index ? 14'h6 : _GEN_828;
  wire [13:0] _GEN_830 = 14'h33e == index ? 14'h6 : _GEN_829;
  wire [13:0] _GEN_831 = 14'h33f == index ? 14'h6 : _GEN_830;
  wire [13:0] _GEN_832 = 14'h340 == index ? 14'h6 : _GEN_831;
  wire [13:0] _GEN_833 = 14'h341 == index ? 14'h6 : _GEN_832;
  wire [13:0] _GEN_834 = 14'h342 == index ? 14'h6 : _GEN_833;
  wire [13:0] _GEN_835 = 14'h343 == index ? 14'h6 : _GEN_834;
  wire [13:0] _GEN_836 = 14'h344 == index ? 14'h6 : _GEN_835;
  wire [13:0] _GEN_837 = 14'h345 == index ? 14'h6 : _GEN_836;
  wire [13:0] _GEN_838 = 14'h346 == index ? 14'h6 : _GEN_837;
  wire [13:0] _GEN_839 = 14'h347 == index ? 14'h6 : _GEN_838;
  wire [13:0] _GEN_840 = 14'h348 == index ? 14'h6 : _GEN_839;
  wire [13:0] _GEN_841 = 14'h349 == index ? 14'h6 : _GEN_840;
  wire [13:0] _GEN_842 = 14'h34a == index ? 14'h6 : _GEN_841;
  wire [13:0] _GEN_843 = 14'h34b == index ? 14'h6 : _GEN_842;
  wire [13:0] _GEN_844 = 14'h34c == index ? 14'h6 : _GEN_843;
  wire [13:0] _GEN_845 = 14'h34d == index ? 14'h6 : _GEN_844;
  wire [13:0] _GEN_846 = 14'h34e == index ? 14'h6 : _GEN_845;
  wire [13:0] _GEN_847 = 14'h34f == index ? 14'h6 : _GEN_846;
  wire [13:0] _GEN_848 = 14'h350 == index ? 14'h6 : _GEN_847;
  wire [13:0] _GEN_849 = 14'h351 == index ? 14'h6 : _GEN_848;
  wire [13:0] _GEN_850 = 14'h352 == index ? 14'h6 : _GEN_849;
  wire [13:0] _GEN_851 = 14'h353 == index ? 14'h6 : _GEN_850;
  wire [13:0] _GEN_852 = 14'h354 == index ? 14'h6 : _GEN_851;
  wire [13:0] _GEN_853 = 14'h355 == index ? 14'h6 : _GEN_852;
  wire [13:0] _GEN_854 = 14'h356 == index ? 14'h6 : _GEN_853;
  wire [13:0] _GEN_855 = 14'h357 == index ? 14'h6 : _GEN_854;
  wire [13:0] _GEN_856 = 14'h358 == index ? 14'h6 : _GEN_855;
  wire [13:0] _GEN_857 = 14'h359 == index ? 14'h6 : _GEN_856;
  wire [13:0] _GEN_858 = 14'h35a == index ? 14'h6 : _GEN_857;
  wire [13:0] _GEN_859 = 14'h35b == index ? 14'h6 : _GEN_858;
  wire [13:0] _GEN_860 = 14'h35c == index ? 14'h6 : _GEN_859;
  wire [13:0] _GEN_861 = 14'h35d == index ? 14'h6 : _GEN_860;
  wire [13:0] _GEN_862 = 14'h35e == index ? 14'h6 : _GEN_861;
  wire [13:0] _GEN_863 = 14'h35f == index ? 14'h6 : _GEN_862;
  wire [13:0] _GEN_864 = 14'h360 == index ? 14'h6 : _GEN_863;
  wire [13:0] _GEN_865 = 14'h361 == index ? 14'h6 : _GEN_864;
  wire [13:0] _GEN_866 = 14'h362 == index ? 14'h6 : _GEN_865;
  wire [13:0] _GEN_867 = 14'h363 == index ? 14'h6 : _GEN_866;
  wire [13:0] _GEN_868 = 14'h364 == index ? 14'h6 : _GEN_867;
  wire [13:0] _GEN_869 = 14'h365 == index ? 14'h6 : _GEN_868;
  wire [13:0] _GEN_870 = 14'h366 == index ? 14'h6 : _GEN_869;
  wire [13:0] _GEN_871 = 14'h367 == index ? 14'h6 : _GEN_870;
  wire [13:0] _GEN_872 = 14'h368 == index ? 14'h6 : _GEN_871;
  wire [13:0] _GEN_873 = 14'h369 == index ? 14'h6 : _GEN_872;
  wire [13:0] _GEN_874 = 14'h36a == index ? 14'h6 : _GEN_873;
  wire [13:0] _GEN_875 = 14'h36b == index ? 14'h6 : _GEN_874;
  wire [13:0] _GEN_876 = 14'h36c == index ? 14'h6 : _GEN_875;
  wire [13:0] _GEN_877 = 14'h36d == index ? 14'h6 : _GEN_876;
  wire [13:0] _GEN_878 = 14'h36e == index ? 14'h6 : _GEN_877;
  wire [13:0] _GEN_879 = 14'h36f == index ? 14'h6 : _GEN_878;
  wire [13:0] _GEN_880 = 14'h370 == index ? 14'h6 : _GEN_879;
  wire [13:0] _GEN_881 = 14'h371 == index ? 14'h6 : _GEN_880;
  wire [13:0] _GEN_882 = 14'h372 == index ? 14'h6 : _GEN_881;
  wire [13:0] _GEN_883 = 14'h373 == index ? 14'h6 : _GEN_882;
  wire [13:0] _GEN_884 = 14'h374 == index ? 14'h6 : _GEN_883;
  wire [13:0] _GEN_885 = 14'h375 == index ? 14'h6 : _GEN_884;
  wire [13:0] _GEN_886 = 14'h376 == index ? 14'h6 : _GEN_885;
  wire [13:0] _GEN_887 = 14'h377 == index ? 14'h6 : _GEN_886;
  wire [13:0] _GEN_888 = 14'h378 == index ? 14'h6 : _GEN_887;
  wire [13:0] _GEN_889 = 14'h379 == index ? 14'h6 : _GEN_888;
  wire [13:0] _GEN_890 = 14'h37a == index ? 14'h6 : _GEN_889;
  wire [13:0] _GEN_891 = 14'h37b == index ? 14'h6 : _GEN_890;
  wire [13:0] _GEN_892 = 14'h37c == index ? 14'h6 : _GEN_891;
  wire [13:0] _GEN_893 = 14'h37d == index ? 14'h6 : _GEN_892;
  wire [13:0] _GEN_894 = 14'h37e == index ? 14'h6 : _GEN_893;
  wire [13:0] _GEN_895 = 14'h37f == index ? 14'h6 : _GEN_894;
  wire [13:0] _GEN_896 = 14'h380 == index ? 14'h0 : _GEN_895;
  wire [13:0] _GEN_897 = 14'h381 == index ? 14'h380 : _GEN_896;
  wire [13:0] _GEN_898 = 14'h382 == index ? 14'h181 : _GEN_897;
  wire [13:0] _GEN_899 = 14'h383 == index ? 14'h101 : _GEN_898;
  wire [13:0] _GEN_900 = 14'h384 == index ? 14'h83 : _GEN_899;
  wire [13:0] _GEN_901 = 14'h385 == index ? 14'h82 : _GEN_900;
  wire [13:0] _GEN_902 = 14'h386 == index ? 14'h81 : _GEN_901;
  wire [13:0] _GEN_903 = 14'h387 == index ? 14'h80 : _GEN_902;
  wire [13:0] _GEN_904 = 14'h388 == index ? 14'h7 : _GEN_903;
  wire [13:0] _GEN_905 = 14'h389 == index ? 14'h7 : _GEN_904;
  wire [13:0] _GEN_906 = 14'h38a == index ? 14'h7 : _GEN_905;
  wire [13:0] _GEN_907 = 14'h38b == index ? 14'h7 : _GEN_906;
  wire [13:0] _GEN_908 = 14'h38c == index ? 14'h7 : _GEN_907;
  wire [13:0] _GEN_909 = 14'h38d == index ? 14'h7 : _GEN_908;
  wire [13:0] _GEN_910 = 14'h38e == index ? 14'h7 : _GEN_909;
  wire [13:0] _GEN_911 = 14'h38f == index ? 14'h7 : _GEN_910;
  wire [13:0] _GEN_912 = 14'h390 == index ? 14'h7 : _GEN_911;
  wire [13:0] _GEN_913 = 14'h391 == index ? 14'h7 : _GEN_912;
  wire [13:0] _GEN_914 = 14'h392 == index ? 14'h7 : _GEN_913;
  wire [13:0] _GEN_915 = 14'h393 == index ? 14'h7 : _GEN_914;
  wire [13:0] _GEN_916 = 14'h394 == index ? 14'h7 : _GEN_915;
  wire [13:0] _GEN_917 = 14'h395 == index ? 14'h7 : _GEN_916;
  wire [13:0] _GEN_918 = 14'h396 == index ? 14'h7 : _GEN_917;
  wire [13:0] _GEN_919 = 14'h397 == index ? 14'h7 : _GEN_918;
  wire [13:0] _GEN_920 = 14'h398 == index ? 14'h7 : _GEN_919;
  wire [13:0] _GEN_921 = 14'h399 == index ? 14'h7 : _GEN_920;
  wire [13:0] _GEN_922 = 14'h39a == index ? 14'h7 : _GEN_921;
  wire [13:0] _GEN_923 = 14'h39b == index ? 14'h7 : _GEN_922;
  wire [13:0] _GEN_924 = 14'h39c == index ? 14'h7 : _GEN_923;
  wire [13:0] _GEN_925 = 14'h39d == index ? 14'h7 : _GEN_924;
  wire [13:0] _GEN_926 = 14'h39e == index ? 14'h7 : _GEN_925;
  wire [13:0] _GEN_927 = 14'h39f == index ? 14'h7 : _GEN_926;
  wire [13:0] _GEN_928 = 14'h3a0 == index ? 14'h7 : _GEN_927;
  wire [13:0] _GEN_929 = 14'h3a1 == index ? 14'h7 : _GEN_928;
  wire [13:0] _GEN_930 = 14'h3a2 == index ? 14'h7 : _GEN_929;
  wire [13:0] _GEN_931 = 14'h3a3 == index ? 14'h7 : _GEN_930;
  wire [13:0] _GEN_932 = 14'h3a4 == index ? 14'h7 : _GEN_931;
  wire [13:0] _GEN_933 = 14'h3a5 == index ? 14'h7 : _GEN_932;
  wire [13:0] _GEN_934 = 14'h3a6 == index ? 14'h7 : _GEN_933;
  wire [13:0] _GEN_935 = 14'h3a7 == index ? 14'h7 : _GEN_934;
  wire [13:0] _GEN_936 = 14'h3a8 == index ? 14'h7 : _GEN_935;
  wire [13:0] _GEN_937 = 14'h3a9 == index ? 14'h7 : _GEN_936;
  wire [13:0] _GEN_938 = 14'h3aa == index ? 14'h7 : _GEN_937;
  wire [13:0] _GEN_939 = 14'h3ab == index ? 14'h7 : _GEN_938;
  wire [13:0] _GEN_940 = 14'h3ac == index ? 14'h7 : _GEN_939;
  wire [13:0] _GEN_941 = 14'h3ad == index ? 14'h7 : _GEN_940;
  wire [13:0] _GEN_942 = 14'h3ae == index ? 14'h7 : _GEN_941;
  wire [13:0] _GEN_943 = 14'h3af == index ? 14'h7 : _GEN_942;
  wire [13:0] _GEN_944 = 14'h3b0 == index ? 14'h7 : _GEN_943;
  wire [13:0] _GEN_945 = 14'h3b1 == index ? 14'h7 : _GEN_944;
  wire [13:0] _GEN_946 = 14'h3b2 == index ? 14'h7 : _GEN_945;
  wire [13:0] _GEN_947 = 14'h3b3 == index ? 14'h7 : _GEN_946;
  wire [13:0] _GEN_948 = 14'h3b4 == index ? 14'h7 : _GEN_947;
  wire [13:0] _GEN_949 = 14'h3b5 == index ? 14'h7 : _GEN_948;
  wire [13:0] _GEN_950 = 14'h3b6 == index ? 14'h7 : _GEN_949;
  wire [13:0] _GEN_951 = 14'h3b7 == index ? 14'h7 : _GEN_950;
  wire [13:0] _GEN_952 = 14'h3b8 == index ? 14'h7 : _GEN_951;
  wire [13:0] _GEN_953 = 14'h3b9 == index ? 14'h7 : _GEN_952;
  wire [13:0] _GEN_954 = 14'h3ba == index ? 14'h7 : _GEN_953;
  wire [13:0] _GEN_955 = 14'h3bb == index ? 14'h7 : _GEN_954;
  wire [13:0] _GEN_956 = 14'h3bc == index ? 14'h7 : _GEN_955;
  wire [13:0] _GEN_957 = 14'h3bd == index ? 14'h7 : _GEN_956;
  wire [13:0] _GEN_958 = 14'h3be == index ? 14'h7 : _GEN_957;
  wire [13:0] _GEN_959 = 14'h3bf == index ? 14'h7 : _GEN_958;
  wire [13:0] _GEN_960 = 14'h3c0 == index ? 14'h7 : _GEN_959;
  wire [13:0] _GEN_961 = 14'h3c1 == index ? 14'h7 : _GEN_960;
  wire [13:0] _GEN_962 = 14'h3c2 == index ? 14'h7 : _GEN_961;
  wire [13:0] _GEN_963 = 14'h3c3 == index ? 14'h7 : _GEN_962;
  wire [13:0] _GEN_964 = 14'h3c4 == index ? 14'h7 : _GEN_963;
  wire [13:0] _GEN_965 = 14'h3c5 == index ? 14'h7 : _GEN_964;
  wire [13:0] _GEN_966 = 14'h3c6 == index ? 14'h7 : _GEN_965;
  wire [13:0] _GEN_967 = 14'h3c7 == index ? 14'h7 : _GEN_966;
  wire [13:0] _GEN_968 = 14'h3c8 == index ? 14'h7 : _GEN_967;
  wire [13:0] _GEN_969 = 14'h3c9 == index ? 14'h7 : _GEN_968;
  wire [13:0] _GEN_970 = 14'h3ca == index ? 14'h7 : _GEN_969;
  wire [13:0] _GEN_971 = 14'h3cb == index ? 14'h7 : _GEN_970;
  wire [13:0] _GEN_972 = 14'h3cc == index ? 14'h7 : _GEN_971;
  wire [13:0] _GEN_973 = 14'h3cd == index ? 14'h7 : _GEN_972;
  wire [13:0] _GEN_974 = 14'h3ce == index ? 14'h7 : _GEN_973;
  wire [13:0] _GEN_975 = 14'h3cf == index ? 14'h7 : _GEN_974;
  wire [13:0] _GEN_976 = 14'h3d0 == index ? 14'h7 : _GEN_975;
  wire [13:0] _GEN_977 = 14'h3d1 == index ? 14'h7 : _GEN_976;
  wire [13:0] _GEN_978 = 14'h3d2 == index ? 14'h7 : _GEN_977;
  wire [13:0] _GEN_979 = 14'h3d3 == index ? 14'h7 : _GEN_978;
  wire [13:0] _GEN_980 = 14'h3d4 == index ? 14'h7 : _GEN_979;
  wire [13:0] _GEN_981 = 14'h3d5 == index ? 14'h7 : _GEN_980;
  wire [13:0] _GEN_982 = 14'h3d6 == index ? 14'h7 : _GEN_981;
  wire [13:0] _GEN_983 = 14'h3d7 == index ? 14'h7 : _GEN_982;
  wire [13:0] _GEN_984 = 14'h3d8 == index ? 14'h7 : _GEN_983;
  wire [13:0] _GEN_985 = 14'h3d9 == index ? 14'h7 : _GEN_984;
  wire [13:0] _GEN_986 = 14'h3da == index ? 14'h7 : _GEN_985;
  wire [13:0] _GEN_987 = 14'h3db == index ? 14'h7 : _GEN_986;
  wire [13:0] _GEN_988 = 14'h3dc == index ? 14'h7 : _GEN_987;
  wire [13:0] _GEN_989 = 14'h3dd == index ? 14'h7 : _GEN_988;
  wire [13:0] _GEN_990 = 14'h3de == index ? 14'h7 : _GEN_989;
  wire [13:0] _GEN_991 = 14'h3df == index ? 14'h7 : _GEN_990;
  wire [13:0] _GEN_992 = 14'h3e0 == index ? 14'h7 : _GEN_991;
  wire [13:0] _GEN_993 = 14'h3e1 == index ? 14'h7 : _GEN_992;
  wire [13:0] _GEN_994 = 14'h3e2 == index ? 14'h7 : _GEN_993;
  wire [13:0] _GEN_995 = 14'h3e3 == index ? 14'h7 : _GEN_994;
  wire [13:0] _GEN_996 = 14'h3e4 == index ? 14'h7 : _GEN_995;
  wire [13:0] _GEN_997 = 14'h3e5 == index ? 14'h7 : _GEN_996;
  wire [13:0] _GEN_998 = 14'h3e6 == index ? 14'h7 : _GEN_997;
  wire [13:0] _GEN_999 = 14'h3e7 == index ? 14'h7 : _GEN_998;
  wire [13:0] _GEN_1000 = 14'h3e8 == index ? 14'h7 : _GEN_999;
  wire [13:0] _GEN_1001 = 14'h3e9 == index ? 14'h7 : _GEN_1000;
  wire [13:0] _GEN_1002 = 14'h3ea == index ? 14'h7 : _GEN_1001;
  wire [13:0] _GEN_1003 = 14'h3eb == index ? 14'h7 : _GEN_1002;
  wire [13:0] _GEN_1004 = 14'h3ec == index ? 14'h7 : _GEN_1003;
  wire [13:0] _GEN_1005 = 14'h3ed == index ? 14'h7 : _GEN_1004;
  wire [13:0] _GEN_1006 = 14'h3ee == index ? 14'h7 : _GEN_1005;
  wire [13:0] _GEN_1007 = 14'h3ef == index ? 14'h7 : _GEN_1006;
  wire [13:0] _GEN_1008 = 14'h3f0 == index ? 14'h7 : _GEN_1007;
  wire [13:0] _GEN_1009 = 14'h3f1 == index ? 14'h7 : _GEN_1008;
  wire [13:0] _GEN_1010 = 14'h3f2 == index ? 14'h7 : _GEN_1009;
  wire [13:0] _GEN_1011 = 14'h3f3 == index ? 14'h7 : _GEN_1010;
  wire [13:0] _GEN_1012 = 14'h3f4 == index ? 14'h7 : _GEN_1011;
  wire [13:0] _GEN_1013 = 14'h3f5 == index ? 14'h7 : _GEN_1012;
  wire [13:0] _GEN_1014 = 14'h3f6 == index ? 14'h7 : _GEN_1013;
  wire [13:0] _GEN_1015 = 14'h3f7 == index ? 14'h7 : _GEN_1014;
  wire [13:0] _GEN_1016 = 14'h3f8 == index ? 14'h7 : _GEN_1015;
  wire [13:0] _GEN_1017 = 14'h3f9 == index ? 14'h7 : _GEN_1016;
  wire [13:0] _GEN_1018 = 14'h3fa == index ? 14'h7 : _GEN_1017;
  wire [13:0] _GEN_1019 = 14'h3fb == index ? 14'h7 : _GEN_1018;
  wire [13:0] _GEN_1020 = 14'h3fc == index ? 14'h7 : _GEN_1019;
  wire [13:0] _GEN_1021 = 14'h3fd == index ? 14'h7 : _GEN_1020;
  wire [13:0] _GEN_1022 = 14'h3fe == index ? 14'h7 : _GEN_1021;
  wire [13:0] _GEN_1023 = 14'h3ff == index ? 14'h7 : _GEN_1022;
  wire [13:0] _GEN_1024 = 14'h400 == index ? 14'h0 : _GEN_1023;
  wire [13:0] _GEN_1025 = 14'h401 == index ? 14'h400 : _GEN_1024;
  wire [13:0] _GEN_1026 = 14'h402 == index ? 14'h200 : _GEN_1025;
  wire [13:0] _GEN_1027 = 14'h403 == index ? 14'h102 : _GEN_1026;
  wire [13:0] _GEN_1028 = 14'h404 == index ? 14'h100 : _GEN_1027;
  wire [13:0] _GEN_1029 = 14'h405 == index ? 14'h83 : _GEN_1028;
  wire [13:0] _GEN_1030 = 14'h406 == index ? 14'h82 : _GEN_1029;
  wire [13:0] _GEN_1031 = 14'h407 == index ? 14'h81 : _GEN_1030;
  wire [13:0] _GEN_1032 = 14'h408 == index ? 14'h80 : _GEN_1031;
  wire [13:0] _GEN_1033 = 14'h409 == index ? 14'h8 : _GEN_1032;
  wire [13:0] _GEN_1034 = 14'h40a == index ? 14'h8 : _GEN_1033;
  wire [13:0] _GEN_1035 = 14'h40b == index ? 14'h8 : _GEN_1034;
  wire [13:0] _GEN_1036 = 14'h40c == index ? 14'h8 : _GEN_1035;
  wire [13:0] _GEN_1037 = 14'h40d == index ? 14'h8 : _GEN_1036;
  wire [13:0] _GEN_1038 = 14'h40e == index ? 14'h8 : _GEN_1037;
  wire [13:0] _GEN_1039 = 14'h40f == index ? 14'h8 : _GEN_1038;
  wire [13:0] _GEN_1040 = 14'h410 == index ? 14'h8 : _GEN_1039;
  wire [13:0] _GEN_1041 = 14'h411 == index ? 14'h8 : _GEN_1040;
  wire [13:0] _GEN_1042 = 14'h412 == index ? 14'h8 : _GEN_1041;
  wire [13:0] _GEN_1043 = 14'h413 == index ? 14'h8 : _GEN_1042;
  wire [13:0] _GEN_1044 = 14'h414 == index ? 14'h8 : _GEN_1043;
  wire [13:0] _GEN_1045 = 14'h415 == index ? 14'h8 : _GEN_1044;
  wire [13:0] _GEN_1046 = 14'h416 == index ? 14'h8 : _GEN_1045;
  wire [13:0] _GEN_1047 = 14'h417 == index ? 14'h8 : _GEN_1046;
  wire [13:0] _GEN_1048 = 14'h418 == index ? 14'h8 : _GEN_1047;
  wire [13:0] _GEN_1049 = 14'h419 == index ? 14'h8 : _GEN_1048;
  wire [13:0] _GEN_1050 = 14'h41a == index ? 14'h8 : _GEN_1049;
  wire [13:0] _GEN_1051 = 14'h41b == index ? 14'h8 : _GEN_1050;
  wire [13:0] _GEN_1052 = 14'h41c == index ? 14'h8 : _GEN_1051;
  wire [13:0] _GEN_1053 = 14'h41d == index ? 14'h8 : _GEN_1052;
  wire [13:0] _GEN_1054 = 14'h41e == index ? 14'h8 : _GEN_1053;
  wire [13:0] _GEN_1055 = 14'h41f == index ? 14'h8 : _GEN_1054;
  wire [13:0] _GEN_1056 = 14'h420 == index ? 14'h8 : _GEN_1055;
  wire [13:0] _GEN_1057 = 14'h421 == index ? 14'h8 : _GEN_1056;
  wire [13:0] _GEN_1058 = 14'h422 == index ? 14'h8 : _GEN_1057;
  wire [13:0] _GEN_1059 = 14'h423 == index ? 14'h8 : _GEN_1058;
  wire [13:0] _GEN_1060 = 14'h424 == index ? 14'h8 : _GEN_1059;
  wire [13:0] _GEN_1061 = 14'h425 == index ? 14'h8 : _GEN_1060;
  wire [13:0] _GEN_1062 = 14'h426 == index ? 14'h8 : _GEN_1061;
  wire [13:0] _GEN_1063 = 14'h427 == index ? 14'h8 : _GEN_1062;
  wire [13:0] _GEN_1064 = 14'h428 == index ? 14'h8 : _GEN_1063;
  wire [13:0] _GEN_1065 = 14'h429 == index ? 14'h8 : _GEN_1064;
  wire [13:0] _GEN_1066 = 14'h42a == index ? 14'h8 : _GEN_1065;
  wire [13:0] _GEN_1067 = 14'h42b == index ? 14'h8 : _GEN_1066;
  wire [13:0] _GEN_1068 = 14'h42c == index ? 14'h8 : _GEN_1067;
  wire [13:0] _GEN_1069 = 14'h42d == index ? 14'h8 : _GEN_1068;
  wire [13:0] _GEN_1070 = 14'h42e == index ? 14'h8 : _GEN_1069;
  wire [13:0] _GEN_1071 = 14'h42f == index ? 14'h8 : _GEN_1070;
  wire [13:0] _GEN_1072 = 14'h430 == index ? 14'h8 : _GEN_1071;
  wire [13:0] _GEN_1073 = 14'h431 == index ? 14'h8 : _GEN_1072;
  wire [13:0] _GEN_1074 = 14'h432 == index ? 14'h8 : _GEN_1073;
  wire [13:0] _GEN_1075 = 14'h433 == index ? 14'h8 : _GEN_1074;
  wire [13:0] _GEN_1076 = 14'h434 == index ? 14'h8 : _GEN_1075;
  wire [13:0] _GEN_1077 = 14'h435 == index ? 14'h8 : _GEN_1076;
  wire [13:0] _GEN_1078 = 14'h436 == index ? 14'h8 : _GEN_1077;
  wire [13:0] _GEN_1079 = 14'h437 == index ? 14'h8 : _GEN_1078;
  wire [13:0] _GEN_1080 = 14'h438 == index ? 14'h8 : _GEN_1079;
  wire [13:0] _GEN_1081 = 14'h439 == index ? 14'h8 : _GEN_1080;
  wire [13:0] _GEN_1082 = 14'h43a == index ? 14'h8 : _GEN_1081;
  wire [13:0] _GEN_1083 = 14'h43b == index ? 14'h8 : _GEN_1082;
  wire [13:0] _GEN_1084 = 14'h43c == index ? 14'h8 : _GEN_1083;
  wire [13:0] _GEN_1085 = 14'h43d == index ? 14'h8 : _GEN_1084;
  wire [13:0] _GEN_1086 = 14'h43e == index ? 14'h8 : _GEN_1085;
  wire [13:0] _GEN_1087 = 14'h43f == index ? 14'h8 : _GEN_1086;
  wire [13:0] _GEN_1088 = 14'h440 == index ? 14'h8 : _GEN_1087;
  wire [13:0] _GEN_1089 = 14'h441 == index ? 14'h8 : _GEN_1088;
  wire [13:0] _GEN_1090 = 14'h442 == index ? 14'h8 : _GEN_1089;
  wire [13:0] _GEN_1091 = 14'h443 == index ? 14'h8 : _GEN_1090;
  wire [13:0] _GEN_1092 = 14'h444 == index ? 14'h8 : _GEN_1091;
  wire [13:0] _GEN_1093 = 14'h445 == index ? 14'h8 : _GEN_1092;
  wire [13:0] _GEN_1094 = 14'h446 == index ? 14'h8 : _GEN_1093;
  wire [13:0] _GEN_1095 = 14'h447 == index ? 14'h8 : _GEN_1094;
  wire [13:0] _GEN_1096 = 14'h448 == index ? 14'h8 : _GEN_1095;
  wire [13:0] _GEN_1097 = 14'h449 == index ? 14'h8 : _GEN_1096;
  wire [13:0] _GEN_1098 = 14'h44a == index ? 14'h8 : _GEN_1097;
  wire [13:0] _GEN_1099 = 14'h44b == index ? 14'h8 : _GEN_1098;
  wire [13:0] _GEN_1100 = 14'h44c == index ? 14'h8 : _GEN_1099;
  wire [13:0] _GEN_1101 = 14'h44d == index ? 14'h8 : _GEN_1100;
  wire [13:0] _GEN_1102 = 14'h44e == index ? 14'h8 : _GEN_1101;
  wire [13:0] _GEN_1103 = 14'h44f == index ? 14'h8 : _GEN_1102;
  wire [13:0] _GEN_1104 = 14'h450 == index ? 14'h8 : _GEN_1103;
  wire [13:0] _GEN_1105 = 14'h451 == index ? 14'h8 : _GEN_1104;
  wire [13:0] _GEN_1106 = 14'h452 == index ? 14'h8 : _GEN_1105;
  wire [13:0] _GEN_1107 = 14'h453 == index ? 14'h8 : _GEN_1106;
  wire [13:0] _GEN_1108 = 14'h454 == index ? 14'h8 : _GEN_1107;
  wire [13:0] _GEN_1109 = 14'h455 == index ? 14'h8 : _GEN_1108;
  wire [13:0] _GEN_1110 = 14'h456 == index ? 14'h8 : _GEN_1109;
  wire [13:0] _GEN_1111 = 14'h457 == index ? 14'h8 : _GEN_1110;
  wire [13:0] _GEN_1112 = 14'h458 == index ? 14'h8 : _GEN_1111;
  wire [13:0] _GEN_1113 = 14'h459 == index ? 14'h8 : _GEN_1112;
  wire [13:0] _GEN_1114 = 14'h45a == index ? 14'h8 : _GEN_1113;
  wire [13:0] _GEN_1115 = 14'h45b == index ? 14'h8 : _GEN_1114;
  wire [13:0] _GEN_1116 = 14'h45c == index ? 14'h8 : _GEN_1115;
  wire [13:0] _GEN_1117 = 14'h45d == index ? 14'h8 : _GEN_1116;
  wire [13:0] _GEN_1118 = 14'h45e == index ? 14'h8 : _GEN_1117;
  wire [13:0] _GEN_1119 = 14'h45f == index ? 14'h8 : _GEN_1118;
  wire [13:0] _GEN_1120 = 14'h460 == index ? 14'h8 : _GEN_1119;
  wire [13:0] _GEN_1121 = 14'h461 == index ? 14'h8 : _GEN_1120;
  wire [13:0] _GEN_1122 = 14'h462 == index ? 14'h8 : _GEN_1121;
  wire [13:0] _GEN_1123 = 14'h463 == index ? 14'h8 : _GEN_1122;
  wire [13:0] _GEN_1124 = 14'h464 == index ? 14'h8 : _GEN_1123;
  wire [13:0] _GEN_1125 = 14'h465 == index ? 14'h8 : _GEN_1124;
  wire [13:0] _GEN_1126 = 14'h466 == index ? 14'h8 : _GEN_1125;
  wire [13:0] _GEN_1127 = 14'h467 == index ? 14'h8 : _GEN_1126;
  wire [13:0] _GEN_1128 = 14'h468 == index ? 14'h8 : _GEN_1127;
  wire [13:0] _GEN_1129 = 14'h469 == index ? 14'h8 : _GEN_1128;
  wire [13:0] _GEN_1130 = 14'h46a == index ? 14'h8 : _GEN_1129;
  wire [13:0] _GEN_1131 = 14'h46b == index ? 14'h8 : _GEN_1130;
  wire [13:0] _GEN_1132 = 14'h46c == index ? 14'h8 : _GEN_1131;
  wire [13:0] _GEN_1133 = 14'h46d == index ? 14'h8 : _GEN_1132;
  wire [13:0] _GEN_1134 = 14'h46e == index ? 14'h8 : _GEN_1133;
  wire [13:0] _GEN_1135 = 14'h46f == index ? 14'h8 : _GEN_1134;
  wire [13:0] _GEN_1136 = 14'h470 == index ? 14'h8 : _GEN_1135;
  wire [13:0] _GEN_1137 = 14'h471 == index ? 14'h8 : _GEN_1136;
  wire [13:0] _GEN_1138 = 14'h472 == index ? 14'h8 : _GEN_1137;
  wire [13:0] _GEN_1139 = 14'h473 == index ? 14'h8 : _GEN_1138;
  wire [13:0] _GEN_1140 = 14'h474 == index ? 14'h8 : _GEN_1139;
  wire [13:0] _GEN_1141 = 14'h475 == index ? 14'h8 : _GEN_1140;
  wire [13:0] _GEN_1142 = 14'h476 == index ? 14'h8 : _GEN_1141;
  wire [13:0] _GEN_1143 = 14'h477 == index ? 14'h8 : _GEN_1142;
  wire [13:0] _GEN_1144 = 14'h478 == index ? 14'h8 : _GEN_1143;
  wire [13:0] _GEN_1145 = 14'h479 == index ? 14'h8 : _GEN_1144;
  wire [13:0] _GEN_1146 = 14'h47a == index ? 14'h8 : _GEN_1145;
  wire [13:0] _GEN_1147 = 14'h47b == index ? 14'h8 : _GEN_1146;
  wire [13:0] _GEN_1148 = 14'h47c == index ? 14'h8 : _GEN_1147;
  wire [13:0] _GEN_1149 = 14'h47d == index ? 14'h8 : _GEN_1148;
  wire [13:0] _GEN_1150 = 14'h47e == index ? 14'h8 : _GEN_1149;
  wire [13:0] _GEN_1151 = 14'h47f == index ? 14'h8 : _GEN_1150;
  wire [13:0] _GEN_1152 = 14'h480 == index ? 14'h0 : _GEN_1151;
  wire [13:0] _GEN_1153 = 14'h481 == index ? 14'h480 : _GEN_1152;
  wire [13:0] _GEN_1154 = 14'h482 == index ? 14'h201 : _GEN_1153;
  wire [13:0] _GEN_1155 = 14'h483 == index ? 14'h180 : _GEN_1154;
  wire [13:0] _GEN_1156 = 14'h484 == index ? 14'h101 : _GEN_1155;
  wire [13:0] _GEN_1157 = 14'h485 == index ? 14'h84 : _GEN_1156;
  wire [13:0] _GEN_1158 = 14'h486 == index ? 14'h83 : _GEN_1157;
  wire [13:0] _GEN_1159 = 14'h487 == index ? 14'h82 : _GEN_1158;
  wire [13:0] _GEN_1160 = 14'h488 == index ? 14'h81 : _GEN_1159;
  wire [13:0] _GEN_1161 = 14'h489 == index ? 14'h80 : _GEN_1160;
  wire [13:0] _GEN_1162 = 14'h48a == index ? 14'h9 : _GEN_1161;
  wire [13:0] _GEN_1163 = 14'h48b == index ? 14'h9 : _GEN_1162;
  wire [13:0] _GEN_1164 = 14'h48c == index ? 14'h9 : _GEN_1163;
  wire [13:0] _GEN_1165 = 14'h48d == index ? 14'h9 : _GEN_1164;
  wire [13:0] _GEN_1166 = 14'h48e == index ? 14'h9 : _GEN_1165;
  wire [13:0] _GEN_1167 = 14'h48f == index ? 14'h9 : _GEN_1166;
  wire [13:0] _GEN_1168 = 14'h490 == index ? 14'h9 : _GEN_1167;
  wire [13:0] _GEN_1169 = 14'h491 == index ? 14'h9 : _GEN_1168;
  wire [13:0] _GEN_1170 = 14'h492 == index ? 14'h9 : _GEN_1169;
  wire [13:0] _GEN_1171 = 14'h493 == index ? 14'h9 : _GEN_1170;
  wire [13:0] _GEN_1172 = 14'h494 == index ? 14'h9 : _GEN_1171;
  wire [13:0] _GEN_1173 = 14'h495 == index ? 14'h9 : _GEN_1172;
  wire [13:0] _GEN_1174 = 14'h496 == index ? 14'h9 : _GEN_1173;
  wire [13:0] _GEN_1175 = 14'h497 == index ? 14'h9 : _GEN_1174;
  wire [13:0] _GEN_1176 = 14'h498 == index ? 14'h9 : _GEN_1175;
  wire [13:0] _GEN_1177 = 14'h499 == index ? 14'h9 : _GEN_1176;
  wire [13:0] _GEN_1178 = 14'h49a == index ? 14'h9 : _GEN_1177;
  wire [13:0] _GEN_1179 = 14'h49b == index ? 14'h9 : _GEN_1178;
  wire [13:0] _GEN_1180 = 14'h49c == index ? 14'h9 : _GEN_1179;
  wire [13:0] _GEN_1181 = 14'h49d == index ? 14'h9 : _GEN_1180;
  wire [13:0] _GEN_1182 = 14'h49e == index ? 14'h9 : _GEN_1181;
  wire [13:0] _GEN_1183 = 14'h49f == index ? 14'h9 : _GEN_1182;
  wire [13:0] _GEN_1184 = 14'h4a0 == index ? 14'h9 : _GEN_1183;
  wire [13:0] _GEN_1185 = 14'h4a1 == index ? 14'h9 : _GEN_1184;
  wire [13:0] _GEN_1186 = 14'h4a2 == index ? 14'h9 : _GEN_1185;
  wire [13:0] _GEN_1187 = 14'h4a3 == index ? 14'h9 : _GEN_1186;
  wire [13:0] _GEN_1188 = 14'h4a4 == index ? 14'h9 : _GEN_1187;
  wire [13:0] _GEN_1189 = 14'h4a5 == index ? 14'h9 : _GEN_1188;
  wire [13:0] _GEN_1190 = 14'h4a6 == index ? 14'h9 : _GEN_1189;
  wire [13:0] _GEN_1191 = 14'h4a7 == index ? 14'h9 : _GEN_1190;
  wire [13:0] _GEN_1192 = 14'h4a8 == index ? 14'h9 : _GEN_1191;
  wire [13:0] _GEN_1193 = 14'h4a9 == index ? 14'h9 : _GEN_1192;
  wire [13:0] _GEN_1194 = 14'h4aa == index ? 14'h9 : _GEN_1193;
  wire [13:0] _GEN_1195 = 14'h4ab == index ? 14'h9 : _GEN_1194;
  wire [13:0] _GEN_1196 = 14'h4ac == index ? 14'h9 : _GEN_1195;
  wire [13:0] _GEN_1197 = 14'h4ad == index ? 14'h9 : _GEN_1196;
  wire [13:0] _GEN_1198 = 14'h4ae == index ? 14'h9 : _GEN_1197;
  wire [13:0] _GEN_1199 = 14'h4af == index ? 14'h9 : _GEN_1198;
  wire [13:0] _GEN_1200 = 14'h4b0 == index ? 14'h9 : _GEN_1199;
  wire [13:0] _GEN_1201 = 14'h4b1 == index ? 14'h9 : _GEN_1200;
  wire [13:0] _GEN_1202 = 14'h4b2 == index ? 14'h9 : _GEN_1201;
  wire [13:0] _GEN_1203 = 14'h4b3 == index ? 14'h9 : _GEN_1202;
  wire [13:0] _GEN_1204 = 14'h4b4 == index ? 14'h9 : _GEN_1203;
  wire [13:0] _GEN_1205 = 14'h4b5 == index ? 14'h9 : _GEN_1204;
  wire [13:0] _GEN_1206 = 14'h4b6 == index ? 14'h9 : _GEN_1205;
  wire [13:0] _GEN_1207 = 14'h4b7 == index ? 14'h9 : _GEN_1206;
  wire [13:0] _GEN_1208 = 14'h4b8 == index ? 14'h9 : _GEN_1207;
  wire [13:0] _GEN_1209 = 14'h4b9 == index ? 14'h9 : _GEN_1208;
  wire [13:0] _GEN_1210 = 14'h4ba == index ? 14'h9 : _GEN_1209;
  wire [13:0] _GEN_1211 = 14'h4bb == index ? 14'h9 : _GEN_1210;
  wire [13:0] _GEN_1212 = 14'h4bc == index ? 14'h9 : _GEN_1211;
  wire [13:0] _GEN_1213 = 14'h4bd == index ? 14'h9 : _GEN_1212;
  wire [13:0] _GEN_1214 = 14'h4be == index ? 14'h9 : _GEN_1213;
  wire [13:0] _GEN_1215 = 14'h4bf == index ? 14'h9 : _GEN_1214;
  wire [13:0] _GEN_1216 = 14'h4c0 == index ? 14'h9 : _GEN_1215;
  wire [13:0] _GEN_1217 = 14'h4c1 == index ? 14'h9 : _GEN_1216;
  wire [13:0] _GEN_1218 = 14'h4c2 == index ? 14'h9 : _GEN_1217;
  wire [13:0] _GEN_1219 = 14'h4c3 == index ? 14'h9 : _GEN_1218;
  wire [13:0] _GEN_1220 = 14'h4c4 == index ? 14'h9 : _GEN_1219;
  wire [13:0] _GEN_1221 = 14'h4c5 == index ? 14'h9 : _GEN_1220;
  wire [13:0] _GEN_1222 = 14'h4c6 == index ? 14'h9 : _GEN_1221;
  wire [13:0] _GEN_1223 = 14'h4c7 == index ? 14'h9 : _GEN_1222;
  wire [13:0] _GEN_1224 = 14'h4c8 == index ? 14'h9 : _GEN_1223;
  wire [13:0] _GEN_1225 = 14'h4c9 == index ? 14'h9 : _GEN_1224;
  wire [13:0] _GEN_1226 = 14'h4ca == index ? 14'h9 : _GEN_1225;
  wire [13:0] _GEN_1227 = 14'h4cb == index ? 14'h9 : _GEN_1226;
  wire [13:0] _GEN_1228 = 14'h4cc == index ? 14'h9 : _GEN_1227;
  wire [13:0] _GEN_1229 = 14'h4cd == index ? 14'h9 : _GEN_1228;
  wire [13:0] _GEN_1230 = 14'h4ce == index ? 14'h9 : _GEN_1229;
  wire [13:0] _GEN_1231 = 14'h4cf == index ? 14'h9 : _GEN_1230;
  wire [13:0] _GEN_1232 = 14'h4d0 == index ? 14'h9 : _GEN_1231;
  wire [13:0] _GEN_1233 = 14'h4d1 == index ? 14'h9 : _GEN_1232;
  wire [13:0] _GEN_1234 = 14'h4d2 == index ? 14'h9 : _GEN_1233;
  wire [13:0] _GEN_1235 = 14'h4d3 == index ? 14'h9 : _GEN_1234;
  wire [13:0] _GEN_1236 = 14'h4d4 == index ? 14'h9 : _GEN_1235;
  wire [13:0] _GEN_1237 = 14'h4d5 == index ? 14'h9 : _GEN_1236;
  wire [13:0] _GEN_1238 = 14'h4d6 == index ? 14'h9 : _GEN_1237;
  wire [13:0] _GEN_1239 = 14'h4d7 == index ? 14'h9 : _GEN_1238;
  wire [13:0] _GEN_1240 = 14'h4d8 == index ? 14'h9 : _GEN_1239;
  wire [13:0] _GEN_1241 = 14'h4d9 == index ? 14'h9 : _GEN_1240;
  wire [13:0] _GEN_1242 = 14'h4da == index ? 14'h9 : _GEN_1241;
  wire [13:0] _GEN_1243 = 14'h4db == index ? 14'h9 : _GEN_1242;
  wire [13:0] _GEN_1244 = 14'h4dc == index ? 14'h9 : _GEN_1243;
  wire [13:0] _GEN_1245 = 14'h4dd == index ? 14'h9 : _GEN_1244;
  wire [13:0] _GEN_1246 = 14'h4de == index ? 14'h9 : _GEN_1245;
  wire [13:0] _GEN_1247 = 14'h4df == index ? 14'h9 : _GEN_1246;
  wire [13:0] _GEN_1248 = 14'h4e0 == index ? 14'h9 : _GEN_1247;
  wire [13:0] _GEN_1249 = 14'h4e1 == index ? 14'h9 : _GEN_1248;
  wire [13:0] _GEN_1250 = 14'h4e2 == index ? 14'h9 : _GEN_1249;
  wire [13:0] _GEN_1251 = 14'h4e3 == index ? 14'h9 : _GEN_1250;
  wire [13:0] _GEN_1252 = 14'h4e4 == index ? 14'h9 : _GEN_1251;
  wire [13:0] _GEN_1253 = 14'h4e5 == index ? 14'h9 : _GEN_1252;
  wire [13:0] _GEN_1254 = 14'h4e6 == index ? 14'h9 : _GEN_1253;
  wire [13:0] _GEN_1255 = 14'h4e7 == index ? 14'h9 : _GEN_1254;
  wire [13:0] _GEN_1256 = 14'h4e8 == index ? 14'h9 : _GEN_1255;
  wire [13:0] _GEN_1257 = 14'h4e9 == index ? 14'h9 : _GEN_1256;
  wire [13:0] _GEN_1258 = 14'h4ea == index ? 14'h9 : _GEN_1257;
  wire [13:0] _GEN_1259 = 14'h4eb == index ? 14'h9 : _GEN_1258;
  wire [13:0] _GEN_1260 = 14'h4ec == index ? 14'h9 : _GEN_1259;
  wire [13:0] _GEN_1261 = 14'h4ed == index ? 14'h9 : _GEN_1260;
  wire [13:0] _GEN_1262 = 14'h4ee == index ? 14'h9 : _GEN_1261;
  wire [13:0] _GEN_1263 = 14'h4ef == index ? 14'h9 : _GEN_1262;
  wire [13:0] _GEN_1264 = 14'h4f0 == index ? 14'h9 : _GEN_1263;
  wire [13:0] _GEN_1265 = 14'h4f1 == index ? 14'h9 : _GEN_1264;
  wire [13:0] _GEN_1266 = 14'h4f2 == index ? 14'h9 : _GEN_1265;
  wire [13:0] _GEN_1267 = 14'h4f3 == index ? 14'h9 : _GEN_1266;
  wire [13:0] _GEN_1268 = 14'h4f4 == index ? 14'h9 : _GEN_1267;
  wire [13:0] _GEN_1269 = 14'h4f5 == index ? 14'h9 : _GEN_1268;
  wire [13:0] _GEN_1270 = 14'h4f6 == index ? 14'h9 : _GEN_1269;
  wire [13:0] _GEN_1271 = 14'h4f7 == index ? 14'h9 : _GEN_1270;
  wire [13:0] _GEN_1272 = 14'h4f8 == index ? 14'h9 : _GEN_1271;
  wire [13:0] _GEN_1273 = 14'h4f9 == index ? 14'h9 : _GEN_1272;
  wire [13:0] _GEN_1274 = 14'h4fa == index ? 14'h9 : _GEN_1273;
  wire [13:0] _GEN_1275 = 14'h4fb == index ? 14'h9 : _GEN_1274;
  wire [13:0] _GEN_1276 = 14'h4fc == index ? 14'h9 : _GEN_1275;
  wire [13:0] _GEN_1277 = 14'h4fd == index ? 14'h9 : _GEN_1276;
  wire [13:0] _GEN_1278 = 14'h4fe == index ? 14'h9 : _GEN_1277;
  wire [13:0] _GEN_1279 = 14'h4ff == index ? 14'h9 : _GEN_1278;
  wire [13:0] _GEN_1280 = 14'h500 == index ? 14'h0 : _GEN_1279;
  wire [13:0] _GEN_1281 = 14'h501 == index ? 14'h500 : _GEN_1280;
  wire [13:0] _GEN_1282 = 14'h502 == index ? 14'h280 : _GEN_1281;
  wire [13:0] _GEN_1283 = 14'h503 == index ? 14'h181 : _GEN_1282;
  wire [13:0] _GEN_1284 = 14'h504 == index ? 14'h102 : _GEN_1283;
  wire [13:0] _GEN_1285 = 14'h505 == index ? 14'h100 : _GEN_1284;
  wire [13:0] _GEN_1286 = 14'h506 == index ? 14'h84 : _GEN_1285;
  wire [13:0] _GEN_1287 = 14'h507 == index ? 14'h83 : _GEN_1286;
  wire [13:0] _GEN_1288 = 14'h508 == index ? 14'h82 : _GEN_1287;
  wire [13:0] _GEN_1289 = 14'h509 == index ? 14'h81 : _GEN_1288;
  wire [13:0] _GEN_1290 = 14'h50a == index ? 14'h80 : _GEN_1289;
  wire [13:0] _GEN_1291 = 14'h50b == index ? 14'ha : _GEN_1290;
  wire [13:0] _GEN_1292 = 14'h50c == index ? 14'ha : _GEN_1291;
  wire [13:0] _GEN_1293 = 14'h50d == index ? 14'ha : _GEN_1292;
  wire [13:0] _GEN_1294 = 14'h50e == index ? 14'ha : _GEN_1293;
  wire [13:0] _GEN_1295 = 14'h50f == index ? 14'ha : _GEN_1294;
  wire [13:0] _GEN_1296 = 14'h510 == index ? 14'ha : _GEN_1295;
  wire [13:0] _GEN_1297 = 14'h511 == index ? 14'ha : _GEN_1296;
  wire [13:0] _GEN_1298 = 14'h512 == index ? 14'ha : _GEN_1297;
  wire [13:0] _GEN_1299 = 14'h513 == index ? 14'ha : _GEN_1298;
  wire [13:0] _GEN_1300 = 14'h514 == index ? 14'ha : _GEN_1299;
  wire [13:0] _GEN_1301 = 14'h515 == index ? 14'ha : _GEN_1300;
  wire [13:0] _GEN_1302 = 14'h516 == index ? 14'ha : _GEN_1301;
  wire [13:0] _GEN_1303 = 14'h517 == index ? 14'ha : _GEN_1302;
  wire [13:0] _GEN_1304 = 14'h518 == index ? 14'ha : _GEN_1303;
  wire [13:0] _GEN_1305 = 14'h519 == index ? 14'ha : _GEN_1304;
  wire [13:0] _GEN_1306 = 14'h51a == index ? 14'ha : _GEN_1305;
  wire [13:0] _GEN_1307 = 14'h51b == index ? 14'ha : _GEN_1306;
  wire [13:0] _GEN_1308 = 14'h51c == index ? 14'ha : _GEN_1307;
  wire [13:0] _GEN_1309 = 14'h51d == index ? 14'ha : _GEN_1308;
  wire [13:0] _GEN_1310 = 14'h51e == index ? 14'ha : _GEN_1309;
  wire [13:0] _GEN_1311 = 14'h51f == index ? 14'ha : _GEN_1310;
  wire [13:0] _GEN_1312 = 14'h520 == index ? 14'ha : _GEN_1311;
  wire [13:0] _GEN_1313 = 14'h521 == index ? 14'ha : _GEN_1312;
  wire [13:0] _GEN_1314 = 14'h522 == index ? 14'ha : _GEN_1313;
  wire [13:0] _GEN_1315 = 14'h523 == index ? 14'ha : _GEN_1314;
  wire [13:0] _GEN_1316 = 14'h524 == index ? 14'ha : _GEN_1315;
  wire [13:0] _GEN_1317 = 14'h525 == index ? 14'ha : _GEN_1316;
  wire [13:0] _GEN_1318 = 14'h526 == index ? 14'ha : _GEN_1317;
  wire [13:0] _GEN_1319 = 14'h527 == index ? 14'ha : _GEN_1318;
  wire [13:0] _GEN_1320 = 14'h528 == index ? 14'ha : _GEN_1319;
  wire [13:0] _GEN_1321 = 14'h529 == index ? 14'ha : _GEN_1320;
  wire [13:0] _GEN_1322 = 14'h52a == index ? 14'ha : _GEN_1321;
  wire [13:0] _GEN_1323 = 14'h52b == index ? 14'ha : _GEN_1322;
  wire [13:0] _GEN_1324 = 14'h52c == index ? 14'ha : _GEN_1323;
  wire [13:0] _GEN_1325 = 14'h52d == index ? 14'ha : _GEN_1324;
  wire [13:0] _GEN_1326 = 14'h52e == index ? 14'ha : _GEN_1325;
  wire [13:0] _GEN_1327 = 14'h52f == index ? 14'ha : _GEN_1326;
  wire [13:0] _GEN_1328 = 14'h530 == index ? 14'ha : _GEN_1327;
  wire [13:0] _GEN_1329 = 14'h531 == index ? 14'ha : _GEN_1328;
  wire [13:0] _GEN_1330 = 14'h532 == index ? 14'ha : _GEN_1329;
  wire [13:0] _GEN_1331 = 14'h533 == index ? 14'ha : _GEN_1330;
  wire [13:0] _GEN_1332 = 14'h534 == index ? 14'ha : _GEN_1331;
  wire [13:0] _GEN_1333 = 14'h535 == index ? 14'ha : _GEN_1332;
  wire [13:0] _GEN_1334 = 14'h536 == index ? 14'ha : _GEN_1333;
  wire [13:0] _GEN_1335 = 14'h537 == index ? 14'ha : _GEN_1334;
  wire [13:0] _GEN_1336 = 14'h538 == index ? 14'ha : _GEN_1335;
  wire [13:0] _GEN_1337 = 14'h539 == index ? 14'ha : _GEN_1336;
  wire [13:0] _GEN_1338 = 14'h53a == index ? 14'ha : _GEN_1337;
  wire [13:0] _GEN_1339 = 14'h53b == index ? 14'ha : _GEN_1338;
  wire [13:0] _GEN_1340 = 14'h53c == index ? 14'ha : _GEN_1339;
  wire [13:0] _GEN_1341 = 14'h53d == index ? 14'ha : _GEN_1340;
  wire [13:0] _GEN_1342 = 14'h53e == index ? 14'ha : _GEN_1341;
  wire [13:0] _GEN_1343 = 14'h53f == index ? 14'ha : _GEN_1342;
  wire [13:0] _GEN_1344 = 14'h540 == index ? 14'ha : _GEN_1343;
  wire [13:0] _GEN_1345 = 14'h541 == index ? 14'ha : _GEN_1344;
  wire [13:0] _GEN_1346 = 14'h542 == index ? 14'ha : _GEN_1345;
  wire [13:0] _GEN_1347 = 14'h543 == index ? 14'ha : _GEN_1346;
  wire [13:0] _GEN_1348 = 14'h544 == index ? 14'ha : _GEN_1347;
  wire [13:0] _GEN_1349 = 14'h545 == index ? 14'ha : _GEN_1348;
  wire [13:0] _GEN_1350 = 14'h546 == index ? 14'ha : _GEN_1349;
  wire [13:0] _GEN_1351 = 14'h547 == index ? 14'ha : _GEN_1350;
  wire [13:0] _GEN_1352 = 14'h548 == index ? 14'ha : _GEN_1351;
  wire [13:0] _GEN_1353 = 14'h549 == index ? 14'ha : _GEN_1352;
  wire [13:0] _GEN_1354 = 14'h54a == index ? 14'ha : _GEN_1353;
  wire [13:0] _GEN_1355 = 14'h54b == index ? 14'ha : _GEN_1354;
  wire [13:0] _GEN_1356 = 14'h54c == index ? 14'ha : _GEN_1355;
  wire [13:0] _GEN_1357 = 14'h54d == index ? 14'ha : _GEN_1356;
  wire [13:0] _GEN_1358 = 14'h54e == index ? 14'ha : _GEN_1357;
  wire [13:0] _GEN_1359 = 14'h54f == index ? 14'ha : _GEN_1358;
  wire [13:0] _GEN_1360 = 14'h550 == index ? 14'ha : _GEN_1359;
  wire [13:0] _GEN_1361 = 14'h551 == index ? 14'ha : _GEN_1360;
  wire [13:0] _GEN_1362 = 14'h552 == index ? 14'ha : _GEN_1361;
  wire [13:0] _GEN_1363 = 14'h553 == index ? 14'ha : _GEN_1362;
  wire [13:0] _GEN_1364 = 14'h554 == index ? 14'ha : _GEN_1363;
  wire [13:0] _GEN_1365 = 14'h555 == index ? 14'ha : _GEN_1364;
  wire [13:0] _GEN_1366 = 14'h556 == index ? 14'ha : _GEN_1365;
  wire [13:0] _GEN_1367 = 14'h557 == index ? 14'ha : _GEN_1366;
  wire [13:0] _GEN_1368 = 14'h558 == index ? 14'ha : _GEN_1367;
  wire [13:0] _GEN_1369 = 14'h559 == index ? 14'ha : _GEN_1368;
  wire [13:0] _GEN_1370 = 14'h55a == index ? 14'ha : _GEN_1369;
  wire [13:0] _GEN_1371 = 14'h55b == index ? 14'ha : _GEN_1370;
  wire [13:0] _GEN_1372 = 14'h55c == index ? 14'ha : _GEN_1371;
  wire [13:0] _GEN_1373 = 14'h55d == index ? 14'ha : _GEN_1372;
  wire [13:0] _GEN_1374 = 14'h55e == index ? 14'ha : _GEN_1373;
  wire [13:0] _GEN_1375 = 14'h55f == index ? 14'ha : _GEN_1374;
  wire [13:0] _GEN_1376 = 14'h560 == index ? 14'ha : _GEN_1375;
  wire [13:0] _GEN_1377 = 14'h561 == index ? 14'ha : _GEN_1376;
  wire [13:0] _GEN_1378 = 14'h562 == index ? 14'ha : _GEN_1377;
  wire [13:0] _GEN_1379 = 14'h563 == index ? 14'ha : _GEN_1378;
  wire [13:0] _GEN_1380 = 14'h564 == index ? 14'ha : _GEN_1379;
  wire [13:0] _GEN_1381 = 14'h565 == index ? 14'ha : _GEN_1380;
  wire [13:0] _GEN_1382 = 14'h566 == index ? 14'ha : _GEN_1381;
  wire [13:0] _GEN_1383 = 14'h567 == index ? 14'ha : _GEN_1382;
  wire [13:0] _GEN_1384 = 14'h568 == index ? 14'ha : _GEN_1383;
  wire [13:0] _GEN_1385 = 14'h569 == index ? 14'ha : _GEN_1384;
  wire [13:0] _GEN_1386 = 14'h56a == index ? 14'ha : _GEN_1385;
  wire [13:0] _GEN_1387 = 14'h56b == index ? 14'ha : _GEN_1386;
  wire [13:0] _GEN_1388 = 14'h56c == index ? 14'ha : _GEN_1387;
  wire [13:0] _GEN_1389 = 14'h56d == index ? 14'ha : _GEN_1388;
  wire [13:0] _GEN_1390 = 14'h56e == index ? 14'ha : _GEN_1389;
  wire [13:0] _GEN_1391 = 14'h56f == index ? 14'ha : _GEN_1390;
  wire [13:0] _GEN_1392 = 14'h570 == index ? 14'ha : _GEN_1391;
  wire [13:0] _GEN_1393 = 14'h571 == index ? 14'ha : _GEN_1392;
  wire [13:0] _GEN_1394 = 14'h572 == index ? 14'ha : _GEN_1393;
  wire [13:0] _GEN_1395 = 14'h573 == index ? 14'ha : _GEN_1394;
  wire [13:0] _GEN_1396 = 14'h574 == index ? 14'ha : _GEN_1395;
  wire [13:0] _GEN_1397 = 14'h575 == index ? 14'ha : _GEN_1396;
  wire [13:0] _GEN_1398 = 14'h576 == index ? 14'ha : _GEN_1397;
  wire [13:0] _GEN_1399 = 14'h577 == index ? 14'ha : _GEN_1398;
  wire [13:0] _GEN_1400 = 14'h578 == index ? 14'ha : _GEN_1399;
  wire [13:0] _GEN_1401 = 14'h579 == index ? 14'ha : _GEN_1400;
  wire [13:0] _GEN_1402 = 14'h57a == index ? 14'ha : _GEN_1401;
  wire [13:0] _GEN_1403 = 14'h57b == index ? 14'ha : _GEN_1402;
  wire [13:0] _GEN_1404 = 14'h57c == index ? 14'ha : _GEN_1403;
  wire [13:0] _GEN_1405 = 14'h57d == index ? 14'ha : _GEN_1404;
  wire [13:0] _GEN_1406 = 14'h57e == index ? 14'ha : _GEN_1405;
  wire [13:0] _GEN_1407 = 14'h57f == index ? 14'ha : _GEN_1406;
  wire [13:0] _GEN_1408 = 14'h580 == index ? 14'h0 : _GEN_1407;
  wire [13:0] _GEN_1409 = 14'h581 == index ? 14'h580 : _GEN_1408;
  wire [13:0] _GEN_1410 = 14'h582 == index ? 14'h281 : _GEN_1409;
  wire [13:0] _GEN_1411 = 14'h583 == index ? 14'h182 : _GEN_1410;
  wire [13:0] _GEN_1412 = 14'h584 == index ? 14'h103 : _GEN_1411;
  wire [13:0] _GEN_1413 = 14'h585 == index ? 14'h101 : _GEN_1412;
  wire [13:0] _GEN_1414 = 14'h586 == index ? 14'h85 : _GEN_1413;
  wire [13:0] _GEN_1415 = 14'h587 == index ? 14'h84 : _GEN_1414;
  wire [13:0] _GEN_1416 = 14'h588 == index ? 14'h83 : _GEN_1415;
  wire [13:0] _GEN_1417 = 14'h589 == index ? 14'h82 : _GEN_1416;
  wire [13:0] _GEN_1418 = 14'h58a == index ? 14'h81 : _GEN_1417;
  wire [13:0] _GEN_1419 = 14'h58b == index ? 14'h80 : _GEN_1418;
  wire [13:0] _GEN_1420 = 14'h58c == index ? 14'hb : _GEN_1419;
  wire [13:0] _GEN_1421 = 14'h58d == index ? 14'hb : _GEN_1420;
  wire [13:0] _GEN_1422 = 14'h58e == index ? 14'hb : _GEN_1421;
  wire [13:0] _GEN_1423 = 14'h58f == index ? 14'hb : _GEN_1422;
  wire [13:0] _GEN_1424 = 14'h590 == index ? 14'hb : _GEN_1423;
  wire [13:0] _GEN_1425 = 14'h591 == index ? 14'hb : _GEN_1424;
  wire [13:0] _GEN_1426 = 14'h592 == index ? 14'hb : _GEN_1425;
  wire [13:0] _GEN_1427 = 14'h593 == index ? 14'hb : _GEN_1426;
  wire [13:0] _GEN_1428 = 14'h594 == index ? 14'hb : _GEN_1427;
  wire [13:0] _GEN_1429 = 14'h595 == index ? 14'hb : _GEN_1428;
  wire [13:0] _GEN_1430 = 14'h596 == index ? 14'hb : _GEN_1429;
  wire [13:0] _GEN_1431 = 14'h597 == index ? 14'hb : _GEN_1430;
  wire [13:0] _GEN_1432 = 14'h598 == index ? 14'hb : _GEN_1431;
  wire [13:0] _GEN_1433 = 14'h599 == index ? 14'hb : _GEN_1432;
  wire [13:0] _GEN_1434 = 14'h59a == index ? 14'hb : _GEN_1433;
  wire [13:0] _GEN_1435 = 14'h59b == index ? 14'hb : _GEN_1434;
  wire [13:0] _GEN_1436 = 14'h59c == index ? 14'hb : _GEN_1435;
  wire [13:0] _GEN_1437 = 14'h59d == index ? 14'hb : _GEN_1436;
  wire [13:0] _GEN_1438 = 14'h59e == index ? 14'hb : _GEN_1437;
  wire [13:0] _GEN_1439 = 14'h59f == index ? 14'hb : _GEN_1438;
  wire [13:0] _GEN_1440 = 14'h5a0 == index ? 14'hb : _GEN_1439;
  wire [13:0] _GEN_1441 = 14'h5a1 == index ? 14'hb : _GEN_1440;
  wire [13:0] _GEN_1442 = 14'h5a2 == index ? 14'hb : _GEN_1441;
  wire [13:0] _GEN_1443 = 14'h5a3 == index ? 14'hb : _GEN_1442;
  wire [13:0] _GEN_1444 = 14'h5a4 == index ? 14'hb : _GEN_1443;
  wire [13:0] _GEN_1445 = 14'h5a5 == index ? 14'hb : _GEN_1444;
  wire [13:0] _GEN_1446 = 14'h5a6 == index ? 14'hb : _GEN_1445;
  wire [13:0] _GEN_1447 = 14'h5a7 == index ? 14'hb : _GEN_1446;
  wire [13:0] _GEN_1448 = 14'h5a8 == index ? 14'hb : _GEN_1447;
  wire [13:0] _GEN_1449 = 14'h5a9 == index ? 14'hb : _GEN_1448;
  wire [13:0] _GEN_1450 = 14'h5aa == index ? 14'hb : _GEN_1449;
  wire [13:0] _GEN_1451 = 14'h5ab == index ? 14'hb : _GEN_1450;
  wire [13:0] _GEN_1452 = 14'h5ac == index ? 14'hb : _GEN_1451;
  wire [13:0] _GEN_1453 = 14'h5ad == index ? 14'hb : _GEN_1452;
  wire [13:0] _GEN_1454 = 14'h5ae == index ? 14'hb : _GEN_1453;
  wire [13:0] _GEN_1455 = 14'h5af == index ? 14'hb : _GEN_1454;
  wire [13:0] _GEN_1456 = 14'h5b0 == index ? 14'hb : _GEN_1455;
  wire [13:0] _GEN_1457 = 14'h5b1 == index ? 14'hb : _GEN_1456;
  wire [13:0] _GEN_1458 = 14'h5b2 == index ? 14'hb : _GEN_1457;
  wire [13:0] _GEN_1459 = 14'h5b3 == index ? 14'hb : _GEN_1458;
  wire [13:0] _GEN_1460 = 14'h5b4 == index ? 14'hb : _GEN_1459;
  wire [13:0] _GEN_1461 = 14'h5b5 == index ? 14'hb : _GEN_1460;
  wire [13:0] _GEN_1462 = 14'h5b6 == index ? 14'hb : _GEN_1461;
  wire [13:0] _GEN_1463 = 14'h5b7 == index ? 14'hb : _GEN_1462;
  wire [13:0] _GEN_1464 = 14'h5b8 == index ? 14'hb : _GEN_1463;
  wire [13:0] _GEN_1465 = 14'h5b9 == index ? 14'hb : _GEN_1464;
  wire [13:0] _GEN_1466 = 14'h5ba == index ? 14'hb : _GEN_1465;
  wire [13:0] _GEN_1467 = 14'h5bb == index ? 14'hb : _GEN_1466;
  wire [13:0] _GEN_1468 = 14'h5bc == index ? 14'hb : _GEN_1467;
  wire [13:0] _GEN_1469 = 14'h5bd == index ? 14'hb : _GEN_1468;
  wire [13:0] _GEN_1470 = 14'h5be == index ? 14'hb : _GEN_1469;
  wire [13:0] _GEN_1471 = 14'h5bf == index ? 14'hb : _GEN_1470;
  wire [13:0] _GEN_1472 = 14'h5c0 == index ? 14'hb : _GEN_1471;
  wire [13:0] _GEN_1473 = 14'h5c1 == index ? 14'hb : _GEN_1472;
  wire [13:0] _GEN_1474 = 14'h5c2 == index ? 14'hb : _GEN_1473;
  wire [13:0] _GEN_1475 = 14'h5c3 == index ? 14'hb : _GEN_1474;
  wire [13:0] _GEN_1476 = 14'h5c4 == index ? 14'hb : _GEN_1475;
  wire [13:0] _GEN_1477 = 14'h5c5 == index ? 14'hb : _GEN_1476;
  wire [13:0] _GEN_1478 = 14'h5c6 == index ? 14'hb : _GEN_1477;
  wire [13:0] _GEN_1479 = 14'h5c7 == index ? 14'hb : _GEN_1478;
  wire [13:0] _GEN_1480 = 14'h5c8 == index ? 14'hb : _GEN_1479;
  wire [13:0] _GEN_1481 = 14'h5c9 == index ? 14'hb : _GEN_1480;
  wire [13:0] _GEN_1482 = 14'h5ca == index ? 14'hb : _GEN_1481;
  wire [13:0] _GEN_1483 = 14'h5cb == index ? 14'hb : _GEN_1482;
  wire [13:0] _GEN_1484 = 14'h5cc == index ? 14'hb : _GEN_1483;
  wire [13:0] _GEN_1485 = 14'h5cd == index ? 14'hb : _GEN_1484;
  wire [13:0] _GEN_1486 = 14'h5ce == index ? 14'hb : _GEN_1485;
  wire [13:0] _GEN_1487 = 14'h5cf == index ? 14'hb : _GEN_1486;
  wire [13:0] _GEN_1488 = 14'h5d0 == index ? 14'hb : _GEN_1487;
  wire [13:0] _GEN_1489 = 14'h5d1 == index ? 14'hb : _GEN_1488;
  wire [13:0] _GEN_1490 = 14'h5d2 == index ? 14'hb : _GEN_1489;
  wire [13:0] _GEN_1491 = 14'h5d3 == index ? 14'hb : _GEN_1490;
  wire [13:0] _GEN_1492 = 14'h5d4 == index ? 14'hb : _GEN_1491;
  wire [13:0] _GEN_1493 = 14'h5d5 == index ? 14'hb : _GEN_1492;
  wire [13:0] _GEN_1494 = 14'h5d6 == index ? 14'hb : _GEN_1493;
  wire [13:0] _GEN_1495 = 14'h5d7 == index ? 14'hb : _GEN_1494;
  wire [13:0] _GEN_1496 = 14'h5d8 == index ? 14'hb : _GEN_1495;
  wire [13:0] _GEN_1497 = 14'h5d9 == index ? 14'hb : _GEN_1496;
  wire [13:0] _GEN_1498 = 14'h5da == index ? 14'hb : _GEN_1497;
  wire [13:0] _GEN_1499 = 14'h5db == index ? 14'hb : _GEN_1498;
  wire [13:0] _GEN_1500 = 14'h5dc == index ? 14'hb : _GEN_1499;
  wire [13:0] _GEN_1501 = 14'h5dd == index ? 14'hb : _GEN_1500;
  wire [13:0] _GEN_1502 = 14'h5de == index ? 14'hb : _GEN_1501;
  wire [13:0] _GEN_1503 = 14'h5df == index ? 14'hb : _GEN_1502;
  wire [13:0] _GEN_1504 = 14'h5e0 == index ? 14'hb : _GEN_1503;
  wire [13:0] _GEN_1505 = 14'h5e1 == index ? 14'hb : _GEN_1504;
  wire [13:0] _GEN_1506 = 14'h5e2 == index ? 14'hb : _GEN_1505;
  wire [13:0] _GEN_1507 = 14'h5e3 == index ? 14'hb : _GEN_1506;
  wire [13:0] _GEN_1508 = 14'h5e4 == index ? 14'hb : _GEN_1507;
  wire [13:0] _GEN_1509 = 14'h5e5 == index ? 14'hb : _GEN_1508;
  wire [13:0] _GEN_1510 = 14'h5e6 == index ? 14'hb : _GEN_1509;
  wire [13:0] _GEN_1511 = 14'h5e7 == index ? 14'hb : _GEN_1510;
  wire [13:0] _GEN_1512 = 14'h5e8 == index ? 14'hb : _GEN_1511;
  wire [13:0] _GEN_1513 = 14'h5e9 == index ? 14'hb : _GEN_1512;
  wire [13:0] _GEN_1514 = 14'h5ea == index ? 14'hb : _GEN_1513;
  wire [13:0] _GEN_1515 = 14'h5eb == index ? 14'hb : _GEN_1514;
  wire [13:0] _GEN_1516 = 14'h5ec == index ? 14'hb : _GEN_1515;
  wire [13:0] _GEN_1517 = 14'h5ed == index ? 14'hb : _GEN_1516;
  wire [13:0] _GEN_1518 = 14'h5ee == index ? 14'hb : _GEN_1517;
  wire [13:0] _GEN_1519 = 14'h5ef == index ? 14'hb : _GEN_1518;
  wire [13:0] _GEN_1520 = 14'h5f0 == index ? 14'hb : _GEN_1519;
  wire [13:0] _GEN_1521 = 14'h5f1 == index ? 14'hb : _GEN_1520;
  wire [13:0] _GEN_1522 = 14'h5f2 == index ? 14'hb : _GEN_1521;
  wire [13:0] _GEN_1523 = 14'h5f3 == index ? 14'hb : _GEN_1522;
  wire [13:0] _GEN_1524 = 14'h5f4 == index ? 14'hb : _GEN_1523;
  wire [13:0] _GEN_1525 = 14'h5f5 == index ? 14'hb : _GEN_1524;
  wire [13:0] _GEN_1526 = 14'h5f6 == index ? 14'hb : _GEN_1525;
  wire [13:0] _GEN_1527 = 14'h5f7 == index ? 14'hb : _GEN_1526;
  wire [13:0] _GEN_1528 = 14'h5f8 == index ? 14'hb : _GEN_1527;
  wire [13:0] _GEN_1529 = 14'h5f9 == index ? 14'hb : _GEN_1528;
  wire [13:0] _GEN_1530 = 14'h5fa == index ? 14'hb : _GEN_1529;
  wire [13:0] _GEN_1531 = 14'h5fb == index ? 14'hb : _GEN_1530;
  wire [13:0] _GEN_1532 = 14'h5fc == index ? 14'hb : _GEN_1531;
  wire [13:0] _GEN_1533 = 14'h5fd == index ? 14'hb : _GEN_1532;
  wire [13:0] _GEN_1534 = 14'h5fe == index ? 14'hb : _GEN_1533;
  wire [13:0] _GEN_1535 = 14'h5ff == index ? 14'hb : _GEN_1534;
  wire [13:0] _GEN_1536 = 14'h600 == index ? 14'h0 : _GEN_1535;
  wire [13:0] _GEN_1537 = 14'h601 == index ? 14'h600 : _GEN_1536;
  wire [13:0] _GEN_1538 = 14'h602 == index ? 14'h300 : _GEN_1537;
  wire [13:0] _GEN_1539 = 14'h603 == index ? 14'h200 : _GEN_1538;
  wire [13:0] _GEN_1540 = 14'h604 == index ? 14'h180 : _GEN_1539;
  wire [13:0] _GEN_1541 = 14'h605 == index ? 14'h102 : _GEN_1540;
  wire [13:0] _GEN_1542 = 14'h606 == index ? 14'h100 : _GEN_1541;
  wire [13:0] _GEN_1543 = 14'h607 == index ? 14'h85 : _GEN_1542;
  wire [13:0] _GEN_1544 = 14'h608 == index ? 14'h84 : _GEN_1543;
  wire [13:0] _GEN_1545 = 14'h609 == index ? 14'h83 : _GEN_1544;
  wire [13:0] _GEN_1546 = 14'h60a == index ? 14'h82 : _GEN_1545;
  wire [13:0] _GEN_1547 = 14'h60b == index ? 14'h81 : _GEN_1546;
  wire [13:0] _GEN_1548 = 14'h60c == index ? 14'h80 : _GEN_1547;
  wire [13:0] _GEN_1549 = 14'h60d == index ? 14'hc : _GEN_1548;
  wire [13:0] _GEN_1550 = 14'h60e == index ? 14'hc : _GEN_1549;
  wire [13:0] _GEN_1551 = 14'h60f == index ? 14'hc : _GEN_1550;
  wire [13:0] _GEN_1552 = 14'h610 == index ? 14'hc : _GEN_1551;
  wire [13:0] _GEN_1553 = 14'h611 == index ? 14'hc : _GEN_1552;
  wire [13:0] _GEN_1554 = 14'h612 == index ? 14'hc : _GEN_1553;
  wire [13:0] _GEN_1555 = 14'h613 == index ? 14'hc : _GEN_1554;
  wire [13:0] _GEN_1556 = 14'h614 == index ? 14'hc : _GEN_1555;
  wire [13:0] _GEN_1557 = 14'h615 == index ? 14'hc : _GEN_1556;
  wire [13:0] _GEN_1558 = 14'h616 == index ? 14'hc : _GEN_1557;
  wire [13:0] _GEN_1559 = 14'h617 == index ? 14'hc : _GEN_1558;
  wire [13:0] _GEN_1560 = 14'h618 == index ? 14'hc : _GEN_1559;
  wire [13:0] _GEN_1561 = 14'h619 == index ? 14'hc : _GEN_1560;
  wire [13:0] _GEN_1562 = 14'h61a == index ? 14'hc : _GEN_1561;
  wire [13:0] _GEN_1563 = 14'h61b == index ? 14'hc : _GEN_1562;
  wire [13:0] _GEN_1564 = 14'h61c == index ? 14'hc : _GEN_1563;
  wire [13:0] _GEN_1565 = 14'h61d == index ? 14'hc : _GEN_1564;
  wire [13:0] _GEN_1566 = 14'h61e == index ? 14'hc : _GEN_1565;
  wire [13:0] _GEN_1567 = 14'h61f == index ? 14'hc : _GEN_1566;
  wire [13:0] _GEN_1568 = 14'h620 == index ? 14'hc : _GEN_1567;
  wire [13:0] _GEN_1569 = 14'h621 == index ? 14'hc : _GEN_1568;
  wire [13:0] _GEN_1570 = 14'h622 == index ? 14'hc : _GEN_1569;
  wire [13:0] _GEN_1571 = 14'h623 == index ? 14'hc : _GEN_1570;
  wire [13:0] _GEN_1572 = 14'h624 == index ? 14'hc : _GEN_1571;
  wire [13:0] _GEN_1573 = 14'h625 == index ? 14'hc : _GEN_1572;
  wire [13:0] _GEN_1574 = 14'h626 == index ? 14'hc : _GEN_1573;
  wire [13:0] _GEN_1575 = 14'h627 == index ? 14'hc : _GEN_1574;
  wire [13:0] _GEN_1576 = 14'h628 == index ? 14'hc : _GEN_1575;
  wire [13:0] _GEN_1577 = 14'h629 == index ? 14'hc : _GEN_1576;
  wire [13:0] _GEN_1578 = 14'h62a == index ? 14'hc : _GEN_1577;
  wire [13:0] _GEN_1579 = 14'h62b == index ? 14'hc : _GEN_1578;
  wire [13:0] _GEN_1580 = 14'h62c == index ? 14'hc : _GEN_1579;
  wire [13:0] _GEN_1581 = 14'h62d == index ? 14'hc : _GEN_1580;
  wire [13:0] _GEN_1582 = 14'h62e == index ? 14'hc : _GEN_1581;
  wire [13:0] _GEN_1583 = 14'h62f == index ? 14'hc : _GEN_1582;
  wire [13:0] _GEN_1584 = 14'h630 == index ? 14'hc : _GEN_1583;
  wire [13:0] _GEN_1585 = 14'h631 == index ? 14'hc : _GEN_1584;
  wire [13:0] _GEN_1586 = 14'h632 == index ? 14'hc : _GEN_1585;
  wire [13:0] _GEN_1587 = 14'h633 == index ? 14'hc : _GEN_1586;
  wire [13:0] _GEN_1588 = 14'h634 == index ? 14'hc : _GEN_1587;
  wire [13:0] _GEN_1589 = 14'h635 == index ? 14'hc : _GEN_1588;
  wire [13:0] _GEN_1590 = 14'h636 == index ? 14'hc : _GEN_1589;
  wire [13:0] _GEN_1591 = 14'h637 == index ? 14'hc : _GEN_1590;
  wire [13:0] _GEN_1592 = 14'h638 == index ? 14'hc : _GEN_1591;
  wire [13:0] _GEN_1593 = 14'h639 == index ? 14'hc : _GEN_1592;
  wire [13:0] _GEN_1594 = 14'h63a == index ? 14'hc : _GEN_1593;
  wire [13:0] _GEN_1595 = 14'h63b == index ? 14'hc : _GEN_1594;
  wire [13:0] _GEN_1596 = 14'h63c == index ? 14'hc : _GEN_1595;
  wire [13:0] _GEN_1597 = 14'h63d == index ? 14'hc : _GEN_1596;
  wire [13:0] _GEN_1598 = 14'h63e == index ? 14'hc : _GEN_1597;
  wire [13:0] _GEN_1599 = 14'h63f == index ? 14'hc : _GEN_1598;
  wire [13:0] _GEN_1600 = 14'h640 == index ? 14'hc : _GEN_1599;
  wire [13:0] _GEN_1601 = 14'h641 == index ? 14'hc : _GEN_1600;
  wire [13:0] _GEN_1602 = 14'h642 == index ? 14'hc : _GEN_1601;
  wire [13:0] _GEN_1603 = 14'h643 == index ? 14'hc : _GEN_1602;
  wire [13:0] _GEN_1604 = 14'h644 == index ? 14'hc : _GEN_1603;
  wire [13:0] _GEN_1605 = 14'h645 == index ? 14'hc : _GEN_1604;
  wire [13:0] _GEN_1606 = 14'h646 == index ? 14'hc : _GEN_1605;
  wire [13:0] _GEN_1607 = 14'h647 == index ? 14'hc : _GEN_1606;
  wire [13:0] _GEN_1608 = 14'h648 == index ? 14'hc : _GEN_1607;
  wire [13:0] _GEN_1609 = 14'h649 == index ? 14'hc : _GEN_1608;
  wire [13:0] _GEN_1610 = 14'h64a == index ? 14'hc : _GEN_1609;
  wire [13:0] _GEN_1611 = 14'h64b == index ? 14'hc : _GEN_1610;
  wire [13:0] _GEN_1612 = 14'h64c == index ? 14'hc : _GEN_1611;
  wire [13:0] _GEN_1613 = 14'h64d == index ? 14'hc : _GEN_1612;
  wire [13:0] _GEN_1614 = 14'h64e == index ? 14'hc : _GEN_1613;
  wire [13:0] _GEN_1615 = 14'h64f == index ? 14'hc : _GEN_1614;
  wire [13:0] _GEN_1616 = 14'h650 == index ? 14'hc : _GEN_1615;
  wire [13:0] _GEN_1617 = 14'h651 == index ? 14'hc : _GEN_1616;
  wire [13:0] _GEN_1618 = 14'h652 == index ? 14'hc : _GEN_1617;
  wire [13:0] _GEN_1619 = 14'h653 == index ? 14'hc : _GEN_1618;
  wire [13:0] _GEN_1620 = 14'h654 == index ? 14'hc : _GEN_1619;
  wire [13:0] _GEN_1621 = 14'h655 == index ? 14'hc : _GEN_1620;
  wire [13:0] _GEN_1622 = 14'h656 == index ? 14'hc : _GEN_1621;
  wire [13:0] _GEN_1623 = 14'h657 == index ? 14'hc : _GEN_1622;
  wire [13:0] _GEN_1624 = 14'h658 == index ? 14'hc : _GEN_1623;
  wire [13:0] _GEN_1625 = 14'h659 == index ? 14'hc : _GEN_1624;
  wire [13:0] _GEN_1626 = 14'h65a == index ? 14'hc : _GEN_1625;
  wire [13:0] _GEN_1627 = 14'h65b == index ? 14'hc : _GEN_1626;
  wire [13:0] _GEN_1628 = 14'h65c == index ? 14'hc : _GEN_1627;
  wire [13:0] _GEN_1629 = 14'h65d == index ? 14'hc : _GEN_1628;
  wire [13:0] _GEN_1630 = 14'h65e == index ? 14'hc : _GEN_1629;
  wire [13:0] _GEN_1631 = 14'h65f == index ? 14'hc : _GEN_1630;
  wire [13:0] _GEN_1632 = 14'h660 == index ? 14'hc : _GEN_1631;
  wire [13:0] _GEN_1633 = 14'h661 == index ? 14'hc : _GEN_1632;
  wire [13:0] _GEN_1634 = 14'h662 == index ? 14'hc : _GEN_1633;
  wire [13:0] _GEN_1635 = 14'h663 == index ? 14'hc : _GEN_1634;
  wire [13:0] _GEN_1636 = 14'h664 == index ? 14'hc : _GEN_1635;
  wire [13:0] _GEN_1637 = 14'h665 == index ? 14'hc : _GEN_1636;
  wire [13:0] _GEN_1638 = 14'h666 == index ? 14'hc : _GEN_1637;
  wire [13:0] _GEN_1639 = 14'h667 == index ? 14'hc : _GEN_1638;
  wire [13:0] _GEN_1640 = 14'h668 == index ? 14'hc : _GEN_1639;
  wire [13:0] _GEN_1641 = 14'h669 == index ? 14'hc : _GEN_1640;
  wire [13:0] _GEN_1642 = 14'h66a == index ? 14'hc : _GEN_1641;
  wire [13:0] _GEN_1643 = 14'h66b == index ? 14'hc : _GEN_1642;
  wire [13:0] _GEN_1644 = 14'h66c == index ? 14'hc : _GEN_1643;
  wire [13:0] _GEN_1645 = 14'h66d == index ? 14'hc : _GEN_1644;
  wire [13:0] _GEN_1646 = 14'h66e == index ? 14'hc : _GEN_1645;
  wire [13:0] _GEN_1647 = 14'h66f == index ? 14'hc : _GEN_1646;
  wire [13:0] _GEN_1648 = 14'h670 == index ? 14'hc : _GEN_1647;
  wire [13:0] _GEN_1649 = 14'h671 == index ? 14'hc : _GEN_1648;
  wire [13:0] _GEN_1650 = 14'h672 == index ? 14'hc : _GEN_1649;
  wire [13:0] _GEN_1651 = 14'h673 == index ? 14'hc : _GEN_1650;
  wire [13:0] _GEN_1652 = 14'h674 == index ? 14'hc : _GEN_1651;
  wire [13:0] _GEN_1653 = 14'h675 == index ? 14'hc : _GEN_1652;
  wire [13:0] _GEN_1654 = 14'h676 == index ? 14'hc : _GEN_1653;
  wire [13:0] _GEN_1655 = 14'h677 == index ? 14'hc : _GEN_1654;
  wire [13:0] _GEN_1656 = 14'h678 == index ? 14'hc : _GEN_1655;
  wire [13:0] _GEN_1657 = 14'h679 == index ? 14'hc : _GEN_1656;
  wire [13:0] _GEN_1658 = 14'h67a == index ? 14'hc : _GEN_1657;
  wire [13:0] _GEN_1659 = 14'h67b == index ? 14'hc : _GEN_1658;
  wire [13:0] _GEN_1660 = 14'h67c == index ? 14'hc : _GEN_1659;
  wire [13:0] _GEN_1661 = 14'h67d == index ? 14'hc : _GEN_1660;
  wire [13:0] _GEN_1662 = 14'h67e == index ? 14'hc : _GEN_1661;
  wire [13:0] _GEN_1663 = 14'h67f == index ? 14'hc : _GEN_1662;
  wire [13:0] _GEN_1664 = 14'h680 == index ? 14'h0 : _GEN_1663;
  wire [13:0] _GEN_1665 = 14'h681 == index ? 14'h680 : _GEN_1664;
  wire [13:0] _GEN_1666 = 14'h682 == index ? 14'h301 : _GEN_1665;
  wire [13:0] _GEN_1667 = 14'h683 == index ? 14'h201 : _GEN_1666;
  wire [13:0] _GEN_1668 = 14'h684 == index ? 14'h181 : _GEN_1667;
  wire [13:0] _GEN_1669 = 14'h685 == index ? 14'h103 : _GEN_1668;
  wire [13:0] _GEN_1670 = 14'h686 == index ? 14'h101 : _GEN_1669;
  wire [13:0] _GEN_1671 = 14'h687 == index ? 14'h86 : _GEN_1670;
  wire [13:0] _GEN_1672 = 14'h688 == index ? 14'h85 : _GEN_1671;
  wire [13:0] _GEN_1673 = 14'h689 == index ? 14'h84 : _GEN_1672;
  wire [13:0] _GEN_1674 = 14'h68a == index ? 14'h83 : _GEN_1673;
  wire [13:0] _GEN_1675 = 14'h68b == index ? 14'h82 : _GEN_1674;
  wire [13:0] _GEN_1676 = 14'h68c == index ? 14'h81 : _GEN_1675;
  wire [13:0] _GEN_1677 = 14'h68d == index ? 14'h80 : _GEN_1676;
  wire [13:0] _GEN_1678 = 14'h68e == index ? 14'hd : _GEN_1677;
  wire [13:0] _GEN_1679 = 14'h68f == index ? 14'hd : _GEN_1678;
  wire [13:0] _GEN_1680 = 14'h690 == index ? 14'hd : _GEN_1679;
  wire [13:0] _GEN_1681 = 14'h691 == index ? 14'hd : _GEN_1680;
  wire [13:0] _GEN_1682 = 14'h692 == index ? 14'hd : _GEN_1681;
  wire [13:0] _GEN_1683 = 14'h693 == index ? 14'hd : _GEN_1682;
  wire [13:0] _GEN_1684 = 14'h694 == index ? 14'hd : _GEN_1683;
  wire [13:0] _GEN_1685 = 14'h695 == index ? 14'hd : _GEN_1684;
  wire [13:0] _GEN_1686 = 14'h696 == index ? 14'hd : _GEN_1685;
  wire [13:0] _GEN_1687 = 14'h697 == index ? 14'hd : _GEN_1686;
  wire [13:0] _GEN_1688 = 14'h698 == index ? 14'hd : _GEN_1687;
  wire [13:0] _GEN_1689 = 14'h699 == index ? 14'hd : _GEN_1688;
  wire [13:0] _GEN_1690 = 14'h69a == index ? 14'hd : _GEN_1689;
  wire [13:0] _GEN_1691 = 14'h69b == index ? 14'hd : _GEN_1690;
  wire [13:0] _GEN_1692 = 14'h69c == index ? 14'hd : _GEN_1691;
  wire [13:0] _GEN_1693 = 14'h69d == index ? 14'hd : _GEN_1692;
  wire [13:0] _GEN_1694 = 14'h69e == index ? 14'hd : _GEN_1693;
  wire [13:0] _GEN_1695 = 14'h69f == index ? 14'hd : _GEN_1694;
  wire [13:0] _GEN_1696 = 14'h6a0 == index ? 14'hd : _GEN_1695;
  wire [13:0] _GEN_1697 = 14'h6a1 == index ? 14'hd : _GEN_1696;
  wire [13:0] _GEN_1698 = 14'h6a2 == index ? 14'hd : _GEN_1697;
  wire [13:0] _GEN_1699 = 14'h6a3 == index ? 14'hd : _GEN_1698;
  wire [13:0] _GEN_1700 = 14'h6a4 == index ? 14'hd : _GEN_1699;
  wire [13:0] _GEN_1701 = 14'h6a5 == index ? 14'hd : _GEN_1700;
  wire [13:0] _GEN_1702 = 14'h6a6 == index ? 14'hd : _GEN_1701;
  wire [13:0] _GEN_1703 = 14'h6a7 == index ? 14'hd : _GEN_1702;
  wire [13:0] _GEN_1704 = 14'h6a8 == index ? 14'hd : _GEN_1703;
  wire [13:0] _GEN_1705 = 14'h6a9 == index ? 14'hd : _GEN_1704;
  wire [13:0] _GEN_1706 = 14'h6aa == index ? 14'hd : _GEN_1705;
  wire [13:0] _GEN_1707 = 14'h6ab == index ? 14'hd : _GEN_1706;
  wire [13:0] _GEN_1708 = 14'h6ac == index ? 14'hd : _GEN_1707;
  wire [13:0] _GEN_1709 = 14'h6ad == index ? 14'hd : _GEN_1708;
  wire [13:0] _GEN_1710 = 14'h6ae == index ? 14'hd : _GEN_1709;
  wire [13:0] _GEN_1711 = 14'h6af == index ? 14'hd : _GEN_1710;
  wire [13:0] _GEN_1712 = 14'h6b0 == index ? 14'hd : _GEN_1711;
  wire [13:0] _GEN_1713 = 14'h6b1 == index ? 14'hd : _GEN_1712;
  wire [13:0] _GEN_1714 = 14'h6b2 == index ? 14'hd : _GEN_1713;
  wire [13:0] _GEN_1715 = 14'h6b3 == index ? 14'hd : _GEN_1714;
  wire [13:0] _GEN_1716 = 14'h6b4 == index ? 14'hd : _GEN_1715;
  wire [13:0] _GEN_1717 = 14'h6b5 == index ? 14'hd : _GEN_1716;
  wire [13:0] _GEN_1718 = 14'h6b6 == index ? 14'hd : _GEN_1717;
  wire [13:0] _GEN_1719 = 14'h6b7 == index ? 14'hd : _GEN_1718;
  wire [13:0] _GEN_1720 = 14'h6b8 == index ? 14'hd : _GEN_1719;
  wire [13:0] _GEN_1721 = 14'h6b9 == index ? 14'hd : _GEN_1720;
  wire [13:0] _GEN_1722 = 14'h6ba == index ? 14'hd : _GEN_1721;
  wire [13:0] _GEN_1723 = 14'h6bb == index ? 14'hd : _GEN_1722;
  wire [13:0] _GEN_1724 = 14'h6bc == index ? 14'hd : _GEN_1723;
  wire [13:0] _GEN_1725 = 14'h6bd == index ? 14'hd : _GEN_1724;
  wire [13:0] _GEN_1726 = 14'h6be == index ? 14'hd : _GEN_1725;
  wire [13:0] _GEN_1727 = 14'h6bf == index ? 14'hd : _GEN_1726;
  wire [13:0] _GEN_1728 = 14'h6c0 == index ? 14'hd : _GEN_1727;
  wire [13:0] _GEN_1729 = 14'h6c1 == index ? 14'hd : _GEN_1728;
  wire [13:0] _GEN_1730 = 14'h6c2 == index ? 14'hd : _GEN_1729;
  wire [13:0] _GEN_1731 = 14'h6c3 == index ? 14'hd : _GEN_1730;
  wire [13:0] _GEN_1732 = 14'h6c4 == index ? 14'hd : _GEN_1731;
  wire [13:0] _GEN_1733 = 14'h6c5 == index ? 14'hd : _GEN_1732;
  wire [13:0] _GEN_1734 = 14'h6c6 == index ? 14'hd : _GEN_1733;
  wire [13:0] _GEN_1735 = 14'h6c7 == index ? 14'hd : _GEN_1734;
  wire [13:0] _GEN_1736 = 14'h6c8 == index ? 14'hd : _GEN_1735;
  wire [13:0] _GEN_1737 = 14'h6c9 == index ? 14'hd : _GEN_1736;
  wire [13:0] _GEN_1738 = 14'h6ca == index ? 14'hd : _GEN_1737;
  wire [13:0] _GEN_1739 = 14'h6cb == index ? 14'hd : _GEN_1738;
  wire [13:0] _GEN_1740 = 14'h6cc == index ? 14'hd : _GEN_1739;
  wire [13:0] _GEN_1741 = 14'h6cd == index ? 14'hd : _GEN_1740;
  wire [13:0] _GEN_1742 = 14'h6ce == index ? 14'hd : _GEN_1741;
  wire [13:0] _GEN_1743 = 14'h6cf == index ? 14'hd : _GEN_1742;
  wire [13:0] _GEN_1744 = 14'h6d0 == index ? 14'hd : _GEN_1743;
  wire [13:0] _GEN_1745 = 14'h6d1 == index ? 14'hd : _GEN_1744;
  wire [13:0] _GEN_1746 = 14'h6d2 == index ? 14'hd : _GEN_1745;
  wire [13:0] _GEN_1747 = 14'h6d3 == index ? 14'hd : _GEN_1746;
  wire [13:0] _GEN_1748 = 14'h6d4 == index ? 14'hd : _GEN_1747;
  wire [13:0] _GEN_1749 = 14'h6d5 == index ? 14'hd : _GEN_1748;
  wire [13:0] _GEN_1750 = 14'h6d6 == index ? 14'hd : _GEN_1749;
  wire [13:0] _GEN_1751 = 14'h6d7 == index ? 14'hd : _GEN_1750;
  wire [13:0] _GEN_1752 = 14'h6d8 == index ? 14'hd : _GEN_1751;
  wire [13:0] _GEN_1753 = 14'h6d9 == index ? 14'hd : _GEN_1752;
  wire [13:0] _GEN_1754 = 14'h6da == index ? 14'hd : _GEN_1753;
  wire [13:0] _GEN_1755 = 14'h6db == index ? 14'hd : _GEN_1754;
  wire [13:0] _GEN_1756 = 14'h6dc == index ? 14'hd : _GEN_1755;
  wire [13:0] _GEN_1757 = 14'h6dd == index ? 14'hd : _GEN_1756;
  wire [13:0] _GEN_1758 = 14'h6de == index ? 14'hd : _GEN_1757;
  wire [13:0] _GEN_1759 = 14'h6df == index ? 14'hd : _GEN_1758;
  wire [13:0] _GEN_1760 = 14'h6e0 == index ? 14'hd : _GEN_1759;
  wire [13:0] _GEN_1761 = 14'h6e1 == index ? 14'hd : _GEN_1760;
  wire [13:0] _GEN_1762 = 14'h6e2 == index ? 14'hd : _GEN_1761;
  wire [13:0] _GEN_1763 = 14'h6e3 == index ? 14'hd : _GEN_1762;
  wire [13:0] _GEN_1764 = 14'h6e4 == index ? 14'hd : _GEN_1763;
  wire [13:0] _GEN_1765 = 14'h6e5 == index ? 14'hd : _GEN_1764;
  wire [13:0] _GEN_1766 = 14'h6e6 == index ? 14'hd : _GEN_1765;
  wire [13:0] _GEN_1767 = 14'h6e7 == index ? 14'hd : _GEN_1766;
  wire [13:0] _GEN_1768 = 14'h6e8 == index ? 14'hd : _GEN_1767;
  wire [13:0] _GEN_1769 = 14'h6e9 == index ? 14'hd : _GEN_1768;
  wire [13:0] _GEN_1770 = 14'h6ea == index ? 14'hd : _GEN_1769;
  wire [13:0] _GEN_1771 = 14'h6eb == index ? 14'hd : _GEN_1770;
  wire [13:0] _GEN_1772 = 14'h6ec == index ? 14'hd : _GEN_1771;
  wire [13:0] _GEN_1773 = 14'h6ed == index ? 14'hd : _GEN_1772;
  wire [13:0] _GEN_1774 = 14'h6ee == index ? 14'hd : _GEN_1773;
  wire [13:0] _GEN_1775 = 14'h6ef == index ? 14'hd : _GEN_1774;
  wire [13:0] _GEN_1776 = 14'h6f0 == index ? 14'hd : _GEN_1775;
  wire [13:0] _GEN_1777 = 14'h6f1 == index ? 14'hd : _GEN_1776;
  wire [13:0] _GEN_1778 = 14'h6f2 == index ? 14'hd : _GEN_1777;
  wire [13:0] _GEN_1779 = 14'h6f3 == index ? 14'hd : _GEN_1778;
  wire [13:0] _GEN_1780 = 14'h6f4 == index ? 14'hd : _GEN_1779;
  wire [13:0] _GEN_1781 = 14'h6f5 == index ? 14'hd : _GEN_1780;
  wire [13:0] _GEN_1782 = 14'h6f6 == index ? 14'hd : _GEN_1781;
  wire [13:0] _GEN_1783 = 14'h6f7 == index ? 14'hd : _GEN_1782;
  wire [13:0] _GEN_1784 = 14'h6f8 == index ? 14'hd : _GEN_1783;
  wire [13:0] _GEN_1785 = 14'h6f9 == index ? 14'hd : _GEN_1784;
  wire [13:0] _GEN_1786 = 14'h6fa == index ? 14'hd : _GEN_1785;
  wire [13:0] _GEN_1787 = 14'h6fb == index ? 14'hd : _GEN_1786;
  wire [13:0] _GEN_1788 = 14'h6fc == index ? 14'hd : _GEN_1787;
  wire [13:0] _GEN_1789 = 14'h6fd == index ? 14'hd : _GEN_1788;
  wire [13:0] _GEN_1790 = 14'h6fe == index ? 14'hd : _GEN_1789;
  wire [13:0] _GEN_1791 = 14'h6ff == index ? 14'hd : _GEN_1790;
  wire [13:0] _GEN_1792 = 14'h700 == index ? 14'h0 : _GEN_1791;
  wire [13:0] _GEN_1793 = 14'h701 == index ? 14'h700 : _GEN_1792;
  wire [13:0] _GEN_1794 = 14'h702 == index ? 14'h380 : _GEN_1793;
  wire [13:0] _GEN_1795 = 14'h703 == index ? 14'h202 : _GEN_1794;
  wire [13:0] _GEN_1796 = 14'h704 == index ? 14'h182 : _GEN_1795;
  wire [13:0] _GEN_1797 = 14'h705 == index ? 14'h104 : _GEN_1796;
  wire [13:0] _GEN_1798 = 14'h706 == index ? 14'h102 : _GEN_1797;
  wire [13:0] _GEN_1799 = 14'h707 == index ? 14'h100 : _GEN_1798;
  wire [13:0] _GEN_1800 = 14'h708 == index ? 14'h86 : _GEN_1799;
  wire [13:0] _GEN_1801 = 14'h709 == index ? 14'h85 : _GEN_1800;
  wire [13:0] _GEN_1802 = 14'h70a == index ? 14'h84 : _GEN_1801;
  wire [13:0] _GEN_1803 = 14'h70b == index ? 14'h83 : _GEN_1802;
  wire [13:0] _GEN_1804 = 14'h70c == index ? 14'h82 : _GEN_1803;
  wire [13:0] _GEN_1805 = 14'h70d == index ? 14'h81 : _GEN_1804;
  wire [13:0] _GEN_1806 = 14'h70e == index ? 14'h80 : _GEN_1805;
  wire [13:0] _GEN_1807 = 14'h70f == index ? 14'he : _GEN_1806;
  wire [13:0] _GEN_1808 = 14'h710 == index ? 14'he : _GEN_1807;
  wire [13:0] _GEN_1809 = 14'h711 == index ? 14'he : _GEN_1808;
  wire [13:0] _GEN_1810 = 14'h712 == index ? 14'he : _GEN_1809;
  wire [13:0] _GEN_1811 = 14'h713 == index ? 14'he : _GEN_1810;
  wire [13:0] _GEN_1812 = 14'h714 == index ? 14'he : _GEN_1811;
  wire [13:0] _GEN_1813 = 14'h715 == index ? 14'he : _GEN_1812;
  wire [13:0] _GEN_1814 = 14'h716 == index ? 14'he : _GEN_1813;
  wire [13:0] _GEN_1815 = 14'h717 == index ? 14'he : _GEN_1814;
  wire [13:0] _GEN_1816 = 14'h718 == index ? 14'he : _GEN_1815;
  wire [13:0] _GEN_1817 = 14'h719 == index ? 14'he : _GEN_1816;
  wire [13:0] _GEN_1818 = 14'h71a == index ? 14'he : _GEN_1817;
  wire [13:0] _GEN_1819 = 14'h71b == index ? 14'he : _GEN_1818;
  wire [13:0] _GEN_1820 = 14'h71c == index ? 14'he : _GEN_1819;
  wire [13:0] _GEN_1821 = 14'h71d == index ? 14'he : _GEN_1820;
  wire [13:0] _GEN_1822 = 14'h71e == index ? 14'he : _GEN_1821;
  wire [13:0] _GEN_1823 = 14'h71f == index ? 14'he : _GEN_1822;
  wire [13:0] _GEN_1824 = 14'h720 == index ? 14'he : _GEN_1823;
  wire [13:0] _GEN_1825 = 14'h721 == index ? 14'he : _GEN_1824;
  wire [13:0] _GEN_1826 = 14'h722 == index ? 14'he : _GEN_1825;
  wire [13:0] _GEN_1827 = 14'h723 == index ? 14'he : _GEN_1826;
  wire [13:0] _GEN_1828 = 14'h724 == index ? 14'he : _GEN_1827;
  wire [13:0] _GEN_1829 = 14'h725 == index ? 14'he : _GEN_1828;
  wire [13:0] _GEN_1830 = 14'h726 == index ? 14'he : _GEN_1829;
  wire [13:0] _GEN_1831 = 14'h727 == index ? 14'he : _GEN_1830;
  wire [13:0] _GEN_1832 = 14'h728 == index ? 14'he : _GEN_1831;
  wire [13:0] _GEN_1833 = 14'h729 == index ? 14'he : _GEN_1832;
  wire [13:0] _GEN_1834 = 14'h72a == index ? 14'he : _GEN_1833;
  wire [13:0] _GEN_1835 = 14'h72b == index ? 14'he : _GEN_1834;
  wire [13:0] _GEN_1836 = 14'h72c == index ? 14'he : _GEN_1835;
  wire [13:0] _GEN_1837 = 14'h72d == index ? 14'he : _GEN_1836;
  wire [13:0] _GEN_1838 = 14'h72e == index ? 14'he : _GEN_1837;
  wire [13:0] _GEN_1839 = 14'h72f == index ? 14'he : _GEN_1838;
  wire [13:0] _GEN_1840 = 14'h730 == index ? 14'he : _GEN_1839;
  wire [13:0] _GEN_1841 = 14'h731 == index ? 14'he : _GEN_1840;
  wire [13:0] _GEN_1842 = 14'h732 == index ? 14'he : _GEN_1841;
  wire [13:0] _GEN_1843 = 14'h733 == index ? 14'he : _GEN_1842;
  wire [13:0] _GEN_1844 = 14'h734 == index ? 14'he : _GEN_1843;
  wire [13:0] _GEN_1845 = 14'h735 == index ? 14'he : _GEN_1844;
  wire [13:0] _GEN_1846 = 14'h736 == index ? 14'he : _GEN_1845;
  wire [13:0] _GEN_1847 = 14'h737 == index ? 14'he : _GEN_1846;
  wire [13:0] _GEN_1848 = 14'h738 == index ? 14'he : _GEN_1847;
  wire [13:0] _GEN_1849 = 14'h739 == index ? 14'he : _GEN_1848;
  wire [13:0] _GEN_1850 = 14'h73a == index ? 14'he : _GEN_1849;
  wire [13:0] _GEN_1851 = 14'h73b == index ? 14'he : _GEN_1850;
  wire [13:0] _GEN_1852 = 14'h73c == index ? 14'he : _GEN_1851;
  wire [13:0] _GEN_1853 = 14'h73d == index ? 14'he : _GEN_1852;
  wire [13:0] _GEN_1854 = 14'h73e == index ? 14'he : _GEN_1853;
  wire [13:0] _GEN_1855 = 14'h73f == index ? 14'he : _GEN_1854;
  wire [13:0] _GEN_1856 = 14'h740 == index ? 14'he : _GEN_1855;
  wire [13:0] _GEN_1857 = 14'h741 == index ? 14'he : _GEN_1856;
  wire [13:0] _GEN_1858 = 14'h742 == index ? 14'he : _GEN_1857;
  wire [13:0] _GEN_1859 = 14'h743 == index ? 14'he : _GEN_1858;
  wire [13:0] _GEN_1860 = 14'h744 == index ? 14'he : _GEN_1859;
  wire [13:0] _GEN_1861 = 14'h745 == index ? 14'he : _GEN_1860;
  wire [13:0] _GEN_1862 = 14'h746 == index ? 14'he : _GEN_1861;
  wire [13:0] _GEN_1863 = 14'h747 == index ? 14'he : _GEN_1862;
  wire [13:0] _GEN_1864 = 14'h748 == index ? 14'he : _GEN_1863;
  wire [13:0] _GEN_1865 = 14'h749 == index ? 14'he : _GEN_1864;
  wire [13:0] _GEN_1866 = 14'h74a == index ? 14'he : _GEN_1865;
  wire [13:0] _GEN_1867 = 14'h74b == index ? 14'he : _GEN_1866;
  wire [13:0] _GEN_1868 = 14'h74c == index ? 14'he : _GEN_1867;
  wire [13:0] _GEN_1869 = 14'h74d == index ? 14'he : _GEN_1868;
  wire [13:0] _GEN_1870 = 14'h74e == index ? 14'he : _GEN_1869;
  wire [13:0] _GEN_1871 = 14'h74f == index ? 14'he : _GEN_1870;
  wire [13:0] _GEN_1872 = 14'h750 == index ? 14'he : _GEN_1871;
  wire [13:0] _GEN_1873 = 14'h751 == index ? 14'he : _GEN_1872;
  wire [13:0] _GEN_1874 = 14'h752 == index ? 14'he : _GEN_1873;
  wire [13:0] _GEN_1875 = 14'h753 == index ? 14'he : _GEN_1874;
  wire [13:0] _GEN_1876 = 14'h754 == index ? 14'he : _GEN_1875;
  wire [13:0] _GEN_1877 = 14'h755 == index ? 14'he : _GEN_1876;
  wire [13:0] _GEN_1878 = 14'h756 == index ? 14'he : _GEN_1877;
  wire [13:0] _GEN_1879 = 14'h757 == index ? 14'he : _GEN_1878;
  wire [13:0] _GEN_1880 = 14'h758 == index ? 14'he : _GEN_1879;
  wire [13:0] _GEN_1881 = 14'h759 == index ? 14'he : _GEN_1880;
  wire [13:0] _GEN_1882 = 14'h75a == index ? 14'he : _GEN_1881;
  wire [13:0] _GEN_1883 = 14'h75b == index ? 14'he : _GEN_1882;
  wire [13:0] _GEN_1884 = 14'h75c == index ? 14'he : _GEN_1883;
  wire [13:0] _GEN_1885 = 14'h75d == index ? 14'he : _GEN_1884;
  wire [13:0] _GEN_1886 = 14'h75e == index ? 14'he : _GEN_1885;
  wire [13:0] _GEN_1887 = 14'h75f == index ? 14'he : _GEN_1886;
  wire [13:0] _GEN_1888 = 14'h760 == index ? 14'he : _GEN_1887;
  wire [13:0] _GEN_1889 = 14'h761 == index ? 14'he : _GEN_1888;
  wire [13:0] _GEN_1890 = 14'h762 == index ? 14'he : _GEN_1889;
  wire [13:0] _GEN_1891 = 14'h763 == index ? 14'he : _GEN_1890;
  wire [13:0] _GEN_1892 = 14'h764 == index ? 14'he : _GEN_1891;
  wire [13:0] _GEN_1893 = 14'h765 == index ? 14'he : _GEN_1892;
  wire [13:0] _GEN_1894 = 14'h766 == index ? 14'he : _GEN_1893;
  wire [13:0] _GEN_1895 = 14'h767 == index ? 14'he : _GEN_1894;
  wire [13:0] _GEN_1896 = 14'h768 == index ? 14'he : _GEN_1895;
  wire [13:0] _GEN_1897 = 14'h769 == index ? 14'he : _GEN_1896;
  wire [13:0] _GEN_1898 = 14'h76a == index ? 14'he : _GEN_1897;
  wire [13:0] _GEN_1899 = 14'h76b == index ? 14'he : _GEN_1898;
  wire [13:0] _GEN_1900 = 14'h76c == index ? 14'he : _GEN_1899;
  wire [13:0] _GEN_1901 = 14'h76d == index ? 14'he : _GEN_1900;
  wire [13:0] _GEN_1902 = 14'h76e == index ? 14'he : _GEN_1901;
  wire [13:0] _GEN_1903 = 14'h76f == index ? 14'he : _GEN_1902;
  wire [13:0] _GEN_1904 = 14'h770 == index ? 14'he : _GEN_1903;
  wire [13:0] _GEN_1905 = 14'h771 == index ? 14'he : _GEN_1904;
  wire [13:0] _GEN_1906 = 14'h772 == index ? 14'he : _GEN_1905;
  wire [13:0] _GEN_1907 = 14'h773 == index ? 14'he : _GEN_1906;
  wire [13:0] _GEN_1908 = 14'h774 == index ? 14'he : _GEN_1907;
  wire [13:0] _GEN_1909 = 14'h775 == index ? 14'he : _GEN_1908;
  wire [13:0] _GEN_1910 = 14'h776 == index ? 14'he : _GEN_1909;
  wire [13:0] _GEN_1911 = 14'h777 == index ? 14'he : _GEN_1910;
  wire [13:0] _GEN_1912 = 14'h778 == index ? 14'he : _GEN_1911;
  wire [13:0] _GEN_1913 = 14'h779 == index ? 14'he : _GEN_1912;
  wire [13:0] _GEN_1914 = 14'h77a == index ? 14'he : _GEN_1913;
  wire [13:0] _GEN_1915 = 14'h77b == index ? 14'he : _GEN_1914;
  wire [13:0] _GEN_1916 = 14'h77c == index ? 14'he : _GEN_1915;
  wire [13:0] _GEN_1917 = 14'h77d == index ? 14'he : _GEN_1916;
  wire [13:0] _GEN_1918 = 14'h77e == index ? 14'he : _GEN_1917;
  wire [13:0] _GEN_1919 = 14'h77f == index ? 14'he : _GEN_1918;
  wire [13:0] _GEN_1920 = 14'h780 == index ? 14'h0 : _GEN_1919;
  wire [13:0] _GEN_1921 = 14'h781 == index ? 14'h780 : _GEN_1920;
  wire [13:0] _GEN_1922 = 14'h782 == index ? 14'h381 : _GEN_1921;
  wire [13:0] _GEN_1923 = 14'h783 == index ? 14'h280 : _GEN_1922;
  wire [13:0] _GEN_1924 = 14'h784 == index ? 14'h183 : _GEN_1923;
  wire [13:0] _GEN_1925 = 14'h785 == index ? 14'h180 : _GEN_1924;
  wire [13:0] _GEN_1926 = 14'h786 == index ? 14'h103 : _GEN_1925;
  wire [13:0] _GEN_1927 = 14'h787 == index ? 14'h101 : _GEN_1926;
  wire [13:0] _GEN_1928 = 14'h788 == index ? 14'h87 : _GEN_1927;
  wire [13:0] _GEN_1929 = 14'h789 == index ? 14'h86 : _GEN_1928;
  wire [13:0] _GEN_1930 = 14'h78a == index ? 14'h85 : _GEN_1929;
  wire [13:0] _GEN_1931 = 14'h78b == index ? 14'h84 : _GEN_1930;
  wire [13:0] _GEN_1932 = 14'h78c == index ? 14'h83 : _GEN_1931;
  wire [13:0] _GEN_1933 = 14'h78d == index ? 14'h82 : _GEN_1932;
  wire [13:0] _GEN_1934 = 14'h78e == index ? 14'h81 : _GEN_1933;
  wire [13:0] _GEN_1935 = 14'h78f == index ? 14'h80 : _GEN_1934;
  wire [13:0] _GEN_1936 = 14'h790 == index ? 14'hf : _GEN_1935;
  wire [13:0] _GEN_1937 = 14'h791 == index ? 14'hf : _GEN_1936;
  wire [13:0] _GEN_1938 = 14'h792 == index ? 14'hf : _GEN_1937;
  wire [13:0] _GEN_1939 = 14'h793 == index ? 14'hf : _GEN_1938;
  wire [13:0] _GEN_1940 = 14'h794 == index ? 14'hf : _GEN_1939;
  wire [13:0] _GEN_1941 = 14'h795 == index ? 14'hf : _GEN_1940;
  wire [13:0] _GEN_1942 = 14'h796 == index ? 14'hf : _GEN_1941;
  wire [13:0] _GEN_1943 = 14'h797 == index ? 14'hf : _GEN_1942;
  wire [13:0] _GEN_1944 = 14'h798 == index ? 14'hf : _GEN_1943;
  wire [13:0] _GEN_1945 = 14'h799 == index ? 14'hf : _GEN_1944;
  wire [13:0] _GEN_1946 = 14'h79a == index ? 14'hf : _GEN_1945;
  wire [13:0] _GEN_1947 = 14'h79b == index ? 14'hf : _GEN_1946;
  wire [13:0] _GEN_1948 = 14'h79c == index ? 14'hf : _GEN_1947;
  wire [13:0] _GEN_1949 = 14'h79d == index ? 14'hf : _GEN_1948;
  wire [13:0] _GEN_1950 = 14'h79e == index ? 14'hf : _GEN_1949;
  wire [13:0] _GEN_1951 = 14'h79f == index ? 14'hf : _GEN_1950;
  wire [13:0] _GEN_1952 = 14'h7a0 == index ? 14'hf : _GEN_1951;
  wire [13:0] _GEN_1953 = 14'h7a1 == index ? 14'hf : _GEN_1952;
  wire [13:0] _GEN_1954 = 14'h7a2 == index ? 14'hf : _GEN_1953;
  wire [13:0] _GEN_1955 = 14'h7a3 == index ? 14'hf : _GEN_1954;
  wire [13:0] _GEN_1956 = 14'h7a4 == index ? 14'hf : _GEN_1955;
  wire [13:0] _GEN_1957 = 14'h7a5 == index ? 14'hf : _GEN_1956;
  wire [13:0] _GEN_1958 = 14'h7a6 == index ? 14'hf : _GEN_1957;
  wire [13:0] _GEN_1959 = 14'h7a7 == index ? 14'hf : _GEN_1958;
  wire [13:0] _GEN_1960 = 14'h7a8 == index ? 14'hf : _GEN_1959;
  wire [13:0] _GEN_1961 = 14'h7a9 == index ? 14'hf : _GEN_1960;
  wire [13:0] _GEN_1962 = 14'h7aa == index ? 14'hf : _GEN_1961;
  wire [13:0] _GEN_1963 = 14'h7ab == index ? 14'hf : _GEN_1962;
  wire [13:0] _GEN_1964 = 14'h7ac == index ? 14'hf : _GEN_1963;
  wire [13:0] _GEN_1965 = 14'h7ad == index ? 14'hf : _GEN_1964;
  wire [13:0] _GEN_1966 = 14'h7ae == index ? 14'hf : _GEN_1965;
  wire [13:0] _GEN_1967 = 14'h7af == index ? 14'hf : _GEN_1966;
  wire [13:0] _GEN_1968 = 14'h7b0 == index ? 14'hf : _GEN_1967;
  wire [13:0] _GEN_1969 = 14'h7b1 == index ? 14'hf : _GEN_1968;
  wire [13:0] _GEN_1970 = 14'h7b2 == index ? 14'hf : _GEN_1969;
  wire [13:0] _GEN_1971 = 14'h7b3 == index ? 14'hf : _GEN_1970;
  wire [13:0] _GEN_1972 = 14'h7b4 == index ? 14'hf : _GEN_1971;
  wire [13:0] _GEN_1973 = 14'h7b5 == index ? 14'hf : _GEN_1972;
  wire [13:0] _GEN_1974 = 14'h7b6 == index ? 14'hf : _GEN_1973;
  wire [13:0] _GEN_1975 = 14'h7b7 == index ? 14'hf : _GEN_1974;
  wire [13:0] _GEN_1976 = 14'h7b8 == index ? 14'hf : _GEN_1975;
  wire [13:0] _GEN_1977 = 14'h7b9 == index ? 14'hf : _GEN_1976;
  wire [13:0] _GEN_1978 = 14'h7ba == index ? 14'hf : _GEN_1977;
  wire [13:0] _GEN_1979 = 14'h7bb == index ? 14'hf : _GEN_1978;
  wire [13:0] _GEN_1980 = 14'h7bc == index ? 14'hf : _GEN_1979;
  wire [13:0] _GEN_1981 = 14'h7bd == index ? 14'hf : _GEN_1980;
  wire [13:0] _GEN_1982 = 14'h7be == index ? 14'hf : _GEN_1981;
  wire [13:0] _GEN_1983 = 14'h7bf == index ? 14'hf : _GEN_1982;
  wire [13:0] _GEN_1984 = 14'h7c0 == index ? 14'hf : _GEN_1983;
  wire [13:0] _GEN_1985 = 14'h7c1 == index ? 14'hf : _GEN_1984;
  wire [13:0] _GEN_1986 = 14'h7c2 == index ? 14'hf : _GEN_1985;
  wire [13:0] _GEN_1987 = 14'h7c3 == index ? 14'hf : _GEN_1986;
  wire [13:0] _GEN_1988 = 14'h7c4 == index ? 14'hf : _GEN_1987;
  wire [13:0] _GEN_1989 = 14'h7c5 == index ? 14'hf : _GEN_1988;
  wire [13:0] _GEN_1990 = 14'h7c6 == index ? 14'hf : _GEN_1989;
  wire [13:0] _GEN_1991 = 14'h7c7 == index ? 14'hf : _GEN_1990;
  wire [13:0] _GEN_1992 = 14'h7c8 == index ? 14'hf : _GEN_1991;
  wire [13:0] _GEN_1993 = 14'h7c9 == index ? 14'hf : _GEN_1992;
  wire [13:0] _GEN_1994 = 14'h7ca == index ? 14'hf : _GEN_1993;
  wire [13:0] _GEN_1995 = 14'h7cb == index ? 14'hf : _GEN_1994;
  wire [13:0] _GEN_1996 = 14'h7cc == index ? 14'hf : _GEN_1995;
  wire [13:0] _GEN_1997 = 14'h7cd == index ? 14'hf : _GEN_1996;
  wire [13:0] _GEN_1998 = 14'h7ce == index ? 14'hf : _GEN_1997;
  wire [13:0] _GEN_1999 = 14'h7cf == index ? 14'hf : _GEN_1998;
  wire [13:0] _GEN_2000 = 14'h7d0 == index ? 14'hf : _GEN_1999;
  wire [13:0] _GEN_2001 = 14'h7d1 == index ? 14'hf : _GEN_2000;
  wire [13:0] _GEN_2002 = 14'h7d2 == index ? 14'hf : _GEN_2001;
  wire [13:0] _GEN_2003 = 14'h7d3 == index ? 14'hf : _GEN_2002;
  wire [13:0] _GEN_2004 = 14'h7d4 == index ? 14'hf : _GEN_2003;
  wire [13:0] _GEN_2005 = 14'h7d5 == index ? 14'hf : _GEN_2004;
  wire [13:0] _GEN_2006 = 14'h7d6 == index ? 14'hf : _GEN_2005;
  wire [13:0] _GEN_2007 = 14'h7d7 == index ? 14'hf : _GEN_2006;
  wire [13:0] _GEN_2008 = 14'h7d8 == index ? 14'hf : _GEN_2007;
  wire [13:0] _GEN_2009 = 14'h7d9 == index ? 14'hf : _GEN_2008;
  wire [13:0] _GEN_2010 = 14'h7da == index ? 14'hf : _GEN_2009;
  wire [13:0] _GEN_2011 = 14'h7db == index ? 14'hf : _GEN_2010;
  wire [13:0] _GEN_2012 = 14'h7dc == index ? 14'hf : _GEN_2011;
  wire [13:0] _GEN_2013 = 14'h7dd == index ? 14'hf : _GEN_2012;
  wire [13:0] _GEN_2014 = 14'h7de == index ? 14'hf : _GEN_2013;
  wire [13:0] _GEN_2015 = 14'h7df == index ? 14'hf : _GEN_2014;
  wire [13:0] _GEN_2016 = 14'h7e0 == index ? 14'hf : _GEN_2015;
  wire [13:0] _GEN_2017 = 14'h7e1 == index ? 14'hf : _GEN_2016;
  wire [13:0] _GEN_2018 = 14'h7e2 == index ? 14'hf : _GEN_2017;
  wire [13:0] _GEN_2019 = 14'h7e3 == index ? 14'hf : _GEN_2018;
  wire [13:0] _GEN_2020 = 14'h7e4 == index ? 14'hf : _GEN_2019;
  wire [13:0] _GEN_2021 = 14'h7e5 == index ? 14'hf : _GEN_2020;
  wire [13:0] _GEN_2022 = 14'h7e6 == index ? 14'hf : _GEN_2021;
  wire [13:0] _GEN_2023 = 14'h7e7 == index ? 14'hf : _GEN_2022;
  wire [13:0] _GEN_2024 = 14'h7e8 == index ? 14'hf : _GEN_2023;
  wire [13:0] _GEN_2025 = 14'h7e9 == index ? 14'hf : _GEN_2024;
  wire [13:0] _GEN_2026 = 14'h7ea == index ? 14'hf : _GEN_2025;
  wire [13:0] _GEN_2027 = 14'h7eb == index ? 14'hf : _GEN_2026;
  wire [13:0] _GEN_2028 = 14'h7ec == index ? 14'hf : _GEN_2027;
  wire [13:0] _GEN_2029 = 14'h7ed == index ? 14'hf : _GEN_2028;
  wire [13:0] _GEN_2030 = 14'h7ee == index ? 14'hf : _GEN_2029;
  wire [13:0] _GEN_2031 = 14'h7ef == index ? 14'hf : _GEN_2030;
  wire [13:0] _GEN_2032 = 14'h7f0 == index ? 14'hf : _GEN_2031;
  wire [13:0] _GEN_2033 = 14'h7f1 == index ? 14'hf : _GEN_2032;
  wire [13:0] _GEN_2034 = 14'h7f2 == index ? 14'hf : _GEN_2033;
  wire [13:0] _GEN_2035 = 14'h7f3 == index ? 14'hf : _GEN_2034;
  wire [13:0] _GEN_2036 = 14'h7f4 == index ? 14'hf : _GEN_2035;
  wire [13:0] _GEN_2037 = 14'h7f5 == index ? 14'hf : _GEN_2036;
  wire [13:0] _GEN_2038 = 14'h7f6 == index ? 14'hf : _GEN_2037;
  wire [13:0] _GEN_2039 = 14'h7f7 == index ? 14'hf : _GEN_2038;
  wire [13:0] _GEN_2040 = 14'h7f8 == index ? 14'hf : _GEN_2039;
  wire [13:0] _GEN_2041 = 14'h7f9 == index ? 14'hf : _GEN_2040;
  wire [13:0] _GEN_2042 = 14'h7fa == index ? 14'hf : _GEN_2041;
  wire [13:0] _GEN_2043 = 14'h7fb == index ? 14'hf : _GEN_2042;
  wire [13:0] _GEN_2044 = 14'h7fc == index ? 14'hf : _GEN_2043;
  wire [13:0] _GEN_2045 = 14'h7fd == index ? 14'hf : _GEN_2044;
  wire [13:0] _GEN_2046 = 14'h7fe == index ? 14'hf : _GEN_2045;
  wire [13:0] _GEN_2047 = 14'h7ff == index ? 14'hf : _GEN_2046;
  wire [13:0] _GEN_2048 = 14'h800 == index ? 14'h0 : _GEN_2047;
  wire [13:0] _GEN_2049 = 14'h801 == index ? 14'h800 : _GEN_2048;
  wire [13:0] _GEN_2050 = 14'h802 == index ? 14'h400 : _GEN_2049;
  wire [13:0] _GEN_2051 = 14'h803 == index ? 14'h281 : _GEN_2050;
  wire [13:0] _GEN_2052 = 14'h804 == index ? 14'h200 : _GEN_2051;
  wire [13:0] _GEN_2053 = 14'h805 == index ? 14'h181 : _GEN_2052;
  wire [13:0] _GEN_2054 = 14'h806 == index ? 14'h104 : _GEN_2053;
  wire [13:0] _GEN_2055 = 14'h807 == index ? 14'h102 : _GEN_2054;
  wire [13:0] _GEN_2056 = 14'h808 == index ? 14'h100 : _GEN_2055;
  wire [13:0] _GEN_2057 = 14'h809 == index ? 14'h87 : _GEN_2056;
  wire [13:0] _GEN_2058 = 14'h80a == index ? 14'h86 : _GEN_2057;
  wire [13:0] _GEN_2059 = 14'h80b == index ? 14'h85 : _GEN_2058;
  wire [13:0] _GEN_2060 = 14'h80c == index ? 14'h84 : _GEN_2059;
  wire [13:0] _GEN_2061 = 14'h80d == index ? 14'h83 : _GEN_2060;
  wire [13:0] _GEN_2062 = 14'h80e == index ? 14'h82 : _GEN_2061;
  wire [13:0] _GEN_2063 = 14'h80f == index ? 14'h81 : _GEN_2062;
  wire [13:0] _GEN_2064 = 14'h810 == index ? 14'h80 : _GEN_2063;
  wire [13:0] _GEN_2065 = 14'h811 == index ? 14'h10 : _GEN_2064;
  wire [13:0] _GEN_2066 = 14'h812 == index ? 14'h10 : _GEN_2065;
  wire [13:0] _GEN_2067 = 14'h813 == index ? 14'h10 : _GEN_2066;
  wire [13:0] _GEN_2068 = 14'h814 == index ? 14'h10 : _GEN_2067;
  wire [13:0] _GEN_2069 = 14'h815 == index ? 14'h10 : _GEN_2068;
  wire [13:0] _GEN_2070 = 14'h816 == index ? 14'h10 : _GEN_2069;
  wire [13:0] _GEN_2071 = 14'h817 == index ? 14'h10 : _GEN_2070;
  wire [13:0] _GEN_2072 = 14'h818 == index ? 14'h10 : _GEN_2071;
  wire [13:0] _GEN_2073 = 14'h819 == index ? 14'h10 : _GEN_2072;
  wire [13:0] _GEN_2074 = 14'h81a == index ? 14'h10 : _GEN_2073;
  wire [13:0] _GEN_2075 = 14'h81b == index ? 14'h10 : _GEN_2074;
  wire [13:0] _GEN_2076 = 14'h81c == index ? 14'h10 : _GEN_2075;
  wire [13:0] _GEN_2077 = 14'h81d == index ? 14'h10 : _GEN_2076;
  wire [13:0] _GEN_2078 = 14'h81e == index ? 14'h10 : _GEN_2077;
  wire [13:0] _GEN_2079 = 14'h81f == index ? 14'h10 : _GEN_2078;
  wire [13:0] _GEN_2080 = 14'h820 == index ? 14'h10 : _GEN_2079;
  wire [13:0] _GEN_2081 = 14'h821 == index ? 14'h10 : _GEN_2080;
  wire [13:0] _GEN_2082 = 14'h822 == index ? 14'h10 : _GEN_2081;
  wire [13:0] _GEN_2083 = 14'h823 == index ? 14'h10 : _GEN_2082;
  wire [13:0] _GEN_2084 = 14'h824 == index ? 14'h10 : _GEN_2083;
  wire [13:0] _GEN_2085 = 14'h825 == index ? 14'h10 : _GEN_2084;
  wire [13:0] _GEN_2086 = 14'h826 == index ? 14'h10 : _GEN_2085;
  wire [13:0] _GEN_2087 = 14'h827 == index ? 14'h10 : _GEN_2086;
  wire [13:0] _GEN_2088 = 14'h828 == index ? 14'h10 : _GEN_2087;
  wire [13:0] _GEN_2089 = 14'h829 == index ? 14'h10 : _GEN_2088;
  wire [13:0] _GEN_2090 = 14'h82a == index ? 14'h10 : _GEN_2089;
  wire [13:0] _GEN_2091 = 14'h82b == index ? 14'h10 : _GEN_2090;
  wire [13:0] _GEN_2092 = 14'h82c == index ? 14'h10 : _GEN_2091;
  wire [13:0] _GEN_2093 = 14'h82d == index ? 14'h10 : _GEN_2092;
  wire [13:0] _GEN_2094 = 14'h82e == index ? 14'h10 : _GEN_2093;
  wire [13:0] _GEN_2095 = 14'h82f == index ? 14'h10 : _GEN_2094;
  wire [13:0] _GEN_2096 = 14'h830 == index ? 14'h10 : _GEN_2095;
  wire [13:0] _GEN_2097 = 14'h831 == index ? 14'h10 : _GEN_2096;
  wire [13:0] _GEN_2098 = 14'h832 == index ? 14'h10 : _GEN_2097;
  wire [13:0] _GEN_2099 = 14'h833 == index ? 14'h10 : _GEN_2098;
  wire [13:0] _GEN_2100 = 14'h834 == index ? 14'h10 : _GEN_2099;
  wire [13:0] _GEN_2101 = 14'h835 == index ? 14'h10 : _GEN_2100;
  wire [13:0] _GEN_2102 = 14'h836 == index ? 14'h10 : _GEN_2101;
  wire [13:0] _GEN_2103 = 14'h837 == index ? 14'h10 : _GEN_2102;
  wire [13:0] _GEN_2104 = 14'h838 == index ? 14'h10 : _GEN_2103;
  wire [13:0] _GEN_2105 = 14'h839 == index ? 14'h10 : _GEN_2104;
  wire [13:0] _GEN_2106 = 14'h83a == index ? 14'h10 : _GEN_2105;
  wire [13:0] _GEN_2107 = 14'h83b == index ? 14'h10 : _GEN_2106;
  wire [13:0] _GEN_2108 = 14'h83c == index ? 14'h10 : _GEN_2107;
  wire [13:0] _GEN_2109 = 14'h83d == index ? 14'h10 : _GEN_2108;
  wire [13:0] _GEN_2110 = 14'h83e == index ? 14'h10 : _GEN_2109;
  wire [13:0] _GEN_2111 = 14'h83f == index ? 14'h10 : _GEN_2110;
  wire [13:0] _GEN_2112 = 14'h840 == index ? 14'h10 : _GEN_2111;
  wire [13:0] _GEN_2113 = 14'h841 == index ? 14'h10 : _GEN_2112;
  wire [13:0] _GEN_2114 = 14'h842 == index ? 14'h10 : _GEN_2113;
  wire [13:0] _GEN_2115 = 14'h843 == index ? 14'h10 : _GEN_2114;
  wire [13:0] _GEN_2116 = 14'h844 == index ? 14'h10 : _GEN_2115;
  wire [13:0] _GEN_2117 = 14'h845 == index ? 14'h10 : _GEN_2116;
  wire [13:0] _GEN_2118 = 14'h846 == index ? 14'h10 : _GEN_2117;
  wire [13:0] _GEN_2119 = 14'h847 == index ? 14'h10 : _GEN_2118;
  wire [13:0] _GEN_2120 = 14'h848 == index ? 14'h10 : _GEN_2119;
  wire [13:0] _GEN_2121 = 14'h849 == index ? 14'h10 : _GEN_2120;
  wire [13:0] _GEN_2122 = 14'h84a == index ? 14'h10 : _GEN_2121;
  wire [13:0] _GEN_2123 = 14'h84b == index ? 14'h10 : _GEN_2122;
  wire [13:0] _GEN_2124 = 14'h84c == index ? 14'h10 : _GEN_2123;
  wire [13:0] _GEN_2125 = 14'h84d == index ? 14'h10 : _GEN_2124;
  wire [13:0] _GEN_2126 = 14'h84e == index ? 14'h10 : _GEN_2125;
  wire [13:0] _GEN_2127 = 14'h84f == index ? 14'h10 : _GEN_2126;
  wire [13:0] _GEN_2128 = 14'h850 == index ? 14'h10 : _GEN_2127;
  wire [13:0] _GEN_2129 = 14'h851 == index ? 14'h10 : _GEN_2128;
  wire [13:0] _GEN_2130 = 14'h852 == index ? 14'h10 : _GEN_2129;
  wire [13:0] _GEN_2131 = 14'h853 == index ? 14'h10 : _GEN_2130;
  wire [13:0] _GEN_2132 = 14'h854 == index ? 14'h10 : _GEN_2131;
  wire [13:0] _GEN_2133 = 14'h855 == index ? 14'h10 : _GEN_2132;
  wire [13:0] _GEN_2134 = 14'h856 == index ? 14'h10 : _GEN_2133;
  wire [13:0] _GEN_2135 = 14'h857 == index ? 14'h10 : _GEN_2134;
  wire [13:0] _GEN_2136 = 14'h858 == index ? 14'h10 : _GEN_2135;
  wire [13:0] _GEN_2137 = 14'h859 == index ? 14'h10 : _GEN_2136;
  wire [13:0] _GEN_2138 = 14'h85a == index ? 14'h10 : _GEN_2137;
  wire [13:0] _GEN_2139 = 14'h85b == index ? 14'h10 : _GEN_2138;
  wire [13:0] _GEN_2140 = 14'h85c == index ? 14'h10 : _GEN_2139;
  wire [13:0] _GEN_2141 = 14'h85d == index ? 14'h10 : _GEN_2140;
  wire [13:0] _GEN_2142 = 14'h85e == index ? 14'h10 : _GEN_2141;
  wire [13:0] _GEN_2143 = 14'h85f == index ? 14'h10 : _GEN_2142;
  wire [13:0] _GEN_2144 = 14'h860 == index ? 14'h10 : _GEN_2143;
  wire [13:0] _GEN_2145 = 14'h861 == index ? 14'h10 : _GEN_2144;
  wire [13:0] _GEN_2146 = 14'h862 == index ? 14'h10 : _GEN_2145;
  wire [13:0] _GEN_2147 = 14'h863 == index ? 14'h10 : _GEN_2146;
  wire [13:0] _GEN_2148 = 14'h864 == index ? 14'h10 : _GEN_2147;
  wire [13:0] _GEN_2149 = 14'h865 == index ? 14'h10 : _GEN_2148;
  wire [13:0] _GEN_2150 = 14'h866 == index ? 14'h10 : _GEN_2149;
  wire [13:0] _GEN_2151 = 14'h867 == index ? 14'h10 : _GEN_2150;
  wire [13:0] _GEN_2152 = 14'h868 == index ? 14'h10 : _GEN_2151;
  wire [13:0] _GEN_2153 = 14'h869 == index ? 14'h10 : _GEN_2152;
  wire [13:0] _GEN_2154 = 14'h86a == index ? 14'h10 : _GEN_2153;
  wire [13:0] _GEN_2155 = 14'h86b == index ? 14'h10 : _GEN_2154;
  wire [13:0] _GEN_2156 = 14'h86c == index ? 14'h10 : _GEN_2155;
  wire [13:0] _GEN_2157 = 14'h86d == index ? 14'h10 : _GEN_2156;
  wire [13:0] _GEN_2158 = 14'h86e == index ? 14'h10 : _GEN_2157;
  wire [13:0] _GEN_2159 = 14'h86f == index ? 14'h10 : _GEN_2158;
  wire [13:0] _GEN_2160 = 14'h870 == index ? 14'h10 : _GEN_2159;
  wire [13:0] _GEN_2161 = 14'h871 == index ? 14'h10 : _GEN_2160;
  wire [13:0] _GEN_2162 = 14'h872 == index ? 14'h10 : _GEN_2161;
  wire [13:0] _GEN_2163 = 14'h873 == index ? 14'h10 : _GEN_2162;
  wire [13:0] _GEN_2164 = 14'h874 == index ? 14'h10 : _GEN_2163;
  wire [13:0] _GEN_2165 = 14'h875 == index ? 14'h10 : _GEN_2164;
  wire [13:0] _GEN_2166 = 14'h876 == index ? 14'h10 : _GEN_2165;
  wire [13:0] _GEN_2167 = 14'h877 == index ? 14'h10 : _GEN_2166;
  wire [13:0] _GEN_2168 = 14'h878 == index ? 14'h10 : _GEN_2167;
  wire [13:0] _GEN_2169 = 14'h879 == index ? 14'h10 : _GEN_2168;
  wire [13:0] _GEN_2170 = 14'h87a == index ? 14'h10 : _GEN_2169;
  wire [13:0] _GEN_2171 = 14'h87b == index ? 14'h10 : _GEN_2170;
  wire [13:0] _GEN_2172 = 14'h87c == index ? 14'h10 : _GEN_2171;
  wire [13:0] _GEN_2173 = 14'h87d == index ? 14'h10 : _GEN_2172;
  wire [13:0] _GEN_2174 = 14'h87e == index ? 14'h10 : _GEN_2173;
  wire [13:0] _GEN_2175 = 14'h87f == index ? 14'h10 : _GEN_2174;
  wire [13:0] _GEN_2176 = 14'h880 == index ? 14'h0 : _GEN_2175;
  wire [13:0] _GEN_2177 = 14'h881 == index ? 14'h880 : _GEN_2176;
  wire [13:0] _GEN_2178 = 14'h882 == index ? 14'h401 : _GEN_2177;
  wire [13:0] _GEN_2179 = 14'h883 == index ? 14'h282 : _GEN_2178;
  wire [13:0] _GEN_2180 = 14'h884 == index ? 14'h201 : _GEN_2179;
  wire [13:0] _GEN_2181 = 14'h885 == index ? 14'h182 : _GEN_2180;
  wire [13:0] _GEN_2182 = 14'h886 == index ? 14'h105 : _GEN_2181;
  wire [13:0] _GEN_2183 = 14'h887 == index ? 14'h103 : _GEN_2182;
  wire [13:0] _GEN_2184 = 14'h888 == index ? 14'h101 : _GEN_2183;
  wire [13:0] _GEN_2185 = 14'h889 == index ? 14'h88 : _GEN_2184;
  wire [13:0] _GEN_2186 = 14'h88a == index ? 14'h87 : _GEN_2185;
  wire [13:0] _GEN_2187 = 14'h88b == index ? 14'h86 : _GEN_2186;
  wire [13:0] _GEN_2188 = 14'h88c == index ? 14'h85 : _GEN_2187;
  wire [13:0] _GEN_2189 = 14'h88d == index ? 14'h84 : _GEN_2188;
  wire [13:0] _GEN_2190 = 14'h88e == index ? 14'h83 : _GEN_2189;
  wire [13:0] _GEN_2191 = 14'h88f == index ? 14'h82 : _GEN_2190;
  wire [13:0] _GEN_2192 = 14'h890 == index ? 14'h81 : _GEN_2191;
  wire [13:0] _GEN_2193 = 14'h891 == index ? 14'h80 : _GEN_2192;
  wire [13:0] _GEN_2194 = 14'h892 == index ? 14'h11 : _GEN_2193;
  wire [13:0] _GEN_2195 = 14'h893 == index ? 14'h11 : _GEN_2194;
  wire [13:0] _GEN_2196 = 14'h894 == index ? 14'h11 : _GEN_2195;
  wire [13:0] _GEN_2197 = 14'h895 == index ? 14'h11 : _GEN_2196;
  wire [13:0] _GEN_2198 = 14'h896 == index ? 14'h11 : _GEN_2197;
  wire [13:0] _GEN_2199 = 14'h897 == index ? 14'h11 : _GEN_2198;
  wire [13:0] _GEN_2200 = 14'h898 == index ? 14'h11 : _GEN_2199;
  wire [13:0] _GEN_2201 = 14'h899 == index ? 14'h11 : _GEN_2200;
  wire [13:0] _GEN_2202 = 14'h89a == index ? 14'h11 : _GEN_2201;
  wire [13:0] _GEN_2203 = 14'h89b == index ? 14'h11 : _GEN_2202;
  wire [13:0] _GEN_2204 = 14'h89c == index ? 14'h11 : _GEN_2203;
  wire [13:0] _GEN_2205 = 14'h89d == index ? 14'h11 : _GEN_2204;
  wire [13:0] _GEN_2206 = 14'h89e == index ? 14'h11 : _GEN_2205;
  wire [13:0] _GEN_2207 = 14'h89f == index ? 14'h11 : _GEN_2206;
  wire [13:0] _GEN_2208 = 14'h8a0 == index ? 14'h11 : _GEN_2207;
  wire [13:0] _GEN_2209 = 14'h8a1 == index ? 14'h11 : _GEN_2208;
  wire [13:0] _GEN_2210 = 14'h8a2 == index ? 14'h11 : _GEN_2209;
  wire [13:0] _GEN_2211 = 14'h8a3 == index ? 14'h11 : _GEN_2210;
  wire [13:0] _GEN_2212 = 14'h8a4 == index ? 14'h11 : _GEN_2211;
  wire [13:0] _GEN_2213 = 14'h8a5 == index ? 14'h11 : _GEN_2212;
  wire [13:0] _GEN_2214 = 14'h8a6 == index ? 14'h11 : _GEN_2213;
  wire [13:0] _GEN_2215 = 14'h8a7 == index ? 14'h11 : _GEN_2214;
  wire [13:0] _GEN_2216 = 14'h8a8 == index ? 14'h11 : _GEN_2215;
  wire [13:0] _GEN_2217 = 14'h8a9 == index ? 14'h11 : _GEN_2216;
  wire [13:0] _GEN_2218 = 14'h8aa == index ? 14'h11 : _GEN_2217;
  wire [13:0] _GEN_2219 = 14'h8ab == index ? 14'h11 : _GEN_2218;
  wire [13:0] _GEN_2220 = 14'h8ac == index ? 14'h11 : _GEN_2219;
  wire [13:0] _GEN_2221 = 14'h8ad == index ? 14'h11 : _GEN_2220;
  wire [13:0] _GEN_2222 = 14'h8ae == index ? 14'h11 : _GEN_2221;
  wire [13:0] _GEN_2223 = 14'h8af == index ? 14'h11 : _GEN_2222;
  wire [13:0] _GEN_2224 = 14'h8b0 == index ? 14'h11 : _GEN_2223;
  wire [13:0] _GEN_2225 = 14'h8b1 == index ? 14'h11 : _GEN_2224;
  wire [13:0] _GEN_2226 = 14'h8b2 == index ? 14'h11 : _GEN_2225;
  wire [13:0] _GEN_2227 = 14'h8b3 == index ? 14'h11 : _GEN_2226;
  wire [13:0] _GEN_2228 = 14'h8b4 == index ? 14'h11 : _GEN_2227;
  wire [13:0] _GEN_2229 = 14'h8b5 == index ? 14'h11 : _GEN_2228;
  wire [13:0] _GEN_2230 = 14'h8b6 == index ? 14'h11 : _GEN_2229;
  wire [13:0] _GEN_2231 = 14'h8b7 == index ? 14'h11 : _GEN_2230;
  wire [13:0] _GEN_2232 = 14'h8b8 == index ? 14'h11 : _GEN_2231;
  wire [13:0] _GEN_2233 = 14'h8b9 == index ? 14'h11 : _GEN_2232;
  wire [13:0] _GEN_2234 = 14'h8ba == index ? 14'h11 : _GEN_2233;
  wire [13:0] _GEN_2235 = 14'h8bb == index ? 14'h11 : _GEN_2234;
  wire [13:0] _GEN_2236 = 14'h8bc == index ? 14'h11 : _GEN_2235;
  wire [13:0] _GEN_2237 = 14'h8bd == index ? 14'h11 : _GEN_2236;
  wire [13:0] _GEN_2238 = 14'h8be == index ? 14'h11 : _GEN_2237;
  wire [13:0] _GEN_2239 = 14'h8bf == index ? 14'h11 : _GEN_2238;
  wire [13:0] _GEN_2240 = 14'h8c0 == index ? 14'h11 : _GEN_2239;
  wire [13:0] _GEN_2241 = 14'h8c1 == index ? 14'h11 : _GEN_2240;
  wire [13:0] _GEN_2242 = 14'h8c2 == index ? 14'h11 : _GEN_2241;
  wire [13:0] _GEN_2243 = 14'h8c3 == index ? 14'h11 : _GEN_2242;
  wire [13:0] _GEN_2244 = 14'h8c4 == index ? 14'h11 : _GEN_2243;
  wire [13:0] _GEN_2245 = 14'h8c5 == index ? 14'h11 : _GEN_2244;
  wire [13:0] _GEN_2246 = 14'h8c6 == index ? 14'h11 : _GEN_2245;
  wire [13:0] _GEN_2247 = 14'h8c7 == index ? 14'h11 : _GEN_2246;
  wire [13:0] _GEN_2248 = 14'h8c8 == index ? 14'h11 : _GEN_2247;
  wire [13:0] _GEN_2249 = 14'h8c9 == index ? 14'h11 : _GEN_2248;
  wire [13:0] _GEN_2250 = 14'h8ca == index ? 14'h11 : _GEN_2249;
  wire [13:0] _GEN_2251 = 14'h8cb == index ? 14'h11 : _GEN_2250;
  wire [13:0] _GEN_2252 = 14'h8cc == index ? 14'h11 : _GEN_2251;
  wire [13:0] _GEN_2253 = 14'h8cd == index ? 14'h11 : _GEN_2252;
  wire [13:0] _GEN_2254 = 14'h8ce == index ? 14'h11 : _GEN_2253;
  wire [13:0] _GEN_2255 = 14'h8cf == index ? 14'h11 : _GEN_2254;
  wire [13:0] _GEN_2256 = 14'h8d0 == index ? 14'h11 : _GEN_2255;
  wire [13:0] _GEN_2257 = 14'h8d1 == index ? 14'h11 : _GEN_2256;
  wire [13:0] _GEN_2258 = 14'h8d2 == index ? 14'h11 : _GEN_2257;
  wire [13:0] _GEN_2259 = 14'h8d3 == index ? 14'h11 : _GEN_2258;
  wire [13:0] _GEN_2260 = 14'h8d4 == index ? 14'h11 : _GEN_2259;
  wire [13:0] _GEN_2261 = 14'h8d5 == index ? 14'h11 : _GEN_2260;
  wire [13:0] _GEN_2262 = 14'h8d6 == index ? 14'h11 : _GEN_2261;
  wire [13:0] _GEN_2263 = 14'h8d7 == index ? 14'h11 : _GEN_2262;
  wire [13:0] _GEN_2264 = 14'h8d8 == index ? 14'h11 : _GEN_2263;
  wire [13:0] _GEN_2265 = 14'h8d9 == index ? 14'h11 : _GEN_2264;
  wire [13:0] _GEN_2266 = 14'h8da == index ? 14'h11 : _GEN_2265;
  wire [13:0] _GEN_2267 = 14'h8db == index ? 14'h11 : _GEN_2266;
  wire [13:0] _GEN_2268 = 14'h8dc == index ? 14'h11 : _GEN_2267;
  wire [13:0] _GEN_2269 = 14'h8dd == index ? 14'h11 : _GEN_2268;
  wire [13:0] _GEN_2270 = 14'h8de == index ? 14'h11 : _GEN_2269;
  wire [13:0] _GEN_2271 = 14'h8df == index ? 14'h11 : _GEN_2270;
  wire [13:0] _GEN_2272 = 14'h8e0 == index ? 14'h11 : _GEN_2271;
  wire [13:0] _GEN_2273 = 14'h8e1 == index ? 14'h11 : _GEN_2272;
  wire [13:0] _GEN_2274 = 14'h8e2 == index ? 14'h11 : _GEN_2273;
  wire [13:0] _GEN_2275 = 14'h8e3 == index ? 14'h11 : _GEN_2274;
  wire [13:0] _GEN_2276 = 14'h8e4 == index ? 14'h11 : _GEN_2275;
  wire [13:0] _GEN_2277 = 14'h8e5 == index ? 14'h11 : _GEN_2276;
  wire [13:0] _GEN_2278 = 14'h8e6 == index ? 14'h11 : _GEN_2277;
  wire [13:0] _GEN_2279 = 14'h8e7 == index ? 14'h11 : _GEN_2278;
  wire [13:0] _GEN_2280 = 14'h8e8 == index ? 14'h11 : _GEN_2279;
  wire [13:0] _GEN_2281 = 14'h8e9 == index ? 14'h11 : _GEN_2280;
  wire [13:0] _GEN_2282 = 14'h8ea == index ? 14'h11 : _GEN_2281;
  wire [13:0] _GEN_2283 = 14'h8eb == index ? 14'h11 : _GEN_2282;
  wire [13:0] _GEN_2284 = 14'h8ec == index ? 14'h11 : _GEN_2283;
  wire [13:0] _GEN_2285 = 14'h8ed == index ? 14'h11 : _GEN_2284;
  wire [13:0] _GEN_2286 = 14'h8ee == index ? 14'h11 : _GEN_2285;
  wire [13:0] _GEN_2287 = 14'h8ef == index ? 14'h11 : _GEN_2286;
  wire [13:0] _GEN_2288 = 14'h8f0 == index ? 14'h11 : _GEN_2287;
  wire [13:0] _GEN_2289 = 14'h8f1 == index ? 14'h11 : _GEN_2288;
  wire [13:0] _GEN_2290 = 14'h8f2 == index ? 14'h11 : _GEN_2289;
  wire [13:0] _GEN_2291 = 14'h8f3 == index ? 14'h11 : _GEN_2290;
  wire [13:0] _GEN_2292 = 14'h8f4 == index ? 14'h11 : _GEN_2291;
  wire [13:0] _GEN_2293 = 14'h8f5 == index ? 14'h11 : _GEN_2292;
  wire [13:0] _GEN_2294 = 14'h8f6 == index ? 14'h11 : _GEN_2293;
  wire [13:0] _GEN_2295 = 14'h8f7 == index ? 14'h11 : _GEN_2294;
  wire [13:0] _GEN_2296 = 14'h8f8 == index ? 14'h11 : _GEN_2295;
  wire [13:0] _GEN_2297 = 14'h8f9 == index ? 14'h11 : _GEN_2296;
  wire [13:0] _GEN_2298 = 14'h8fa == index ? 14'h11 : _GEN_2297;
  wire [13:0] _GEN_2299 = 14'h8fb == index ? 14'h11 : _GEN_2298;
  wire [13:0] _GEN_2300 = 14'h8fc == index ? 14'h11 : _GEN_2299;
  wire [13:0] _GEN_2301 = 14'h8fd == index ? 14'h11 : _GEN_2300;
  wire [13:0] _GEN_2302 = 14'h8fe == index ? 14'h11 : _GEN_2301;
  wire [13:0] _GEN_2303 = 14'h8ff == index ? 14'h11 : _GEN_2302;
  wire [13:0] _GEN_2304 = 14'h900 == index ? 14'h0 : _GEN_2303;
  wire [13:0] _GEN_2305 = 14'h901 == index ? 14'h900 : _GEN_2304;
  wire [13:0] _GEN_2306 = 14'h902 == index ? 14'h480 : _GEN_2305;
  wire [13:0] _GEN_2307 = 14'h903 == index ? 14'h300 : _GEN_2306;
  wire [13:0] _GEN_2308 = 14'h904 == index ? 14'h202 : _GEN_2307;
  wire [13:0] _GEN_2309 = 14'h905 == index ? 14'h183 : _GEN_2308;
  wire [13:0] _GEN_2310 = 14'h906 == index ? 14'h180 : _GEN_2309;
  wire [13:0] _GEN_2311 = 14'h907 == index ? 14'h104 : _GEN_2310;
  wire [13:0] _GEN_2312 = 14'h908 == index ? 14'h102 : _GEN_2311;
  wire [13:0] _GEN_2313 = 14'h909 == index ? 14'h100 : _GEN_2312;
  wire [13:0] _GEN_2314 = 14'h90a == index ? 14'h88 : _GEN_2313;
  wire [13:0] _GEN_2315 = 14'h90b == index ? 14'h87 : _GEN_2314;
  wire [13:0] _GEN_2316 = 14'h90c == index ? 14'h86 : _GEN_2315;
  wire [13:0] _GEN_2317 = 14'h90d == index ? 14'h85 : _GEN_2316;
  wire [13:0] _GEN_2318 = 14'h90e == index ? 14'h84 : _GEN_2317;
  wire [13:0] _GEN_2319 = 14'h90f == index ? 14'h83 : _GEN_2318;
  wire [13:0] _GEN_2320 = 14'h910 == index ? 14'h82 : _GEN_2319;
  wire [13:0] _GEN_2321 = 14'h911 == index ? 14'h81 : _GEN_2320;
  wire [13:0] _GEN_2322 = 14'h912 == index ? 14'h80 : _GEN_2321;
  wire [13:0] _GEN_2323 = 14'h913 == index ? 14'h12 : _GEN_2322;
  wire [13:0] _GEN_2324 = 14'h914 == index ? 14'h12 : _GEN_2323;
  wire [13:0] _GEN_2325 = 14'h915 == index ? 14'h12 : _GEN_2324;
  wire [13:0] _GEN_2326 = 14'h916 == index ? 14'h12 : _GEN_2325;
  wire [13:0] _GEN_2327 = 14'h917 == index ? 14'h12 : _GEN_2326;
  wire [13:0] _GEN_2328 = 14'h918 == index ? 14'h12 : _GEN_2327;
  wire [13:0] _GEN_2329 = 14'h919 == index ? 14'h12 : _GEN_2328;
  wire [13:0] _GEN_2330 = 14'h91a == index ? 14'h12 : _GEN_2329;
  wire [13:0] _GEN_2331 = 14'h91b == index ? 14'h12 : _GEN_2330;
  wire [13:0] _GEN_2332 = 14'h91c == index ? 14'h12 : _GEN_2331;
  wire [13:0] _GEN_2333 = 14'h91d == index ? 14'h12 : _GEN_2332;
  wire [13:0] _GEN_2334 = 14'h91e == index ? 14'h12 : _GEN_2333;
  wire [13:0] _GEN_2335 = 14'h91f == index ? 14'h12 : _GEN_2334;
  wire [13:0] _GEN_2336 = 14'h920 == index ? 14'h12 : _GEN_2335;
  wire [13:0] _GEN_2337 = 14'h921 == index ? 14'h12 : _GEN_2336;
  wire [13:0] _GEN_2338 = 14'h922 == index ? 14'h12 : _GEN_2337;
  wire [13:0] _GEN_2339 = 14'h923 == index ? 14'h12 : _GEN_2338;
  wire [13:0] _GEN_2340 = 14'h924 == index ? 14'h12 : _GEN_2339;
  wire [13:0] _GEN_2341 = 14'h925 == index ? 14'h12 : _GEN_2340;
  wire [13:0] _GEN_2342 = 14'h926 == index ? 14'h12 : _GEN_2341;
  wire [13:0] _GEN_2343 = 14'h927 == index ? 14'h12 : _GEN_2342;
  wire [13:0] _GEN_2344 = 14'h928 == index ? 14'h12 : _GEN_2343;
  wire [13:0] _GEN_2345 = 14'h929 == index ? 14'h12 : _GEN_2344;
  wire [13:0] _GEN_2346 = 14'h92a == index ? 14'h12 : _GEN_2345;
  wire [13:0] _GEN_2347 = 14'h92b == index ? 14'h12 : _GEN_2346;
  wire [13:0] _GEN_2348 = 14'h92c == index ? 14'h12 : _GEN_2347;
  wire [13:0] _GEN_2349 = 14'h92d == index ? 14'h12 : _GEN_2348;
  wire [13:0] _GEN_2350 = 14'h92e == index ? 14'h12 : _GEN_2349;
  wire [13:0] _GEN_2351 = 14'h92f == index ? 14'h12 : _GEN_2350;
  wire [13:0] _GEN_2352 = 14'h930 == index ? 14'h12 : _GEN_2351;
  wire [13:0] _GEN_2353 = 14'h931 == index ? 14'h12 : _GEN_2352;
  wire [13:0] _GEN_2354 = 14'h932 == index ? 14'h12 : _GEN_2353;
  wire [13:0] _GEN_2355 = 14'h933 == index ? 14'h12 : _GEN_2354;
  wire [13:0] _GEN_2356 = 14'h934 == index ? 14'h12 : _GEN_2355;
  wire [13:0] _GEN_2357 = 14'h935 == index ? 14'h12 : _GEN_2356;
  wire [13:0] _GEN_2358 = 14'h936 == index ? 14'h12 : _GEN_2357;
  wire [13:0] _GEN_2359 = 14'h937 == index ? 14'h12 : _GEN_2358;
  wire [13:0] _GEN_2360 = 14'h938 == index ? 14'h12 : _GEN_2359;
  wire [13:0] _GEN_2361 = 14'h939 == index ? 14'h12 : _GEN_2360;
  wire [13:0] _GEN_2362 = 14'h93a == index ? 14'h12 : _GEN_2361;
  wire [13:0] _GEN_2363 = 14'h93b == index ? 14'h12 : _GEN_2362;
  wire [13:0] _GEN_2364 = 14'h93c == index ? 14'h12 : _GEN_2363;
  wire [13:0] _GEN_2365 = 14'h93d == index ? 14'h12 : _GEN_2364;
  wire [13:0] _GEN_2366 = 14'h93e == index ? 14'h12 : _GEN_2365;
  wire [13:0] _GEN_2367 = 14'h93f == index ? 14'h12 : _GEN_2366;
  wire [13:0] _GEN_2368 = 14'h940 == index ? 14'h12 : _GEN_2367;
  wire [13:0] _GEN_2369 = 14'h941 == index ? 14'h12 : _GEN_2368;
  wire [13:0] _GEN_2370 = 14'h942 == index ? 14'h12 : _GEN_2369;
  wire [13:0] _GEN_2371 = 14'h943 == index ? 14'h12 : _GEN_2370;
  wire [13:0] _GEN_2372 = 14'h944 == index ? 14'h12 : _GEN_2371;
  wire [13:0] _GEN_2373 = 14'h945 == index ? 14'h12 : _GEN_2372;
  wire [13:0] _GEN_2374 = 14'h946 == index ? 14'h12 : _GEN_2373;
  wire [13:0] _GEN_2375 = 14'h947 == index ? 14'h12 : _GEN_2374;
  wire [13:0] _GEN_2376 = 14'h948 == index ? 14'h12 : _GEN_2375;
  wire [13:0] _GEN_2377 = 14'h949 == index ? 14'h12 : _GEN_2376;
  wire [13:0] _GEN_2378 = 14'h94a == index ? 14'h12 : _GEN_2377;
  wire [13:0] _GEN_2379 = 14'h94b == index ? 14'h12 : _GEN_2378;
  wire [13:0] _GEN_2380 = 14'h94c == index ? 14'h12 : _GEN_2379;
  wire [13:0] _GEN_2381 = 14'h94d == index ? 14'h12 : _GEN_2380;
  wire [13:0] _GEN_2382 = 14'h94e == index ? 14'h12 : _GEN_2381;
  wire [13:0] _GEN_2383 = 14'h94f == index ? 14'h12 : _GEN_2382;
  wire [13:0] _GEN_2384 = 14'h950 == index ? 14'h12 : _GEN_2383;
  wire [13:0] _GEN_2385 = 14'h951 == index ? 14'h12 : _GEN_2384;
  wire [13:0] _GEN_2386 = 14'h952 == index ? 14'h12 : _GEN_2385;
  wire [13:0] _GEN_2387 = 14'h953 == index ? 14'h12 : _GEN_2386;
  wire [13:0] _GEN_2388 = 14'h954 == index ? 14'h12 : _GEN_2387;
  wire [13:0] _GEN_2389 = 14'h955 == index ? 14'h12 : _GEN_2388;
  wire [13:0] _GEN_2390 = 14'h956 == index ? 14'h12 : _GEN_2389;
  wire [13:0] _GEN_2391 = 14'h957 == index ? 14'h12 : _GEN_2390;
  wire [13:0] _GEN_2392 = 14'h958 == index ? 14'h12 : _GEN_2391;
  wire [13:0] _GEN_2393 = 14'h959 == index ? 14'h12 : _GEN_2392;
  wire [13:0] _GEN_2394 = 14'h95a == index ? 14'h12 : _GEN_2393;
  wire [13:0] _GEN_2395 = 14'h95b == index ? 14'h12 : _GEN_2394;
  wire [13:0] _GEN_2396 = 14'h95c == index ? 14'h12 : _GEN_2395;
  wire [13:0] _GEN_2397 = 14'h95d == index ? 14'h12 : _GEN_2396;
  wire [13:0] _GEN_2398 = 14'h95e == index ? 14'h12 : _GEN_2397;
  wire [13:0] _GEN_2399 = 14'h95f == index ? 14'h12 : _GEN_2398;
  wire [13:0] _GEN_2400 = 14'h960 == index ? 14'h12 : _GEN_2399;
  wire [13:0] _GEN_2401 = 14'h961 == index ? 14'h12 : _GEN_2400;
  wire [13:0] _GEN_2402 = 14'h962 == index ? 14'h12 : _GEN_2401;
  wire [13:0] _GEN_2403 = 14'h963 == index ? 14'h12 : _GEN_2402;
  wire [13:0] _GEN_2404 = 14'h964 == index ? 14'h12 : _GEN_2403;
  wire [13:0] _GEN_2405 = 14'h965 == index ? 14'h12 : _GEN_2404;
  wire [13:0] _GEN_2406 = 14'h966 == index ? 14'h12 : _GEN_2405;
  wire [13:0] _GEN_2407 = 14'h967 == index ? 14'h12 : _GEN_2406;
  wire [13:0] _GEN_2408 = 14'h968 == index ? 14'h12 : _GEN_2407;
  wire [13:0] _GEN_2409 = 14'h969 == index ? 14'h12 : _GEN_2408;
  wire [13:0] _GEN_2410 = 14'h96a == index ? 14'h12 : _GEN_2409;
  wire [13:0] _GEN_2411 = 14'h96b == index ? 14'h12 : _GEN_2410;
  wire [13:0] _GEN_2412 = 14'h96c == index ? 14'h12 : _GEN_2411;
  wire [13:0] _GEN_2413 = 14'h96d == index ? 14'h12 : _GEN_2412;
  wire [13:0] _GEN_2414 = 14'h96e == index ? 14'h12 : _GEN_2413;
  wire [13:0] _GEN_2415 = 14'h96f == index ? 14'h12 : _GEN_2414;
  wire [13:0] _GEN_2416 = 14'h970 == index ? 14'h12 : _GEN_2415;
  wire [13:0] _GEN_2417 = 14'h971 == index ? 14'h12 : _GEN_2416;
  wire [13:0] _GEN_2418 = 14'h972 == index ? 14'h12 : _GEN_2417;
  wire [13:0] _GEN_2419 = 14'h973 == index ? 14'h12 : _GEN_2418;
  wire [13:0] _GEN_2420 = 14'h974 == index ? 14'h12 : _GEN_2419;
  wire [13:0] _GEN_2421 = 14'h975 == index ? 14'h12 : _GEN_2420;
  wire [13:0] _GEN_2422 = 14'h976 == index ? 14'h12 : _GEN_2421;
  wire [13:0] _GEN_2423 = 14'h977 == index ? 14'h12 : _GEN_2422;
  wire [13:0] _GEN_2424 = 14'h978 == index ? 14'h12 : _GEN_2423;
  wire [13:0] _GEN_2425 = 14'h979 == index ? 14'h12 : _GEN_2424;
  wire [13:0] _GEN_2426 = 14'h97a == index ? 14'h12 : _GEN_2425;
  wire [13:0] _GEN_2427 = 14'h97b == index ? 14'h12 : _GEN_2426;
  wire [13:0] _GEN_2428 = 14'h97c == index ? 14'h12 : _GEN_2427;
  wire [13:0] _GEN_2429 = 14'h97d == index ? 14'h12 : _GEN_2428;
  wire [13:0] _GEN_2430 = 14'h97e == index ? 14'h12 : _GEN_2429;
  wire [13:0] _GEN_2431 = 14'h97f == index ? 14'h12 : _GEN_2430;
  wire [13:0] _GEN_2432 = 14'h980 == index ? 14'h0 : _GEN_2431;
  wire [13:0] _GEN_2433 = 14'h981 == index ? 14'h980 : _GEN_2432;
  wire [13:0] _GEN_2434 = 14'h982 == index ? 14'h481 : _GEN_2433;
  wire [13:0] _GEN_2435 = 14'h983 == index ? 14'h301 : _GEN_2434;
  wire [13:0] _GEN_2436 = 14'h984 == index ? 14'h203 : _GEN_2435;
  wire [13:0] _GEN_2437 = 14'h985 == index ? 14'h184 : _GEN_2436;
  wire [13:0] _GEN_2438 = 14'h986 == index ? 14'h181 : _GEN_2437;
  wire [13:0] _GEN_2439 = 14'h987 == index ? 14'h105 : _GEN_2438;
  wire [13:0] _GEN_2440 = 14'h988 == index ? 14'h103 : _GEN_2439;
  wire [13:0] _GEN_2441 = 14'h989 == index ? 14'h101 : _GEN_2440;
  wire [13:0] _GEN_2442 = 14'h98a == index ? 14'h89 : _GEN_2441;
  wire [13:0] _GEN_2443 = 14'h98b == index ? 14'h88 : _GEN_2442;
  wire [13:0] _GEN_2444 = 14'h98c == index ? 14'h87 : _GEN_2443;
  wire [13:0] _GEN_2445 = 14'h98d == index ? 14'h86 : _GEN_2444;
  wire [13:0] _GEN_2446 = 14'h98e == index ? 14'h85 : _GEN_2445;
  wire [13:0] _GEN_2447 = 14'h98f == index ? 14'h84 : _GEN_2446;
  wire [13:0] _GEN_2448 = 14'h990 == index ? 14'h83 : _GEN_2447;
  wire [13:0] _GEN_2449 = 14'h991 == index ? 14'h82 : _GEN_2448;
  wire [13:0] _GEN_2450 = 14'h992 == index ? 14'h81 : _GEN_2449;
  wire [13:0] _GEN_2451 = 14'h993 == index ? 14'h80 : _GEN_2450;
  wire [13:0] _GEN_2452 = 14'h994 == index ? 14'h13 : _GEN_2451;
  wire [13:0] _GEN_2453 = 14'h995 == index ? 14'h13 : _GEN_2452;
  wire [13:0] _GEN_2454 = 14'h996 == index ? 14'h13 : _GEN_2453;
  wire [13:0] _GEN_2455 = 14'h997 == index ? 14'h13 : _GEN_2454;
  wire [13:0] _GEN_2456 = 14'h998 == index ? 14'h13 : _GEN_2455;
  wire [13:0] _GEN_2457 = 14'h999 == index ? 14'h13 : _GEN_2456;
  wire [13:0] _GEN_2458 = 14'h99a == index ? 14'h13 : _GEN_2457;
  wire [13:0] _GEN_2459 = 14'h99b == index ? 14'h13 : _GEN_2458;
  wire [13:0] _GEN_2460 = 14'h99c == index ? 14'h13 : _GEN_2459;
  wire [13:0] _GEN_2461 = 14'h99d == index ? 14'h13 : _GEN_2460;
  wire [13:0] _GEN_2462 = 14'h99e == index ? 14'h13 : _GEN_2461;
  wire [13:0] _GEN_2463 = 14'h99f == index ? 14'h13 : _GEN_2462;
  wire [13:0] _GEN_2464 = 14'h9a0 == index ? 14'h13 : _GEN_2463;
  wire [13:0] _GEN_2465 = 14'h9a1 == index ? 14'h13 : _GEN_2464;
  wire [13:0] _GEN_2466 = 14'h9a2 == index ? 14'h13 : _GEN_2465;
  wire [13:0] _GEN_2467 = 14'h9a3 == index ? 14'h13 : _GEN_2466;
  wire [13:0] _GEN_2468 = 14'h9a4 == index ? 14'h13 : _GEN_2467;
  wire [13:0] _GEN_2469 = 14'h9a5 == index ? 14'h13 : _GEN_2468;
  wire [13:0] _GEN_2470 = 14'h9a6 == index ? 14'h13 : _GEN_2469;
  wire [13:0] _GEN_2471 = 14'h9a7 == index ? 14'h13 : _GEN_2470;
  wire [13:0] _GEN_2472 = 14'h9a8 == index ? 14'h13 : _GEN_2471;
  wire [13:0] _GEN_2473 = 14'h9a9 == index ? 14'h13 : _GEN_2472;
  wire [13:0] _GEN_2474 = 14'h9aa == index ? 14'h13 : _GEN_2473;
  wire [13:0] _GEN_2475 = 14'h9ab == index ? 14'h13 : _GEN_2474;
  wire [13:0] _GEN_2476 = 14'h9ac == index ? 14'h13 : _GEN_2475;
  wire [13:0] _GEN_2477 = 14'h9ad == index ? 14'h13 : _GEN_2476;
  wire [13:0] _GEN_2478 = 14'h9ae == index ? 14'h13 : _GEN_2477;
  wire [13:0] _GEN_2479 = 14'h9af == index ? 14'h13 : _GEN_2478;
  wire [13:0] _GEN_2480 = 14'h9b0 == index ? 14'h13 : _GEN_2479;
  wire [13:0] _GEN_2481 = 14'h9b1 == index ? 14'h13 : _GEN_2480;
  wire [13:0] _GEN_2482 = 14'h9b2 == index ? 14'h13 : _GEN_2481;
  wire [13:0] _GEN_2483 = 14'h9b3 == index ? 14'h13 : _GEN_2482;
  wire [13:0] _GEN_2484 = 14'h9b4 == index ? 14'h13 : _GEN_2483;
  wire [13:0] _GEN_2485 = 14'h9b5 == index ? 14'h13 : _GEN_2484;
  wire [13:0] _GEN_2486 = 14'h9b6 == index ? 14'h13 : _GEN_2485;
  wire [13:0] _GEN_2487 = 14'h9b7 == index ? 14'h13 : _GEN_2486;
  wire [13:0] _GEN_2488 = 14'h9b8 == index ? 14'h13 : _GEN_2487;
  wire [13:0] _GEN_2489 = 14'h9b9 == index ? 14'h13 : _GEN_2488;
  wire [13:0] _GEN_2490 = 14'h9ba == index ? 14'h13 : _GEN_2489;
  wire [13:0] _GEN_2491 = 14'h9bb == index ? 14'h13 : _GEN_2490;
  wire [13:0] _GEN_2492 = 14'h9bc == index ? 14'h13 : _GEN_2491;
  wire [13:0] _GEN_2493 = 14'h9bd == index ? 14'h13 : _GEN_2492;
  wire [13:0] _GEN_2494 = 14'h9be == index ? 14'h13 : _GEN_2493;
  wire [13:0] _GEN_2495 = 14'h9bf == index ? 14'h13 : _GEN_2494;
  wire [13:0] _GEN_2496 = 14'h9c0 == index ? 14'h13 : _GEN_2495;
  wire [13:0] _GEN_2497 = 14'h9c1 == index ? 14'h13 : _GEN_2496;
  wire [13:0] _GEN_2498 = 14'h9c2 == index ? 14'h13 : _GEN_2497;
  wire [13:0] _GEN_2499 = 14'h9c3 == index ? 14'h13 : _GEN_2498;
  wire [13:0] _GEN_2500 = 14'h9c4 == index ? 14'h13 : _GEN_2499;
  wire [13:0] _GEN_2501 = 14'h9c5 == index ? 14'h13 : _GEN_2500;
  wire [13:0] _GEN_2502 = 14'h9c6 == index ? 14'h13 : _GEN_2501;
  wire [13:0] _GEN_2503 = 14'h9c7 == index ? 14'h13 : _GEN_2502;
  wire [13:0] _GEN_2504 = 14'h9c8 == index ? 14'h13 : _GEN_2503;
  wire [13:0] _GEN_2505 = 14'h9c9 == index ? 14'h13 : _GEN_2504;
  wire [13:0] _GEN_2506 = 14'h9ca == index ? 14'h13 : _GEN_2505;
  wire [13:0] _GEN_2507 = 14'h9cb == index ? 14'h13 : _GEN_2506;
  wire [13:0] _GEN_2508 = 14'h9cc == index ? 14'h13 : _GEN_2507;
  wire [13:0] _GEN_2509 = 14'h9cd == index ? 14'h13 : _GEN_2508;
  wire [13:0] _GEN_2510 = 14'h9ce == index ? 14'h13 : _GEN_2509;
  wire [13:0] _GEN_2511 = 14'h9cf == index ? 14'h13 : _GEN_2510;
  wire [13:0] _GEN_2512 = 14'h9d0 == index ? 14'h13 : _GEN_2511;
  wire [13:0] _GEN_2513 = 14'h9d1 == index ? 14'h13 : _GEN_2512;
  wire [13:0] _GEN_2514 = 14'h9d2 == index ? 14'h13 : _GEN_2513;
  wire [13:0] _GEN_2515 = 14'h9d3 == index ? 14'h13 : _GEN_2514;
  wire [13:0] _GEN_2516 = 14'h9d4 == index ? 14'h13 : _GEN_2515;
  wire [13:0] _GEN_2517 = 14'h9d5 == index ? 14'h13 : _GEN_2516;
  wire [13:0] _GEN_2518 = 14'h9d6 == index ? 14'h13 : _GEN_2517;
  wire [13:0] _GEN_2519 = 14'h9d7 == index ? 14'h13 : _GEN_2518;
  wire [13:0] _GEN_2520 = 14'h9d8 == index ? 14'h13 : _GEN_2519;
  wire [13:0] _GEN_2521 = 14'h9d9 == index ? 14'h13 : _GEN_2520;
  wire [13:0] _GEN_2522 = 14'h9da == index ? 14'h13 : _GEN_2521;
  wire [13:0] _GEN_2523 = 14'h9db == index ? 14'h13 : _GEN_2522;
  wire [13:0] _GEN_2524 = 14'h9dc == index ? 14'h13 : _GEN_2523;
  wire [13:0] _GEN_2525 = 14'h9dd == index ? 14'h13 : _GEN_2524;
  wire [13:0] _GEN_2526 = 14'h9de == index ? 14'h13 : _GEN_2525;
  wire [13:0] _GEN_2527 = 14'h9df == index ? 14'h13 : _GEN_2526;
  wire [13:0] _GEN_2528 = 14'h9e0 == index ? 14'h13 : _GEN_2527;
  wire [13:0] _GEN_2529 = 14'h9e1 == index ? 14'h13 : _GEN_2528;
  wire [13:0] _GEN_2530 = 14'h9e2 == index ? 14'h13 : _GEN_2529;
  wire [13:0] _GEN_2531 = 14'h9e3 == index ? 14'h13 : _GEN_2530;
  wire [13:0] _GEN_2532 = 14'h9e4 == index ? 14'h13 : _GEN_2531;
  wire [13:0] _GEN_2533 = 14'h9e5 == index ? 14'h13 : _GEN_2532;
  wire [13:0] _GEN_2534 = 14'h9e6 == index ? 14'h13 : _GEN_2533;
  wire [13:0] _GEN_2535 = 14'h9e7 == index ? 14'h13 : _GEN_2534;
  wire [13:0] _GEN_2536 = 14'h9e8 == index ? 14'h13 : _GEN_2535;
  wire [13:0] _GEN_2537 = 14'h9e9 == index ? 14'h13 : _GEN_2536;
  wire [13:0] _GEN_2538 = 14'h9ea == index ? 14'h13 : _GEN_2537;
  wire [13:0] _GEN_2539 = 14'h9eb == index ? 14'h13 : _GEN_2538;
  wire [13:0] _GEN_2540 = 14'h9ec == index ? 14'h13 : _GEN_2539;
  wire [13:0] _GEN_2541 = 14'h9ed == index ? 14'h13 : _GEN_2540;
  wire [13:0] _GEN_2542 = 14'h9ee == index ? 14'h13 : _GEN_2541;
  wire [13:0] _GEN_2543 = 14'h9ef == index ? 14'h13 : _GEN_2542;
  wire [13:0] _GEN_2544 = 14'h9f0 == index ? 14'h13 : _GEN_2543;
  wire [13:0] _GEN_2545 = 14'h9f1 == index ? 14'h13 : _GEN_2544;
  wire [13:0] _GEN_2546 = 14'h9f2 == index ? 14'h13 : _GEN_2545;
  wire [13:0] _GEN_2547 = 14'h9f3 == index ? 14'h13 : _GEN_2546;
  wire [13:0] _GEN_2548 = 14'h9f4 == index ? 14'h13 : _GEN_2547;
  wire [13:0] _GEN_2549 = 14'h9f5 == index ? 14'h13 : _GEN_2548;
  wire [13:0] _GEN_2550 = 14'h9f6 == index ? 14'h13 : _GEN_2549;
  wire [13:0] _GEN_2551 = 14'h9f7 == index ? 14'h13 : _GEN_2550;
  wire [13:0] _GEN_2552 = 14'h9f8 == index ? 14'h13 : _GEN_2551;
  wire [13:0] _GEN_2553 = 14'h9f9 == index ? 14'h13 : _GEN_2552;
  wire [13:0] _GEN_2554 = 14'h9fa == index ? 14'h13 : _GEN_2553;
  wire [13:0] _GEN_2555 = 14'h9fb == index ? 14'h13 : _GEN_2554;
  wire [13:0] _GEN_2556 = 14'h9fc == index ? 14'h13 : _GEN_2555;
  wire [13:0] _GEN_2557 = 14'h9fd == index ? 14'h13 : _GEN_2556;
  wire [13:0] _GEN_2558 = 14'h9fe == index ? 14'h13 : _GEN_2557;
  wire [13:0] _GEN_2559 = 14'h9ff == index ? 14'h13 : _GEN_2558;
  wire [13:0] _GEN_2560 = 14'ha00 == index ? 14'h0 : _GEN_2559;
  wire [13:0] _GEN_2561 = 14'ha01 == index ? 14'ha00 : _GEN_2560;
  wire [13:0] _GEN_2562 = 14'ha02 == index ? 14'h500 : _GEN_2561;
  wire [13:0] _GEN_2563 = 14'ha03 == index ? 14'h302 : _GEN_2562;
  wire [13:0] _GEN_2564 = 14'ha04 == index ? 14'h280 : _GEN_2563;
  wire [13:0] _GEN_2565 = 14'ha05 == index ? 14'h200 : _GEN_2564;
  wire [13:0] _GEN_2566 = 14'ha06 == index ? 14'h182 : _GEN_2565;
  wire [13:0] _GEN_2567 = 14'ha07 == index ? 14'h106 : _GEN_2566;
  wire [13:0] _GEN_2568 = 14'ha08 == index ? 14'h104 : _GEN_2567;
  wire [13:0] _GEN_2569 = 14'ha09 == index ? 14'h102 : _GEN_2568;
  wire [13:0] _GEN_2570 = 14'ha0a == index ? 14'h100 : _GEN_2569;
  wire [13:0] _GEN_2571 = 14'ha0b == index ? 14'h89 : _GEN_2570;
  wire [13:0] _GEN_2572 = 14'ha0c == index ? 14'h88 : _GEN_2571;
  wire [13:0] _GEN_2573 = 14'ha0d == index ? 14'h87 : _GEN_2572;
  wire [13:0] _GEN_2574 = 14'ha0e == index ? 14'h86 : _GEN_2573;
  wire [13:0] _GEN_2575 = 14'ha0f == index ? 14'h85 : _GEN_2574;
  wire [13:0] _GEN_2576 = 14'ha10 == index ? 14'h84 : _GEN_2575;
  wire [13:0] _GEN_2577 = 14'ha11 == index ? 14'h83 : _GEN_2576;
  wire [13:0] _GEN_2578 = 14'ha12 == index ? 14'h82 : _GEN_2577;
  wire [13:0] _GEN_2579 = 14'ha13 == index ? 14'h81 : _GEN_2578;
  wire [13:0] _GEN_2580 = 14'ha14 == index ? 14'h80 : _GEN_2579;
  wire [13:0] _GEN_2581 = 14'ha15 == index ? 14'h14 : _GEN_2580;
  wire [13:0] _GEN_2582 = 14'ha16 == index ? 14'h14 : _GEN_2581;
  wire [13:0] _GEN_2583 = 14'ha17 == index ? 14'h14 : _GEN_2582;
  wire [13:0] _GEN_2584 = 14'ha18 == index ? 14'h14 : _GEN_2583;
  wire [13:0] _GEN_2585 = 14'ha19 == index ? 14'h14 : _GEN_2584;
  wire [13:0] _GEN_2586 = 14'ha1a == index ? 14'h14 : _GEN_2585;
  wire [13:0] _GEN_2587 = 14'ha1b == index ? 14'h14 : _GEN_2586;
  wire [13:0] _GEN_2588 = 14'ha1c == index ? 14'h14 : _GEN_2587;
  wire [13:0] _GEN_2589 = 14'ha1d == index ? 14'h14 : _GEN_2588;
  wire [13:0] _GEN_2590 = 14'ha1e == index ? 14'h14 : _GEN_2589;
  wire [13:0] _GEN_2591 = 14'ha1f == index ? 14'h14 : _GEN_2590;
  wire [13:0] _GEN_2592 = 14'ha20 == index ? 14'h14 : _GEN_2591;
  wire [13:0] _GEN_2593 = 14'ha21 == index ? 14'h14 : _GEN_2592;
  wire [13:0] _GEN_2594 = 14'ha22 == index ? 14'h14 : _GEN_2593;
  wire [13:0] _GEN_2595 = 14'ha23 == index ? 14'h14 : _GEN_2594;
  wire [13:0] _GEN_2596 = 14'ha24 == index ? 14'h14 : _GEN_2595;
  wire [13:0] _GEN_2597 = 14'ha25 == index ? 14'h14 : _GEN_2596;
  wire [13:0] _GEN_2598 = 14'ha26 == index ? 14'h14 : _GEN_2597;
  wire [13:0] _GEN_2599 = 14'ha27 == index ? 14'h14 : _GEN_2598;
  wire [13:0] _GEN_2600 = 14'ha28 == index ? 14'h14 : _GEN_2599;
  wire [13:0] _GEN_2601 = 14'ha29 == index ? 14'h14 : _GEN_2600;
  wire [13:0] _GEN_2602 = 14'ha2a == index ? 14'h14 : _GEN_2601;
  wire [13:0] _GEN_2603 = 14'ha2b == index ? 14'h14 : _GEN_2602;
  wire [13:0] _GEN_2604 = 14'ha2c == index ? 14'h14 : _GEN_2603;
  wire [13:0] _GEN_2605 = 14'ha2d == index ? 14'h14 : _GEN_2604;
  wire [13:0] _GEN_2606 = 14'ha2e == index ? 14'h14 : _GEN_2605;
  wire [13:0] _GEN_2607 = 14'ha2f == index ? 14'h14 : _GEN_2606;
  wire [13:0] _GEN_2608 = 14'ha30 == index ? 14'h14 : _GEN_2607;
  wire [13:0] _GEN_2609 = 14'ha31 == index ? 14'h14 : _GEN_2608;
  wire [13:0] _GEN_2610 = 14'ha32 == index ? 14'h14 : _GEN_2609;
  wire [13:0] _GEN_2611 = 14'ha33 == index ? 14'h14 : _GEN_2610;
  wire [13:0] _GEN_2612 = 14'ha34 == index ? 14'h14 : _GEN_2611;
  wire [13:0] _GEN_2613 = 14'ha35 == index ? 14'h14 : _GEN_2612;
  wire [13:0] _GEN_2614 = 14'ha36 == index ? 14'h14 : _GEN_2613;
  wire [13:0] _GEN_2615 = 14'ha37 == index ? 14'h14 : _GEN_2614;
  wire [13:0] _GEN_2616 = 14'ha38 == index ? 14'h14 : _GEN_2615;
  wire [13:0] _GEN_2617 = 14'ha39 == index ? 14'h14 : _GEN_2616;
  wire [13:0] _GEN_2618 = 14'ha3a == index ? 14'h14 : _GEN_2617;
  wire [13:0] _GEN_2619 = 14'ha3b == index ? 14'h14 : _GEN_2618;
  wire [13:0] _GEN_2620 = 14'ha3c == index ? 14'h14 : _GEN_2619;
  wire [13:0] _GEN_2621 = 14'ha3d == index ? 14'h14 : _GEN_2620;
  wire [13:0] _GEN_2622 = 14'ha3e == index ? 14'h14 : _GEN_2621;
  wire [13:0] _GEN_2623 = 14'ha3f == index ? 14'h14 : _GEN_2622;
  wire [13:0] _GEN_2624 = 14'ha40 == index ? 14'h14 : _GEN_2623;
  wire [13:0] _GEN_2625 = 14'ha41 == index ? 14'h14 : _GEN_2624;
  wire [13:0] _GEN_2626 = 14'ha42 == index ? 14'h14 : _GEN_2625;
  wire [13:0] _GEN_2627 = 14'ha43 == index ? 14'h14 : _GEN_2626;
  wire [13:0] _GEN_2628 = 14'ha44 == index ? 14'h14 : _GEN_2627;
  wire [13:0] _GEN_2629 = 14'ha45 == index ? 14'h14 : _GEN_2628;
  wire [13:0] _GEN_2630 = 14'ha46 == index ? 14'h14 : _GEN_2629;
  wire [13:0] _GEN_2631 = 14'ha47 == index ? 14'h14 : _GEN_2630;
  wire [13:0] _GEN_2632 = 14'ha48 == index ? 14'h14 : _GEN_2631;
  wire [13:0] _GEN_2633 = 14'ha49 == index ? 14'h14 : _GEN_2632;
  wire [13:0] _GEN_2634 = 14'ha4a == index ? 14'h14 : _GEN_2633;
  wire [13:0] _GEN_2635 = 14'ha4b == index ? 14'h14 : _GEN_2634;
  wire [13:0] _GEN_2636 = 14'ha4c == index ? 14'h14 : _GEN_2635;
  wire [13:0] _GEN_2637 = 14'ha4d == index ? 14'h14 : _GEN_2636;
  wire [13:0] _GEN_2638 = 14'ha4e == index ? 14'h14 : _GEN_2637;
  wire [13:0] _GEN_2639 = 14'ha4f == index ? 14'h14 : _GEN_2638;
  wire [13:0] _GEN_2640 = 14'ha50 == index ? 14'h14 : _GEN_2639;
  wire [13:0] _GEN_2641 = 14'ha51 == index ? 14'h14 : _GEN_2640;
  wire [13:0] _GEN_2642 = 14'ha52 == index ? 14'h14 : _GEN_2641;
  wire [13:0] _GEN_2643 = 14'ha53 == index ? 14'h14 : _GEN_2642;
  wire [13:0] _GEN_2644 = 14'ha54 == index ? 14'h14 : _GEN_2643;
  wire [13:0] _GEN_2645 = 14'ha55 == index ? 14'h14 : _GEN_2644;
  wire [13:0] _GEN_2646 = 14'ha56 == index ? 14'h14 : _GEN_2645;
  wire [13:0] _GEN_2647 = 14'ha57 == index ? 14'h14 : _GEN_2646;
  wire [13:0] _GEN_2648 = 14'ha58 == index ? 14'h14 : _GEN_2647;
  wire [13:0] _GEN_2649 = 14'ha59 == index ? 14'h14 : _GEN_2648;
  wire [13:0] _GEN_2650 = 14'ha5a == index ? 14'h14 : _GEN_2649;
  wire [13:0] _GEN_2651 = 14'ha5b == index ? 14'h14 : _GEN_2650;
  wire [13:0] _GEN_2652 = 14'ha5c == index ? 14'h14 : _GEN_2651;
  wire [13:0] _GEN_2653 = 14'ha5d == index ? 14'h14 : _GEN_2652;
  wire [13:0] _GEN_2654 = 14'ha5e == index ? 14'h14 : _GEN_2653;
  wire [13:0] _GEN_2655 = 14'ha5f == index ? 14'h14 : _GEN_2654;
  wire [13:0] _GEN_2656 = 14'ha60 == index ? 14'h14 : _GEN_2655;
  wire [13:0] _GEN_2657 = 14'ha61 == index ? 14'h14 : _GEN_2656;
  wire [13:0] _GEN_2658 = 14'ha62 == index ? 14'h14 : _GEN_2657;
  wire [13:0] _GEN_2659 = 14'ha63 == index ? 14'h14 : _GEN_2658;
  wire [13:0] _GEN_2660 = 14'ha64 == index ? 14'h14 : _GEN_2659;
  wire [13:0] _GEN_2661 = 14'ha65 == index ? 14'h14 : _GEN_2660;
  wire [13:0] _GEN_2662 = 14'ha66 == index ? 14'h14 : _GEN_2661;
  wire [13:0] _GEN_2663 = 14'ha67 == index ? 14'h14 : _GEN_2662;
  wire [13:0] _GEN_2664 = 14'ha68 == index ? 14'h14 : _GEN_2663;
  wire [13:0] _GEN_2665 = 14'ha69 == index ? 14'h14 : _GEN_2664;
  wire [13:0] _GEN_2666 = 14'ha6a == index ? 14'h14 : _GEN_2665;
  wire [13:0] _GEN_2667 = 14'ha6b == index ? 14'h14 : _GEN_2666;
  wire [13:0] _GEN_2668 = 14'ha6c == index ? 14'h14 : _GEN_2667;
  wire [13:0] _GEN_2669 = 14'ha6d == index ? 14'h14 : _GEN_2668;
  wire [13:0] _GEN_2670 = 14'ha6e == index ? 14'h14 : _GEN_2669;
  wire [13:0] _GEN_2671 = 14'ha6f == index ? 14'h14 : _GEN_2670;
  wire [13:0] _GEN_2672 = 14'ha70 == index ? 14'h14 : _GEN_2671;
  wire [13:0] _GEN_2673 = 14'ha71 == index ? 14'h14 : _GEN_2672;
  wire [13:0] _GEN_2674 = 14'ha72 == index ? 14'h14 : _GEN_2673;
  wire [13:0] _GEN_2675 = 14'ha73 == index ? 14'h14 : _GEN_2674;
  wire [13:0] _GEN_2676 = 14'ha74 == index ? 14'h14 : _GEN_2675;
  wire [13:0] _GEN_2677 = 14'ha75 == index ? 14'h14 : _GEN_2676;
  wire [13:0] _GEN_2678 = 14'ha76 == index ? 14'h14 : _GEN_2677;
  wire [13:0] _GEN_2679 = 14'ha77 == index ? 14'h14 : _GEN_2678;
  wire [13:0] _GEN_2680 = 14'ha78 == index ? 14'h14 : _GEN_2679;
  wire [13:0] _GEN_2681 = 14'ha79 == index ? 14'h14 : _GEN_2680;
  wire [13:0] _GEN_2682 = 14'ha7a == index ? 14'h14 : _GEN_2681;
  wire [13:0] _GEN_2683 = 14'ha7b == index ? 14'h14 : _GEN_2682;
  wire [13:0] _GEN_2684 = 14'ha7c == index ? 14'h14 : _GEN_2683;
  wire [13:0] _GEN_2685 = 14'ha7d == index ? 14'h14 : _GEN_2684;
  wire [13:0] _GEN_2686 = 14'ha7e == index ? 14'h14 : _GEN_2685;
  wire [13:0] _GEN_2687 = 14'ha7f == index ? 14'h14 : _GEN_2686;
  wire [13:0] _GEN_2688 = 14'ha80 == index ? 14'h0 : _GEN_2687;
  wire [13:0] _GEN_2689 = 14'ha81 == index ? 14'ha80 : _GEN_2688;
  wire [13:0] _GEN_2690 = 14'ha82 == index ? 14'h501 : _GEN_2689;
  wire [13:0] _GEN_2691 = 14'ha83 == index ? 14'h380 : _GEN_2690;
  wire [13:0] _GEN_2692 = 14'ha84 == index ? 14'h281 : _GEN_2691;
  wire [13:0] _GEN_2693 = 14'ha85 == index ? 14'h201 : _GEN_2692;
  wire [13:0] _GEN_2694 = 14'ha86 == index ? 14'h183 : _GEN_2693;
  wire [13:0] _GEN_2695 = 14'ha87 == index ? 14'h180 : _GEN_2694;
  wire [13:0] _GEN_2696 = 14'ha88 == index ? 14'h105 : _GEN_2695;
  wire [13:0] _GEN_2697 = 14'ha89 == index ? 14'h103 : _GEN_2696;
  wire [13:0] _GEN_2698 = 14'ha8a == index ? 14'h101 : _GEN_2697;
  wire [13:0] _GEN_2699 = 14'ha8b == index ? 14'h8a : _GEN_2698;
  wire [13:0] _GEN_2700 = 14'ha8c == index ? 14'h89 : _GEN_2699;
  wire [13:0] _GEN_2701 = 14'ha8d == index ? 14'h88 : _GEN_2700;
  wire [13:0] _GEN_2702 = 14'ha8e == index ? 14'h87 : _GEN_2701;
  wire [13:0] _GEN_2703 = 14'ha8f == index ? 14'h86 : _GEN_2702;
  wire [13:0] _GEN_2704 = 14'ha90 == index ? 14'h85 : _GEN_2703;
  wire [13:0] _GEN_2705 = 14'ha91 == index ? 14'h84 : _GEN_2704;
  wire [13:0] _GEN_2706 = 14'ha92 == index ? 14'h83 : _GEN_2705;
  wire [13:0] _GEN_2707 = 14'ha93 == index ? 14'h82 : _GEN_2706;
  wire [13:0] _GEN_2708 = 14'ha94 == index ? 14'h81 : _GEN_2707;
  wire [13:0] _GEN_2709 = 14'ha95 == index ? 14'h80 : _GEN_2708;
  wire [13:0] _GEN_2710 = 14'ha96 == index ? 14'h15 : _GEN_2709;
  wire [13:0] _GEN_2711 = 14'ha97 == index ? 14'h15 : _GEN_2710;
  wire [13:0] _GEN_2712 = 14'ha98 == index ? 14'h15 : _GEN_2711;
  wire [13:0] _GEN_2713 = 14'ha99 == index ? 14'h15 : _GEN_2712;
  wire [13:0] _GEN_2714 = 14'ha9a == index ? 14'h15 : _GEN_2713;
  wire [13:0] _GEN_2715 = 14'ha9b == index ? 14'h15 : _GEN_2714;
  wire [13:0] _GEN_2716 = 14'ha9c == index ? 14'h15 : _GEN_2715;
  wire [13:0] _GEN_2717 = 14'ha9d == index ? 14'h15 : _GEN_2716;
  wire [13:0] _GEN_2718 = 14'ha9e == index ? 14'h15 : _GEN_2717;
  wire [13:0] _GEN_2719 = 14'ha9f == index ? 14'h15 : _GEN_2718;
  wire [13:0] _GEN_2720 = 14'haa0 == index ? 14'h15 : _GEN_2719;
  wire [13:0] _GEN_2721 = 14'haa1 == index ? 14'h15 : _GEN_2720;
  wire [13:0] _GEN_2722 = 14'haa2 == index ? 14'h15 : _GEN_2721;
  wire [13:0] _GEN_2723 = 14'haa3 == index ? 14'h15 : _GEN_2722;
  wire [13:0] _GEN_2724 = 14'haa4 == index ? 14'h15 : _GEN_2723;
  wire [13:0] _GEN_2725 = 14'haa5 == index ? 14'h15 : _GEN_2724;
  wire [13:0] _GEN_2726 = 14'haa6 == index ? 14'h15 : _GEN_2725;
  wire [13:0] _GEN_2727 = 14'haa7 == index ? 14'h15 : _GEN_2726;
  wire [13:0] _GEN_2728 = 14'haa8 == index ? 14'h15 : _GEN_2727;
  wire [13:0] _GEN_2729 = 14'haa9 == index ? 14'h15 : _GEN_2728;
  wire [13:0] _GEN_2730 = 14'haaa == index ? 14'h15 : _GEN_2729;
  wire [13:0] _GEN_2731 = 14'haab == index ? 14'h15 : _GEN_2730;
  wire [13:0] _GEN_2732 = 14'haac == index ? 14'h15 : _GEN_2731;
  wire [13:0] _GEN_2733 = 14'haad == index ? 14'h15 : _GEN_2732;
  wire [13:0] _GEN_2734 = 14'haae == index ? 14'h15 : _GEN_2733;
  wire [13:0] _GEN_2735 = 14'haaf == index ? 14'h15 : _GEN_2734;
  wire [13:0] _GEN_2736 = 14'hab0 == index ? 14'h15 : _GEN_2735;
  wire [13:0] _GEN_2737 = 14'hab1 == index ? 14'h15 : _GEN_2736;
  wire [13:0] _GEN_2738 = 14'hab2 == index ? 14'h15 : _GEN_2737;
  wire [13:0] _GEN_2739 = 14'hab3 == index ? 14'h15 : _GEN_2738;
  wire [13:0] _GEN_2740 = 14'hab4 == index ? 14'h15 : _GEN_2739;
  wire [13:0] _GEN_2741 = 14'hab5 == index ? 14'h15 : _GEN_2740;
  wire [13:0] _GEN_2742 = 14'hab6 == index ? 14'h15 : _GEN_2741;
  wire [13:0] _GEN_2743 = 14'hab7 == index ? 14'h15 : _GEN_2742;
  wire [13:0] _GEN_2744 = 14'hab8 == index ? 14'h15 : _GEN_2743;
  wire [13:0] _GEN_2745 = 14'hab9 == index ? 14'h15 : _GEN_2744;
  wire [13:0] _GEN_2746 = 14'haba == index ? 14'h15 : _GEN_2745;
  wire [13:0] _GEN_2747 = 14'habb == index ? 14'h15 : _GEN_2746;
  wire [13:0] _GEN_2748 = 14'habc == index ? 14'h15 : _GEN_2747;
  wire [13:0] _GEN_2749 = 14'habd == index ? 14'h15 : _GEN_2748;
  wire [13:0] _GEN_2750 = 14'habe == index ? 14'h15 : _GEN_2749;
  wire [13:0] _GEN_2751 = 14'habf == index ? 14'h15 : _GEN_2750;
  wire [13:0] _GEN_2752 = 14'hac0 == index ? 14'h15 : _GEN_2751;
  wire [13:0] _GEN_2753 = 14'hac1 == index ? 14'h15 : _GEN_2752;
  wire [13:0] _GEN_2754 = 14'hac2 == index ? 14'h15 : _GEN_2753;
  wire [13:0] _GEN_2755 = 14'hac3 == index ? 14'h15 : _GEN_2754;
  wire [13:0] _GEN_2756 = 14'hac4 == index ? 14'h15 : _GEN_2755;
  wire [13:0] _GEN_2757 = 14'hac5 == index ? 14'h15 : _GEN_2756;
  wire [13:0] _GEN_2758 = 14'hac6 == index ? 14'h15 : _GEN_2757;
  wire [13:0] _GEN_2759 = 14'hac7 == index ? 14'h15 : _GEN_2758;
  wire [13:0] _GEN_2760 = 14'hac8 == index ? 14'h15 : _GEN_2759;
  wire [13:0] _GEN_2761 = 14'hac9 == index ? 14'h15 : _GEN_2760;
  wire [13:0] _GEN_2762 = 14'haca == index ? 14'h15 : _GEN_2761;
  wire [13:0] _GEN_2763 = 14'hacb == index ? 14'h15 : _GEN_2762;
  wire [13:0] _GEN_2764 = 14'hacc == index ? 14'h15 : _GEN_2763;
  wire [13:0] _GEN_2765 = 14'hacd == index ? 14'h15 : _GEN_2764;
  wire [13:0] _GEN_2766 = 14'hace == index ? 14'h15 : _GEN_2765;
  wire [13:0] _GEN_2767 = 14'hacf == index ? 14'h15 : _GEN_2766;
  wire [13:0] _GEN_2768 = 14'had0 == index ? 14'h15 : _GEN_2767;
  wire [13:0] _GEN_2769 = 14'had1 == index ? 14'h15 : _GEN_2768;
  wire [13:0] _GEN_2770 = 14'had2 == index ? 14'h15 : _GEN_2769;
  wire [13:0] _GEN_2771 = 14'had3 == index ? 14'h15 : _GEN_2770;
  wire [13:0] _GEN_2772 = 14'had4 == index ? 14'h15 : _GEN_2771;
  wire [13:0] _GEN_2773 = 14'had5 == index ? 14'h15 : _GEN_2772;
  wire [13:0] _GEN_2774 = 14'had6 == index ? 14'h15 : _GEN_2773;
  wire [13:0] _GEN_2775 = 14'had7 == index ? 14'h15 : _GEN_2774;
  wire [13:0] _GEN_2776 = 14'had8 == index ? 14'h15 : _GEN_2775;
  wire [13:0] _GEN_2777 = 14'had9 == index ? 14'h15 : _GEN_2776;
  wire [13:0] _GEN_2778 = 14'hada == index ? 14'h15 : _GEN_2777;
  wire [13:0] _GEN_2779 = 14'hadb == index ? 14'h15 : _GEN_2778;
  wire [13:0] _GEN_2780 = 14'hadc == index ? 14'h15 : _GEN_2779;
  wire [13:0] _GEN_2781 = 14'hadd == index ? 14'h15 : _GEN_2780;
  wire [13:0] _GEN_2782 = 14'hade == index ? 14'h15 : _GEN_2781;
  wire [13:0] _GEN_2783 = 14'hadf == index ? 14'h15 : _GEN_2782;
  wire [13:0] _GEN_2784 = 14'hae0 == index ? 14'h15 : _GEN_2783;
  wire [13:0] _GEN_2785 = 14'hae1 == index ? 14'h15 : _GEN_2784;
  wire [13:0] _GEN_2786 = 14'hae2 == index ? 14'h15 : _GEN_2785;
  wire [13:0] _GEN_2787 = 14'hae3 == index ? 14'h15 : _GEN_2786;
  wire [13:0] _GEN_2788 = 14'hae4 == index ? 14'h15 : _GEN_2787;
  wire [13:0] _GEN_2789 = 14'hae5 == index ? 14'h15 : _GEN_2788;
  wire [13:0] _GEN_2790 = 14'hae6 == index ? 14'h15 : _GEN_2789;
  wire [13:0] _GEN_2791 = 14'hae7 == index ? 14'h15 : _GEN_2790;
  wire [13:0] _GEN_2792 = 14'hae8 == index ? 14'h15 : _GEN_2791;
  wire [13:0] _GEN_2793 = 14'hae9 == index ? 14'h15 : _GEN_2792;
  wire [13:0] _GEN_2794 = 14'haea == index ? 14'h15 : _GEN_2793;
  wire [13:0] _GEN_2795 = 14'haeb == index ? 14'h15 : _GEN_2794;
  wire [13:0] _GEN_2796 = 14'haec == index ? 14'h15 : _GEN_2795;
  wire [13:0] _GEN_2797 = 14'haed == index ? 14'h15 : _GEN_2796;
  wire [13:0] _GEN_2798 = 14'haee == index ? 14'h15 : _GEN_2797;
  wire [13:0] _GEN_2799 = 14'haef == index ? 14'h15 : _GEN_2798;
  wire [13:0] _GEN_2800 = 14'haf0 == index ? 14'h15 : _GEN_2799;
  wire [13:0] _GEN_2801 = 14'haf1 == index ? 14'h15 : _GEN_2800;
  wire [13:0] _GEN_2802 = 14'haf2 == index ? 14'h15 : _GEN_2801;
  wire [13:0] _GEN_2803 = 14'haf3 == index ? 14'h15 : _GEN_2802;
  wire [13:0] _GEN_2804 = 14'haf4 == index ? 14'h15 : _GEN_2803;
  wire [13:0] _GEN_2805 = 14'haf5 == index ? 14'h15 : _GEN_2804;
  wire [13:0] _GEN_2806 = 14'haf6 == index ? 14'h15 : _GEN_2805;
  wire [13:0] _GEN_2807 = 14'haf7 == index ? 14'h15 : _GEN_2806;
  wire [13:0] _GEN_2808 = 14'haf8 == index ? 14'h15 : _GEN_2807;
  wire [13:0] _GEN_2809 = 14'haf9 == index ? 14'h15 : _GEN_2808;
  wire [13:0] _GEN_2810 = 14'hafa == index ? 14'h15 : _GEN_2809;
  wire [13:0] _GEN_2811 = 14'hafb == index ? 14'h15 : _GEN_2810;
  wire [13:0] _GEN_2812 = 14'hafc == index ? 14'h15 : _GEN_2811;
  wire [13:0] _GEN_2813 = 14'hafd == index ? 14'h15 : _GEN_2812;
  wire [13:0] _GEN_2814 = 14'hafe == index ? 14'h15 : _GEN_2813;
  wire [13:0] _GEN_2815 = 14'haff == index ? 14'h15 : _GEN_2814;
  wire [13:0] _GEN_2816 = 14'hb00 == index ? 14'h0 : _GEN_2815;
  wire [13:0] _GEN_2817 = 14'hb01 == index ? 14'hb00 : _GEN_2816;
  wire [13:0] _GEN_2818 = 14'hb02 == index ? 14'h580 : _GEN_2817;
  wire [13:0] _GEN_2819 = 14'hb03 == index ? 14'h381 : _GEN_2818;
  wire [13:0] _GEN_2820 = 14'hb04 == index ? 14'h282 : _GEN_2819;
  wire [13:0] _GEN_2821 = 14'hb05 == index ? 14'h202 : _GEN_2820;
  wire [13:0] _GEN_2822 = 14'hb06 == index ? 14'h184 : _GEN_2821;
  wire [13:0] _GEN_2823 = 14'hb07 == index ? 14'h181 : _GEN_2822;
  wire [13:0] _GEN_2824 = 14'hb08 == index ? 14'h106 : _GEN_2823;
  wire [13:0] _GEN_2825 = 14'hb09 == index ? 14'h104 : _GEN_2824;
  wire [13:0] _GEN_2826 = 14'hb0a == index ? 14'h102 : _GEN_2825;
  wire [13:0] _GEN_2827 = 14'hb0b == index ? 14'h100 : _GEN_2826;
  wire [13:0] _GEN_2828 = 14'hb0c == index ? 14'h8a : _GEN_2827;
  wire [13:0] _GEN_2829 = 14'hb0d == index ? 14'h89 : _GEN_2828;
  wire [13:0] _GEN_2830 = 14'hb0e == index ? 14'h88 : _GEN_2829;
  wire [13:0] _GEN_2831 = 14'hb0f == index ? 14'h87 : _GEN_2830;
  wire [13:0] _GEN_2832 = 14'hb10 == index ? 14'h86 : _GEN_2831;
  wire [13:0] _GEN_2833 = 14'hb11 == index ? 14'h85 : _GEN_2832;
  wire [13:0] _GEN_2834 = 14'hb12 == index ? 14'h84 : _GEN_2833;
  wire [13:0] _GEN_2835 = 14'hb13 == index ? 14'h83 : _GEN_2834;
  wire [13:0] _GEN_2836 = 14'hb14 == index ? 14'h82 : _GEN_2835;
  wire [13:0] _GEN_2837 = 14'hb15 == index ? 14'h81 : _GEN_2836;
  wire [13:0] _GEN_2838 = 14'hb16 == index ? 14'h80 : _GEN_2837;
  wire [13:0] _GEN_2839 = 14'hb17 == index ? 14'h16 : _GEN_2838;
  wire [13:0] _GEN_2840 = 14'hb18 == index ? 14'h16 : _GEN_2839;
  wire [13:0] _GEN_2841 = 14'hb19 == index ? 14'h16 : _GEN_2840;
  wire [13:0] _GEN_2842 = 14'hb1a == index ? 14'h16 : _GEN_2841;
  wire [13:0] _GEN_2843 = 14'hb1b == index ? 14'h16 : _GEN_2842;
  wire [13:0] _GEN_2844 = 14'hb1c == index ? 14'h16 : _GEN_2843;
  wire [13:0] _GEN_2845 = 14'hb1d == index ? 14'h16 : _GEN_2844;
  wire [13:0] _GEN_2846 = 14'hb1e == index ? 14'h16 : _GEN_2845;
  wire [13:0] _GEN_2847 = 14'hb1f == index ? 14'h16 : _GEN_2846;
  wire [13:0] _GEN_2848 = 14'hb20 == index ? 14'h16 : _GEN_2847;
  wire [13:0] _GEN_2849 = 14'hb21 == index ? 14'h16 : _GEN_2848;
  wire [13:0] _GEN_2850 = 14'hb22 == index ? 14'h16 : _GEN_2849;
  wire [13:0] _GEN_2851 = 14'hb23 == index ? 14'h16 : _GEN_2850;
  wire [13:0] _GEN_2852 = 14'hb24 == index ? 14'h16 : _GEN_2851;
  wire [13:0] _GEN_2853 = 14'hb25 == index ? 14'h16 : _GEN_2852;
  wire [13:0] _GEN_2854 = 14'hb26 == index ? 14'h16 : _GEN_2853;
  wire [13:0] _GEN_2855 = 14'hb27 == index ? 14'h16 : _GEN_2854;
  wire [13:0] _GEN_2856 = 14'hb28 == index ? 14'h16 : _GEN_2855;
  wire [13:0] _GEN_2857 = 14'hb29 == index ? 14'h16 : _GEN_2856;
  wire [13:0] _GEN_2858 = 14'hb2a == index ? 14'h16 : _GEN_2857;
  wire [13:0] _GEN_2859 = 14'hb2b == index ? 14'h16 : _GEN_2858;
  wire [13:0] _GEN_2860 = 14'hb2c == index ? 14'h16 : _GEN_2859;
  wire [13:0] _GEN_2861 = 14'hb2d == index ? 14'h16 : _GEN_2860;
  wire [13:0] _GEN_2862 = 14'hb2e == index ? 14'h16 : _GEN_2861;
  wire [13:0] _GEN_2863 = 14'hb2f == index ? 14'h16 : _GEN_2862;
  wire [13:0] _GEN_2864 = 14'hb30 == index ? 14'h16 : _GEN_2863;
  wire [13:0] _GEN_2865 = 14'hb31 == index ? 14'h16 : _GEN_2864;
  wire [13:0] _GEN_2866 = 14'hb32 == index ? 14'h16 : _GEN_2865;
  wire [13:0] _GEN_2867 = 14'hb33 == index ? 14'h16 : _GEN_2866;
  wire [13:0] _GEN_2868 = 14'hb34 == index ? 14'h16 : _GEN_2867;
  wire [13:0] _GEN_2869 = 14'hb35 == index ? 14'h16 : _GEN_2868;
  wire [13:0] _GEN_2870 = 14'hb36 == index ? 14'h16 : _GEN_2869;
  wire [13:0] _GEN_2871 = 14'hb37 == index ? 14'h16 : _GEN_2870;
  wire [13:0] _GEN_2872 = 14'hb38 == index ? 14'h16 : _GEN_2871;
  wire [13:0] _GEN_2873 = 14'hb39 == index ? 14'h16 : _GEN_2872;
  wire [13:0] _GEN_2874 = 14'hb3a == index ? 14'h16 : _GEN_2873;
  wire [13:0] _GEN_2875 = 14'hb3b == index ? 14'h16 : _GEN_2874;
  wire [13:0] _GEN_2876 = 14'hb3c == index ? 14'h16 : _GEN_2875;
  wire [13:0] _GEN_2877 = 14'hb3d == index ? 14'h16 : _GEN_2876;
  wire [13:0] _GEN_2878 = 14'hb3e == index ? 14'h16 : _GEN_2877;
  wire [13:0] _GEN_2879 = 14'hb3f == index ? 14'h16 : _GEN_2878;
  wire [13:0] _GEN_2880 = 14'hb40 == index ? 14'h16 : _GEN_2879;
  wire [13:0] _GEN_2881 = 14'hb41 == index ? 14'h16 : _GEN_2880;
  wire [13:0] _GEN_2882 = 14'hb42 == index ? 14'h16 : _GEN_2881;
  wire [13:0] _GEN_2883 = 14'hb43 == index ? 14'h16 : _GEN_2882;
  wire [13:0] _GEN_2884 = 14'hb44 == index ? 14'h16 : _GEN_2883;
  wire [13:0] _GEN_2885 = 14'hb45 == index ? 14'h16 : _GEN_2884;
  wire [13:0] _GEN_2886 = 14'hb46 == index ? 14'h16 : _GEN_2885;
  wire [13:0] _GEN_2887 = 14'hb47 == index ? 14'h16 : _GEN_2886;
  wire [13:0] _GEN_2888 = 14'hb48 == index ? 14'h16 : _GEN_2887;
  wire [13:0] _GEN_2889 = 14'hb49 == index ? 14'h16 : _GEN_2888;
  wire [13:0] _GEN_2890 = 14'hb4a == index ? 14'h16 : _GEN_2889;
  wire [13:0] _GEN_2891 = 14'hb4b == index ? 14'h16 : _GEN_2890;
  wire [13:0] _GEN_2892 = 14'hb4c == index ? 14'h16 : _GEN_2891;
  wire [13:0] _GEN_2893 = 14'hb4d == index ? 14'h16 : _GEN_2892;
  wire [13:0] _GEN_2894 = 14'hb4e == index ? 14'h16 : _GEN_2893;
  wire [13:0] _GEN_2895 = 14'hb4f == index ? 14'h16 : _GEN_2894;
  wire [13:0] _GEN_2896 = 14'hb50 == index ? 14'h16 : _GEN_2895;
  wire [13:0] _GEN_2897 = 14'hb51 == index ? 14'h16 : _GEN_2896;
  wire [13:0] _GEN_2898 = 14'hb52 == index ? 14'h16 : _GEN_2897;
  wire [13:0] _GEN_2899 = 14'hb53 == index ? 14'h16 : _GEN_2898;
  wire [13:0] _GEN_2900 = 14'hb54 == index ? 14'h16 : _GEN_2899;
  wire [13:0] _GEN_2901 = 14'hb55 == index ? 14'h16 : _GEN_2900;
  wire [13:0] _GEN_2902 = 14'hb56 == index ? 14'h16 : _GEN_2901;
  wire [13:0] _GEN_2903 = 14'hb57 == index ? 14'h16 : _GEN_2902;
  wire [13:0] _GEN_2904 = 14'hb58 == index ? 14'h16 : _GEN_2903;
  wire [13:0] _GEN_2905 = 14'hb59 == index ? 14'h16 : _GEN_2904;
  wire [13:0] _GEN_2906 = 14'hb5a == index ? 14'h16 : _GEN_2905;
  wire [13:0] _GEN_2907 = 14'hb5b == index ? 14'h16 : _GEN_2906;
  wire [13:0] _GEN_2908 = 14'hb5c == index ? 14'h16 : _GEN_2907;
  wire [13:0] _GEN_2909 = 14'hb5d == index ? 14'h16 : _GEN_2908;
  wire [13:0] _GEN_2910 = 14'hb5e == index ? 14'h16 : _GEN_2909;
  wire [13:0] _GEN_2911 = 14'hb5f == index ? 14'h16 : _GEN_2910;
  wire [13:0] _GEN_2912 = 14'hb60 == index ? 14'h16 : _GEN_2911;
  wire [13:0] _GEN_2913 = 14'hb61 == index ? 14'h16 : _GEN_2912;
  wire [13:0] _GEN_2914 = 14'hb62 == index ? 14'h16 : _GEN_2913;
  wire [13:0] _GEN_2915 = 14'hb63 == index ? 14'h16 : _GEN_2914;
  wire [13:0] _GEN_2916 = 14'hb64 == index ? 14'h16 : _GEN_2915;
  wire [13:0] _GEN_2917 = 14'hb65 == index ? 14'h16 : _GEN_2916;
  wire [13:0] _GEN_2918 = 14'hb66 == index ? 14'h16 : _GEN_2917;
  wire [13:0] _GEN_2919 = 14'hb67 == index ? 14'h16 : _GEN_2918;
  wire [13:0] _GEN_2920 = 14'hb68 == index ? 14'h16 : _GEN_2919;
  wire [13:0] _GEN_2921 = 14'hb69 == index ? 14'h16 : _GEN_2920;
  wire [13:0] _GEN_2922 = 14'hb6a == index ? 14'h16 : _GEN_2921;
  wire [13:0] _GEN_2923 = 14'hb6b == index ? 14'h16 : _GEN_2922;
  wire [13:0] _GEN_2924 = 14'hb6c == index ? 14'h16 : _GEN_2923;
  wire [13:0] _GEN_2925 = 14'hb6d == index ? 14'h16 : _GEN_2924;
  wire [13:0] _GEN_2926 = 14'hb6e == index ? 14'h16 : _GEN_2925;
  wire [13:0] _GEN_2927 = 14'hb6f == index ? 14'h16 : _GEN_2926;
  wire [13:0] _GEN_2928 = 14'hb70 == index ? 14'h16 : _GEN_2927;
  wire [13:0] _GEN_2929 = 14'hb71 == index ? 14'h16 : _GEN_2928;
  wire [13:0] _GEN_2930 = 14'hb72 == index ? 14'h16 : _GEN_2929;
  wire [13:0] _GEN_2931 = 14'hb73 == index ? 14'h16 : _GEN_2930;
  wire [13:0] _GEN_2932 = 14'hb74 == index ? 14'h16 : _GEN_2931;
  wire [13:0] _GEN_2933 = 14'hb75 == index ? 14'h16 : _GEN_2932;
  wire [13:0] _GEN_2934 = 14'hb76 == index ? 14'h16 : _GEN_2933;
  wire [13:0] _GEN_2935 = 14'hb77 == index ? 14'h16 : _GEN_2934;
  wire [13:0] _GEN_2936 = 14'hb78 == index ? 14'h16 : _GEN_2935;
  wire [13:0] _GEN_2937 = 14'hb79 == index ? 14'h16 : _GEN_2936;
  wire [13:0] _GEN_2938 = 14'hb7a == index ? 14'h16 : _GEN_2937;
  wire [13:0] _GEN_2939 = 14'hb7b == index ? 14'h16 : _GEN_2938;
  wire [13:0] _GEN_2940 = 14'hb7c == index ? 14'h16 : _GEN_2939;
  wire [13:0] _GEN_2941 = 14'hb7d == index ? 14'h16 : _GEN_2940;
  wire [13:0] _GEN_2942 = 14'hb7e == index ? 14'h16 : _GEN_2941;
  wire [13:0] _GEN_2943 = 14'hb7f == index ? 14'h16 : _GEN_2942;
  wire [13:0] _GEN_2944 = 14'hb80 == index ? 14'h0 : _GEN_2943;
  wire [13:0] _GEN_2945 = 14'hb81 == index ? 14'hb80 : _GEN_2944;
  wire [13:0] _GEN_2946 = 14'hb82 == index ? 14'h581 : _GEN_2945;
  wire [13:0] _GEN_2947 = 14'hb83 == index ? 14'h382 : _GEN_2946;
  wire [13:0] _GEN_2948 = 14'hb84 == index ? 14'h283 : _GEN_2947;
  wire [13:0] _GEN_2949 = 14'hb85 == index ? 14'h203 : _GEN_2948;
  wire [13:0] _GEN_2950 = 14'hb86 == index ? 14'h185 : _GEN_2949;
  wire [13:0] _GEN_2951 = 14'hb87 == index ? 14'h182 : _GEN_2950;
  wire [13:0] _GEN_2952 = 14'hb88 == index ? 14'h107 : _GEN_2951;
  wire [13:0] _GEN_2953 = 14'hb89 == index ? 14'h105 : _GEN_2952;
  wire [13:0] _GEN_2954 = 14'hb8a == index ? 14'h103 : _GEN_2953;
  wire [13:0] _GEN_2955 = 14'hb8b == index ? 14'h101 : _GEN_2954;
  wire [13:0] _GEN_2956 = 14'hb8c == index ? 14'h8b : _GEN_2955;
  wire [13:0] _GEN_2957 = 14'hb8d == index ? 14'h8a : _GEN_2956;
  wire [13:0] _GEN_2958 = 14'hb8e == index ? 14'h89 : _GEN_2957;
  wire [13:0] _GEN_2959 = 14'hb8f == index ? 14'h88 : _GEN_2958;
  wire [13:0] _GEN_2960 = 14'hb90 == index ? 14'h87 : _GEN_2959;
  wire [13:0] _GEN_2961 = 14'hb91 == index ? 14'h86 : _GEN_2960;
  wire [13:0] _GEN_2962 = 14'hb92 == index ? 14'h85 : _GEN_2961;
  wire [13:0] _GEN_2963 = 14'hb93 == index ? 14'h84 : _GEN_2962;
  wire [13:0] _GEN_2964 = 14'hb94 == index ? 14'h83 : _GEN_2963;
  wire [13:0] _GEN_2965 = 14'hb95 == index ? 14'h82 : _GEN_2964;
  wire [13:0] _GEN_2966 = 14'hb96 == index ? 14'h81 : _GEN_2965;
  wire [13:0] _GEN_2967 = 14'hb97 == index ? 14'h80 : _GEN_2966;
  wire [13:0] _GEN_2968 = 14'hb98 == index ? 14'h17 : _GEN_2967;
  wire [13:0] _GEN_2969 = 14'hb99 == index ? 14'h17 : _GEN_2968;
  wire [13:0] _GEN_2970 = 14'hb9a == index ? 14'h17 : _GEN_2969;
  wire [13:0] _GEN_2971 = 14'hb9b == index ? 14'h17 : _GEN_2970;
  wire [13:0] _GEN_2972 = 14'hb9c == index ? 14'h17 : _GEN_2971;
  wire [13:0] _GEN_2973 = 14'hb9d == index ? 14'h17 : _GEN_2972;
  wire [13:0] _GEN_2974 = 14'hb9e == index ? 14'h17 : _GEN_2973;
  wire [13:0] _GEN_2975 = 14'hb9f == index ? 14'h17 : _GEN_2974;
  wire [13:0] _GEN_2976 = 14'hba0 == index ? 14'h17 : _GEN_2975;
  wire [13:0] _GEN_2977 = 14'hba1 == index ? 14'h17 : _GEN_2976;
  wire [13:0] _GEN_2978 = 14'hba2 == index ? 14'h17 : _GEN_2977;
  wire [13:0] _GEN_2979 = 14'hba3 == index ? 14'h17 : _GEN_2978;
  wire [13:0] _GEN_2980 = 14'hba4 == index ? 14'h17 : _GEN_2979;
  wire [13:0] _GEN_2981 = 14'hba5 == index ? 14'h17 : _GEN_2980;
  wire [13:0] _GEN_2982 = 14'hba6 == index ? 14'h17 : _GEN_2981;
  wire [13:0] _GEN_2983 = 14'hba7 == index ? 14'h17 : _GEN_2982;
  wire [13:0] _GEN_2984 = 14'hba8 == index ? 14'h17 : _GEN_2983;
  wire [13:0] _GEN_2985 = 14'hba9 == index ? 14'h17 : _GEN_2984;
  wire [13:0] _GEN_2986 = 14'hbaa == index ? 14'h17 : _GEN_2985;
  wire [13:0] _GEN_2987 = 14'hbab == index ? 14'h17 : _GEN_2986;
  wire [13:0] _GEN_2988 = 14'hbac == index ? 14'h17 : _GEN_2987;
  wire [13:0] _GEN_2989 = 14'hbad == index ? 14'h17 : _GEN_2988;
  wire [13:0] _GEN_2990 = 14'hbae == index ? 14'h17 : _GEN_2989;
  wire [13:0] _GEN_2991 = 14'hbaf == index ? 14'h17 : _GEN_2990;
  wire [13:0] _GEN_2992 = 14'hbb0 == index ? 14'h17 : _GEN_2991;
  wire [13:0] _GEN_2993 = 14'hbb1 == index ? 14'h17 : _GEN_2992;
  wire [13:0] _GEN_2994 = 14'hbb2 == index ? 14'h17 : _GEN_2993;
  wire [13:0] _GEN_2995 = 14'hbb3 == index ? 14'h17 : _GEN_2994;
  wire [13:0] _GEN_2996 = 14'hbb4 == index ? 14'h17 : _GEN_2995;
  wire [13:0] _GEN_2997 = 14'hbb5 == index ? 14'h17 : _GEN_2996;
  wire [13:0] _GEN_2998 = 14'hbb6 == index ? 14'h17 : _GEN_2997;
  wire [13:0] _GEN_2999 = 14'hbb7 == index ? 14'h17 : _GEN_2998;
  wire [13:0] _GEN_3000 = 14'hbb8 == index ? 14'h17 : _GEN_2999;
  wire [13:0] _GEN_3001 = 14'hbb9 == index ? 14'h17 : _GEN_3000;
  wire [13:0] _GEN_3002 = 14'hbba == index ? 14'h17 : _GEN_3001;
  wire [13:0] _GEN_3003 = 14'hbbb == index ? 14'h17 : _GEN_3002;
  wire [13:0] _GEN_3004 = 14'hbbc == index ? 14'h17 : _GEN_3003;
  wire [13:0] _GEN_3005 = 14'hbbd == index ? 14'h17 : _GEN_3004;
  wire [13:0] _GEN_3006 = 14'hbbe == index ? 14'h17 : _GEN_3005;
  wire [13:0] _GEN_3007 = 14'hbbf == index ? 14'h17 : _GEN_3006;
  wire [13:0] _GEN_3008 = 14'hbc0 == index ? 14'h17 : _GEN_3007;
  wire [13:0] _GEN_3009 = 14'hbc1 == index ? 14'h17 : _GEN_3008;
  wire [13:0] _GEN_3010 = 14'hbc2 == index ? 14'h17 : _GEN_3009;
  wire [13:0] _GEN_3011 = 14'hbc3 == index ? 14'h17 : _GEN_3010;
  wire [13:0] _GEN_3012 = 14'hbc4 == index ? 14'h17 : _GEN_3011;
  wire [13:0] _GEN_3013 = 14'hbc5 == index ? 14'h17 : _GEN_3012;
  wire [13:0] _GEN_3014 = 14'hbc6 == index ? 14'h17 : _GEN_3013;
  wire [13:0] _GEN_3015 = 14'hbc7 == index ? 14'h17 : _GEN_3014;
  wire [13:0] _GEN_3016 = 14'hbc8 == index ? 14'h17 : _GEN_3015;
  wire [13:0] _GEN_3017 = 14'hbc9 == index ? 14'h17 : _GEN_3016;
  wire [13:0] _GEN_3018 = 14'hbca == index ? 14'h17 : _GEN_3017;
  wire [13:0] _GEN_3019 = 14'hbcb == index ? 14'h17 : _GEN_3018;
  wire [13:0] _GEN_3020 = 14'hbcc == index ? 14'h17 : _GEN_3019;
  wire [13:0] _GEN_3021 = 14'hbcd == index ? 14'h17 : _GEN_3020;
  wire [13:0] _GEN_3022 = 14'hbce == index ? 14'h17 : _GEN_3021;
  wire [13:0] _GEN_3023 = 14'hbcf == index ? 14'h17 : _GEN_3022;
  wire [13:0] _GEN_3024 = 14'hbd0 == index ? 14'h17 : _GEN_3023;
  wire [13:0] _GEN_3025 = 14'hbd1 == index ? 14'h17 : _GEN_3024;
  wire [13:0] _GEN_3026 = 14'hbd2 == index ? 14'h17 : _GEN_3025;
  wire [13:0] _GEN_3027 = 14'hbd3 == index ? 14'h17 : _GEN_3026;
  wire [13:0] _GEN_3028 = 14'hbd4 == index ? 14'h17 : _GEN_3027;
  wire [13:0] _GEN_3029 = 14'hbd5 == index ? 14'h17 : _GEN_3028;
  wire [13:0] _GEN_3030 = 14'hbd6 == index ? 14'h17 : _GEN_3029;
  wire [13:0] _GEN_3031 = 14'hbd7 == index ? 14'h17 : _GEN_3030;
  wire [13:0] _GEN_3032 = 14'hbd8 == index ? 14'h17 : _GEN_3031;
  wire [13:0] _GEN_3033 = 14'hbd9 == index ? 14'h17 : _GEN_3032;
  wire [13:0] _GEN_3034 = 14'hbda == index ? 14'h17 : _GEN_3033;
  wire [13:0] _GEN_3035 = 14'hbdb == index ? 14'h17 : _GEN_3034;
  wire [13:0] _GEN_3036 = 14'hbdc == index ? 14'h17 : _GEN_3035;
  wire [13:0] _GEN_3037 = 14'hbdd == index ? 14'h17 : _GEN_3036;
  wire [13:0] _GEN_3038 = 14'hbde == index ? 14'h17 : _GEN_3037;
  wire [13:0] _GEN_3039 = 14'hbdf == index ? 14'h17 : _GEN_3038;
  wire [13:0] _GEN_3040 = 14'hbe0 == index ? 14'h17 : _GEN_3039;
  wire [13:0] _GEN_3041 = 14'hbe1 == index ? 14'h17 : _GEN_3040;
  wire [13:0] _GEN_3042 = 14'hbe2 == index ? 14'h17 : _GEN_3041;
  wire [13:0] _GEN_3043 = 14'hbe3 == index ? 14'h17 : _GEN_3042;
  wire [13:0] _GEN_3044 = 14'hbe4 == index ? 14'h17 : _GEN_3043;
  wire [13:0] _GEN_3045 = 14'hbe5 == index ? 14'h17 : _GEN_3044;
  wire [13:0] _GEN_3046 = 14'hbe6 == index ? 14'h17 : _GEN_3045;
  wire [13:0] _GEN_3047 = 14'hbe7 == index ? 14'h17 : _GEN_3046;
  wire [13:0] _GEN_3048 = 14'hbe8 == index ? 14'h17 : _GEN_3047;
  wire [13:0] _GEN_3049 = 14'hbe9 == index ? 14'h17 : _GEN_3048;
  wire [13:0] _GEN_3050 = 14'hbea == index ? 14'h17 : _GEN_3049;
  wire [13:0] _GEN_3051 = 14'hbeb == index ? 14'h17 : _GEN_3050;
  wire [13:0] _GEN_3052 = 14'hbec == index ? 14'h17 : _GEN_3051;
  wire [13:0] _GEN_3053 = 14'hbed == index ? 14'h17 : _GEN_3052;
  wire [13:0] _GEN_3054 = 14'hbee == index ? 14'h17 : _GEN_3053;
  wire [13:0] _GEN_3055 = 14'hbef == index ? 14'h17 : _GEN_3054;
  wire [13:0] _GEN_3056 = 14'hbf0 == index ? 14'h17 : _GEN_3055;
  wire [13:0] _GEN_3057 = 14'hbf1 == index ? 14'h17 : _GEN_3056;
  wire [13:0] _GEN_3058 = 14'hbf2 == index ? 14'h17 : _GEN_3057;
  wire [13:0] _GEN_3059 = 14'hbf3 == index ? 14'h17 : _GEN_3058;
  wire [13:0] _GEN_3060 = 14'hbf4 == index ? 14'h17 : _GEN_3059;
  wire [13:0] _GEN_3061 = 14'hbf5 == index ? 14'h17 : _GEN_3060;
  wire [13:0] _GEN_3062 = 14'hbf6 == index ? 14'h17 : _GEN_3061;
  wire [13:0] _GEN_3063 = 14'hbf7 == index ? 14'h17 : _GEN_3062;
  wire [13:0] _GEN_3064 = 14'hbf8 == index ? 14'h17 : _GEN_3063;
  wire [13:0] _GEN_3065 = 14'hbf9 == index ? 14'h17 : _GEN_3064;
  wire [13:0] _GEN_3066 = 14'hbfa == index ? 14'h17 : _GEN_3065;
  wire [13:0] _GEN_3067 = 14'hbfb == index ? 14'h17 : _GEN_3066;
  wire [13:0] _GEN_3068 = 14'hbfc == index ? 14'h17 : _GEN_3067;
  wire [13:0] _GEN_3069 = 14'hbfd == index ? 14'h17 : _GEN_3068;
  wire [13:0] _GEN_3070 = 14'hbfe == index ? 14'h17 : _GEN_3069;
  wire [13:0] _GEN_3071 = 14'hbff == index ? 14'h17 : _GEN_3070;
  wire [13:0] _GEN_3072 = 14'hc00 == index ? 14'h0 : _GEN_3071;
  wire [13:0] _GEN_3073 = 14'hc01 == index ? 14'hc00 : _GEN_3072;
  wire [13:0] _GEN_3074 = 14'hc02 == index ? 14'h600 : _GEN_3073;
  wire [13:0] _GEN_3075 = 14'hc03 == index ? 14'h400 : _GEN_3074;
  wire [13:0] _GEN_3076 = 14'hc04 == index ? 14'h300 : _GEN_3075;
  wire [13:0] _GEN_3077 = 14'hc05 == index ? 14'h204 : _GEN_3076;
  wire [13:0] _GEN_3078 = 14'hc06 == index ? 14'h200 : _GEN_3077;
  wire [13:0] _GEN_3079 = 14'hc07 == index ? 14'h183 : _GEN_3078;
  wire [13:0] _GEN_3080 = 14'hc08 == index ? 14'h180 : _GEN_3079;
  wire [13:0] _GEN_3081 = 14'hc09 == index ? 14'h106 : _GEN_3080;
  wire [13:0] _GEN_3082 = 14'hc0a == index ? 14'h104 : _GEN_3081;
  wire [13:0] _GEN_3083 = 14'hc0b == index ? 14'h102 : _GEN_3082;
  wire [13:0] _GEN_3084 = 14'hc0c == index ? 14'h100 : _GEN_3083;
  wire [13:0] _GEN_3085 = 14'hc0d == index ? 14'h8b : _GEN_3084;
  wire [13:0] _GEN_3086 = 14'hc0e == index ? 14'h8a : _GEN_3085;
  wire [13:0] _GEN_3087 = 14'hc0f == index ? 14'h89 : _GEN_3086;
  wire [13:0] _GEN_3088 = 14'hc10 == index ? 14'h88 : _GEN_3087;
  wire [13:0] _GEN_3089 = 14'hc11 == index ? 14'h87 : _GEN_3088;
  wire [13:0] _GEN_3090 = 14'hc12 == index ? 14'h86 : _GEN_3089;
  wire [13:0] _GEN_3091 = 14'hc13 == index ? 14'h85 : _GEN_3090;
  wire [13:0] _GEN_3092 = 14'hc14 == index ? 14'h84 : _GEN_3091;
  wire [13:0] _GEN_3093 = 14'hc15 == index ? 14'h83 : _GEN_3092;
  wire [13:0] _GEN_3094 = 14'hc16 == index ? 14'h82 : _GEN_3093;
  wire [13:0] _GEN_3095 = 14'hc17 == index ? 14'h81 : _GEN_3094;
  wire [13:0] _GEN_3096 = 14'hc18 == index ? 14'h80 : _GEN_3095;
  wire [13:0] _GEN_3097 = 14'hc19 == index ? 14'h18 : _GEN_3096;
  wire [13:0] _GEN_3098 = 14'hc1a == index ? 14'h18 : _GEN_3097;
  wire [13:0] _GEN_3099 = 14'hc1b == index ? 14'h18 : _GEN_3098;
  wire [13:0] _GEN_3100 = 14'hc1c == index ? 14'h18 : _GEN_3099;
  wire [13:0] _GEN_3101 = 14'hc1d == index ? 14'h18 : _GEN_3100;
  wire [13:0] _GEN_3102 = 14'hc1e == index ? 14'h18 : _GEN_3101;
  wire [13:0] _GEN_3103 = 14'hc1f == index ? 14'h18 : _GEN_3102;
  wire [13:0] _GEN_3104 = 14'hc20 == index ? 14'h18 : _GEN_3103;
  wire [13:0] _GEN_3105 = 14'hc21 == index ? 14'h18 : _GEN_3104;
  wire [13:0] _GEN_3106 = 14'hc22 == index ? 14'h18 : _GEN_3105;
  wire [13:0] _GEN_3107 = 14'hc23 == index ? 14'h18 : _GEN_3106;
  wire [13:0] _GEN_3108 = 14'hc24 == index ? 14'h18 : _GEN_3107;
  wire [13:0] _GEN_3109 = 14'hc25 == index ? 14'h18 : _GEN_3108;
  wire [13:0] _GEN_3110 = 14'hc26 == index ? 14'h18 : _GEN_3109;
  wire [13:0] _GEN_3111 = 14'hc27 == index ? 14'h18 : _GEN_3110;
  wire [13:0] _GEN_3112 = 14'hc28 == index ? 14'h18 : _GEN_3111;
  wire [13:0] _GEN_3113 = 14'hc29 == index ? 14'h18 : _GEN_3112;
  wire [13:0] _GEN_3114 = 14'hc2a == index ? 14'h18 : _GEN_3113;
  wire [13:0] _GEN_3115 = 14'hc2b == index ? 14'h18 : _GEN_3114;
  wire [13:0] _GEN_3116 = 14'hc2c == index ? 14'h18 : _GEN_3115;
  wire [13:0] _GEN_3117 = 14'hc2d == index ? 14'h18 : _GEN_3116;
  wire [13:0] _GEN_3118 = 14'hc2e == index ? 14'h18 : _GEN_3117;
  wire [13:0] _GEN_3119 = 14'hc2f == index ? 14'h18 : _GEN_3118;
  wire [13:0] _GEN_3120 = 14'hc30 == index ? 14'h18 : _GEN_3119;
  wire [13:0] _GEN_3121 = 14'hc31 == index ? 14'h18 : _GEN_3120;
  wire [13:0] _GEN_3122 = 14'hc32 == index ? 14'h18 : _GEN_3121;
  wire [13:0] _GEN_3123 = 14'hc33 == index ? 14'h18 : _GEN_3122;
  wire [13:0] _GEN_3124 = 14'hc34 == index ? 14'h18 : _GEN_3123;
  wire [13:0] _GEN_3125 = 14'hc35 == index ? 14'h18 : _GEN_3124;
  wire [13:0] _GEN_3126 = 14'hc36 == index ? 14'h18 : _GEN_3125;
  wire [13:0] _GEN_3127 = 14'hc37 == index ? 14'h18 : _GEN_3126;
  wire [13:0] _GEN_3128 = 14'hc38 == index ? 14'h18 : _GEN_3127;
  wire [13:0] _GEN_3129 = 14'hc39 == index ? 14'h18 : _GEN_3128;
  wire [13:0] _GEN_3130 = 14'hc3a == index ? 14'h18 : _GEN_3129;
  wire [13:0] _GEN_3131 = 14'hc3b == index ? 14'h18 : _GEN_3130;
  wire [13:0] _GEN_3132 = 14'hc3c == index ? 14'h18 : _GEN_3131;
  wire [13:0] _GEN_3133 = 14'hc3d == index ? 14'h18 : _GEN_3132;
  wire [13:0] _GEN_3134 = 14'hc3e == index ? 14'h18 : _GEN_3133;
  wire [13:0] _GEN_3135 = 14'hc3f == index ? 14'h18 : _GEN_3134;
  wire [13:0] _GEN_3136 = 14'hc40 == index ? 14'h18 : _GEN_3135;
  wire [13:0] _GEN_3137 = 14'hc41 == index ? 14'h18 : _GEN_3136;
  wire [13:0] _GEN_3138 = 14'hc42 == index ? 14'h18 : _GEN_3137;
  wire [13:0] _GEN_3139 = 14'hc43 == index ? 14'h18 : _GEN_3138;
  wire [13:0] _GEN_3140 = 14'hc44 == index ? 14'h18 : _GEN_3139;
  wire [13:0] _GEN_3141 = 14'hc45 == index ? 14'h18 : _GEN_3140;
  wire [13:0] _GEN_3142 = 14'hc46 == index ? 14'h18 : _GEN_3141;
  wire [13:0] _GEN_3143 = 14'hc47 == index ? 14'h18 : _GEN_3142;
  wire [13:0] _GEN_3144 = 14'hc48 == index ? 14'h18 : _GEN_3143;
  wire [13:0] _GEN_3145 = 14'hc49 == index ? 14'h18 : _GEN_3144;
  wire [13:0] _GEN_3146 = 14'hc4a == index ? 14'h18 : _GEN_3145;
  wire [13:0] _GEN_3147 = 14'hc4b == index ? 14'h18 : _GEN_3146;
  wire [13:0] _GEN_3148 = 14'hc4c == index ? 14'h18 : _GEN_3147;
  wire [13:0] _GEN_3149 = 14'hc4d == index ? 14'h18 : _GEN_3148;
  wire [13:0] _GEN_3150 = 14'hc4e == index ? 14'h18 : _GEN_3149;
  wire [13:0] _GEN_3151 = 14'hc4f == index ? 14'h18 : _GEN_3150;
  wire [13:0] _GEN_3152 = 14'hc50 == index ? 14'h18 : _GEN_3151;
  wire [13:0] _GEN_3153 = 14'hc51 == index ? 14'h18 : _GEN_3152;
  wire [13:0] _GEN_3154 = 14'hc52 == index ? 14'h18 : _GEN_3153;
  wire [13:0] _GEN_3155 = 14'hc53 == index ? 14'h18 : _GEN_3154;
  wire [13:0] _GEN_3156 = 14'hc54 == index ? 14'h18 : _GEN_3155;
  wire [13:0] _GEN_3157 = 14'hc55 == index ? 14'h18 : _GEN_3156;
  wire [13:0] _GEN_3158 = 14'hc56 == index ? 14'h18 : _GEN_3157;
  wire [13:0] _GEN_3159 = 14'hc57 == index ? 14'h18 : _GEN_3158;
  wire [13:0] _GEN_3160 = 14'hc58 == index ? 14'h18 : _GEN_3159;
  wire [13:0] _GEN_3161 = 14'hc59 == index ? 14'h18 : _GEN_3160;
  wire [13:0] _GEN_3162 = 14'hc5a == index ? 14'h18 : _GEN_3161;
  wire [13:0] _GEN_3163 = 14'hc5b == index ? 14'h18 : _GEN_3162;
  wire [13:0] _GEN_3164 = 14'hc5c == index ? 14'h18 : _GEN_3163;
  wire [13:0] _GEN_3165 = 14'hc5d == index ? 14'h18 : _GEN_3164;
  wire [13:0] _GEN_3166 = 14'hc5e == index ? 14'h18 : _GEN_3165;
  wire [13:0] _GEN_3167 = 14'hc5f == index ? 14'h18 : _GEN_3166;
  wire [13:0] _GEN_3168 = 14'hc60 == index ? 14'h18 : _GEN_3167;
  wire [13:0] _GEN_3169 = 14'hc61 == index ? 14'h18 : _GEN_3168;
  wire [13:0] _GEN_3170 = 14'hc62 == index ? 14'h18 : _GEN_3169;
  wire [13:0] _GEN_3171 = 14'hc63 == index ? 14'h18 : _GEN_3170;
  wire [13:0] _GEN_3172 = 14'hc64 == index ? 14'h18 : _GEN_3171;
  wire [13:0] _GEN_3173 = 14'hc65 == index ? 14'h18 : _GEN_3172;
  wire [13:0] _GEN_3174 = 14'hc66 == index ? 14'h18 : _GEN_3173;
  wire [13:0] _GEN_3175 = 14'hc67 == index ? 14'h18 : _GEN_3174;
  wire [13:0] _GEN_3176 = 14'hc68 == index ? 14'h18 : _GEN_3175;
  wire [13:0] _GEN_3177 = 14'hc69 == index ? 14'h18 : _GEN_3176;
  wire [13:0] _GEN_3178 = 14'hc6a == index ? 14'h18 : _GEN_3177;
  wire [13:0] _GEN_3179 = 14'hc6b == index ? 14'h18 : _GEN_3178;
  wire [13:0] _GEN_3180 = 14'hc6c == index ? 14'h18 : _GEN_3179;
  wire [13:0] _GEN_3181 = 14'hc6d == index ? 14'h18 : _GEN_3180;
  wire [13:0] _GEN_3182 = 14'hc6e == index ? 14'h18 : _GEN_3181;
  wire [13:0] _GEN_3183 = 14'hc6f == index ? 14'h18 : _GEN_3182;
  wire [13:0] _GEN_3184 = 14'hc70 == index ? 14'h18 : _GEN_3183;
  wire [13:0] _GEN_3185 = 14'hc71 == index ? 14'h18 : _GEN_3184;
  wire [13:0] _GEN_3186 = 14'hc72 == index ? 14'h18 : _GEN_3185;
  wire [13:0] _GEN_3187 = 14'hc73 == index ? 14'h18 : _GEN_3186;
  wire [13:0] _GEN_3188 = 14'hc74 == index ? 14'h18 : _GEN_3187;
  wire [13:0] _GEN_3189 = 14'hc75 == index ? 14'h18 : _GEN_3188;
  wire [13:0] _GEN_3190 = 14'hc76 == index ? 14'h18 : _GEN_3189;
  wire [13:0] _GEN_3191 = 14'hc77 == index ? 14'h18 : _GEN_3190;
  wire [13:0] _GEN_3192 = 14'hc78 == index ? 14'h18 : _GEN_3191;
  wire [13:0] _GEN_3193 = 14'hc79 == index ? 14'h18 : _GEN_3192;
  wire [13:0] _GEN_3194 = 14'hc7a == index ? 14'h18 : _GEN_3193;
  wire [13:0] _GEN_3195 = 14'hc7b == index ? 14'h18 : _GEN_3194;
  wire [13:0] _GEN_3196 = 14'hc7c == index ? 14'h18 : _GEN_3195;
  wire [13:0] _GEN_3197 = 14'hc7d == index ? 14'h18 : _GEN_3196;
  wire [13:0] _GEN_3198 = 14'hc7e == index ? 14'h18 : _GEN_3197;
  wire [13:0] _GEN_3199 = 14'hc7f == index ? 14'h18 : _GEN_3198;
  wire [13:0] _GEN_3200 = 14'hc80 == index ? 14'h0 : _GEN_3199;
  wire [13:0] _GEN_3201 = 14'hc81 == index ? 14'hc80 : _GEN_3200;
  wire [13:0] _GEN_3202 = 14'hc82 == index ? 14'h601 : _GEN_3201;
  wire [13:0] _GEN_3203 = 14'hc83 == index ? 14'h401 : _GEN_3202;
  wire [13:0] _GEN_3204 = 14'hc84 == index ? 14'h301 : _GEN_3203;
  wire [13:0] _GEN_3205 = 14'hc85 == index ? 14'h280 : _GEN_3204;
  wire [13:0] _GEN_3206 = 14'hc86 == index ? 14'h201 : _GEN_3205;
  wire [13:0] _GEN_3207 = 14'hc87 == index ? 14'h184 : _GEN_3206;
  wire [13:0] _GEN_3208 = 14'hc88 == index ? 14'h181 : _GEN_3207;
  wire [13:0] _GEN_3209 = 14'hc89 == index ? 14'h107 : _GEN_3208;
  wire [13:0] _GEN_3210 = 14'hc8a == index ? 14'h105 : _GEN_3209;
  wire [13:0] _GEN_3211 = 14'hc8b == index ? 14'h103 : _GEN_3210;
  wire [13:0] _GEN_3212 = 14'hc8c == index ? 14'h101 : _GEN_3211;
  wire [13:0] _GEN_3213 = 14'hc8d == index ? 14'h8c : _GEN_3212;
  wire [13:0] _GEN_3214 = 14'hc8e == index ? 14'h8b : _GEN_3213;
  wire [13:0] _GEN_3215 = 14'hc8f == index ? 14'h8a : _GEN_3214;
  wire [13:0] _GEN_3216 = 14'hc90 == index ? 14'h89 : _GEN_3215;
  wire [13:0] _GEN_3217 = 14'hc91 == index ? 14'h88 : _GEN_3216;
  wire [13:0] _GEN_3218 = 14'hc92 == index ? 14'h87 : _GEN_3217;
  wire [13:0] _GEN_3219 = 14'hc93 == index ? 14'h86 : _GEN_3218;
  wire [13:0] _GEN_3220 = 14'hc94 == index ? 14'h85 : _GEN_3219;
  wire [13:0] _GEN_3221 = 14'hc95 == index ? 14'h84 : _GEN_3220;
  wire [13:0] _GEN_3222 = 14'hc96 == index ? 14'h83 : _GEN_3221;
  wire [13:0] _GEN_3223 = 14'hc97 == index ? 14'h82 : _GEN_3222;
  wire [13:0] _GEN_3224 = 14'hc98 == index ? 14'h81 : _GEN_3223;
  wire [13:0] _GEN_3225 = 14'hc99 == index ? 14'h80 : _GEN_3224;
  wire [13:0] _GEN_3226 = 14'hc9a == index ? 14'h19 : _GEN_3225;
  wire [13:0] _GEN_3227 = 14'hc9b == index ? 14'h19 : _GEN_3226;
  wire [13:0] _GEN_3228 = 14'hc9c == index ? 14'h19 : _GEN_3227;
  wire [13:0] _GEN_3229 = 14'hc9d == index ? 14'h19 : _GEN_3228;
  wire [13:0] _GEN_3230 = 14'hc9e == index ? 14'h19 : _GEN_3229;
  wire [13:0] _GEN_3231 = 14'hc9f == index ? 14'h19 : _GEN_3230;
  wire [13:0] _GEN_3232 = 14'hca0 == index ? 14'h19 : _GEN_3231;
  wire [13:0] _GEN_3233 = 14'hca1 == index ? 14'h19 : _GEN_3232;
  wire [13:0] _GEN_3234 = 14'hca2 == index ? 14'h19 : _GEN_3233;
  wire [13:0] _GEN_3235 = 14'hca3 == index ? 14'h19 : _GEN_3234;
  wire [13:0] _GEN_3236 = 14'hca4 == index ? 14'h19 : _GEN_3235;
  wire [13:0] _GEN_3237 = 14'hca5 == index ? 14'h19 : _GEN_3236;
  wire [13:0] _GEN_3238 = 14'hca6 == index ? 14'h19 : _GEN_3237;
  wire [13:0] _GEN_3239 = 14'hca7 == index ? 14'h19 : _GEN_3238;
  wire [13:0] _GEN_3240 = 14'hca8 == index ? 14'h19 : _GEN_3239;
  wire [13:0] _GEN_3241 = 14'hca9 == index ? 14'h19 : _GEN_3240;
  wire [13:0] _GEN_3242 = 14'hcaa == index ? 14'h19 : _GEN_3241;
  wire [13:0] _GEN_3243 = 14'hcab == index ? 14'h19 : _GEN_3242;
  wire [13:0] _GEN_3244 = 14'hcac == index ? 14'h19 : _GEN_3243;
  wire [13:0] _GEN_3245 = 14'hcad == index ? 14'h19 : _GEN_3244;
  wire [13:0] _GEN_3246 = 14'hcae == index ? 14'h19 : _GEN_3245;
  wire [13:0] _GEN_3247 = 14'hcaf == index ? 14'h19 : _GEN_3246;
  wire [13:0] _GEN_3248 = 14'hcb0 == index ? 14'h19 : _GEN_3247;
  wire [13:0] _GEN_3249 = 14'hcb1 == index ? 14'h19 : _GEN_3248;
  wire [13:0] _GEN_3250 = 14'hcb2 == index ? 14'h19 : _GEN_3249;
  wire [13:0] _GEN_3251 = 14'hcb3 == index ? 14'h19 : _GEN_3250;
  wire [13:0] _GEN_3252 = 14'hcb4 == index ? 14'h19 : _GEN_3251;
  wire [13:0] _GEN_3253 = 14'hcb5 == index ? 14'h19 : _GEN_3252;
  wire [13:0] _GEN_3254 = 14'hcb6 == index ? 14'h19 : _GEN_3253;
  wire [13:0] _GEN_3255 = 14'hcb7 == index ? 14'h19 : _GEN_3254;
  wire [13:0] _GEN_3256 = 14'hcb8 == index ? 14'h19 : _GEN_3255;
  wire [13:0] _GEN_3257 = 14'hcb9 == index ? 14'h19 : _GEN_3256;
  wire [13:0] _GEN_3258 = 14'hcba == index ? 14'h19 : _GEN_3257;
  wire [13:0] _GEN_3259 = 14'hcbb == index ? 14'h19 : _GEN_3258;
  wire [13:0] _GEN_3260 = 14'hcbc == index ? 14'h19 : _GEN_3259;
  wire [13:0] _GEN_3261 = 14'hcbd == index ? 14'h19 : _GEN_3260;
  wire [13:0] _GEN_3262 = 14'hcbe == index ? 14'h19 : _GEN_3261;
  wire [13:0] _GEN_3263 = 14'hcbf == index ? 14'h19 : _GEN_3262;
  wire [13:0] _GEN_3264 = 14'hcc0 == index ? 14'h19 : _GEN_3263;
  wire [13:0] _GEN_3265 = 14'hcc1 == index ? 14'h19 : _GEN_3264;
  wire [13:0] _GEN_3266 = 14'hcc2 == index ? 14'h19 : _GEN_3265;
  wire [13:0] _GEN_3267 = 14'hcc3 == index ? 14'h19 : _GEN_3266;
  wire [13:0] _GEN_3268 = 14'hcc4 == index ? 14'h19 : _GEN_3267;
  wire [13:0] _GEN_3269 = 14'hcc5 == index ? 14'h19 : _GEN_3268;
  wire [13:0] _GEN_3270 = 14'hcc6 == index ? 14'h19 : _GEN_3269;
  wire [13:0] _GEN_3271 = 14'hcc7 == index ? 14'h19 : _GEN_3270;
  wire [13:0] _GEN_3272 = 14'hcc8 == index ? 14'h19 : _GEN_3271;
  wire [13:0] _GEN_3273 = 14'hcc9 == index ? 14'h19 : _GEN_3272;
  wire [13:0] _GEN_3274 = 14'hcca == index ? 14'h19 : _GEN_3273;
  wire [13:0] _GEN_3275 = 14'hccb == index ? 14'h19 : _GEN_3274;
  wire [13:0] _GEN_3276 = 14'hccc == index ? 14'h19 : _GEN_3275;
  wire [13:0] _GEN_3277 = 14'hccd == index ? 14'h19 : _GEN_3276;
  wire [13:0] _GEN_3278 = 14'hcce == index ? 14'h19 : _GEN_3277;
  wire [13:0] _GEN_3279 = 14'hccf == index ? 14'h19 : _GEN_3278;
  wire [13:0] _GEN_3280 = 14'hcd0 == index ? 14'h19 : _GEN_3279;
  wire [13:0] _GEN_3281 = 14'hcd1 == index ? 14'h19 : _GEN_3280;
  wire [13:0] _GEN_3282 = 14'hcd2 == index ? 14'h19 : _GEN_3281;
  wire [13:0] _GEN_3283 = 14'hcd3 == index ? 14'h19 : _GEN_3282;
  wire [13:0] _GEN_3284 = 14'hcd4 == index ? 14'h19 : _GEN_3283;
  wire [13:0] _GEN_3285 = 14'hcd5 == index ? 14'h19 : _GEN_3284;
  wire [13:0] _GEN_3286 = 14'hcd6 == index ? 14'h19 : _GEN_3285;
  wire [13:0] _GEN_3287 = 14'hcd7 == index ? 14'h19 : _GEN_3286;
  wire [13:0] _GEN_3288 = 14'hcd8 == index ? 14'h19 : _GEN_3287;
  wire [13:0] _GEN_3289 = 14'hcd9 == index ? 14'h19 : _GEN_3288;
  wire [13:0] _GEN_3290 = 14'hcda == index ? 14'h19 : _GEN_3289;
  wire [13:0] _GEN_3291 = 14'hcdb == index ? 14'h19 : _GEN_3290;
  wire [13:0] _GEN_3292 = 14'hcdc == index ? 14'h19 : _GEN_3291;
  wire [13:0] _GEN_3293 = 14'hcdd == index ? 14'h19 : _GEN_3292;
  wire [13:0] _GEN_3294 = 14'hcde == index ? 14'h19 : _GEN_3293;
  wire [13:0] _GEN_3295 = 14'hcdf == index ? 14'h19 : _GEN_3294;
  wire [13:0] _GEN_3296 = 14'hce0 == index ? 14'h19 : _GEN_3295;
  wire [13:0] _GEN_3297 = 14'hce1 == index ? 14'h19 : _GEN_3296;
  wire [13:0] _GEN_3298 = 14'hce2 == index ? 14'h19 : _GEN_3297;
  wire [13:0] _GEN_3299 = 14'hce3 == index ? 14'h19 : _GEN_3298;
  wire [13:0] _GEN_3300 = 14'hce4 == index ? 14'h19 : _GEN_3299;
  wire [13:0] _GEN_3301 = 14'hce5 == index ? 14'h19 : _GEN_3300;
  wire [13:0] _GEN_3302 = 14'hce6 == index ? 14'h19 : _GEN_3301;
  wire [13:0] _GEN_3303 = 14'hce7 == index ? 14'h19 : _GEN_3302;
  wire [13:0] _GEN_3304 = 14'hce8 == index ? 14'h19 : _GEN_3303;
  wire [13:0] _GEN_3305 = 14'hce9 == index ? 14'h19 : _GEN_3304;
  wire [13:0] _GEN_3306 = 14'hcea == index ? 14'h19 : _GEN_3305;
  wire [13:0] _GEN_3307 = 14'hceb == index ? 14'h19 : _GEN_3306;
  wire [13:0] _GEN_3308 = 14'hcec == index ? 14'h19 : _GEN_3307;
  wire [13:0] _GEN_3309 = 14'hced == index ? 14'h19 : _GEN_3308;
  wire [13:0] _GEN_3310 = 14'hcee == index ? 14'h19 : _GEN_3309;
  wire [13:0] _GEN_3311 = 14'hcef == index ? 14'h19 : _GEN_3310;
  wire [13:0] _GEN_3312 = 14'hcf0 == index ? 14'h19 : _GEN_3311;
  wire [13:0] _GEN_3313 = 14'hcf1 == index ? 14'h19 : _GEN_3312;
  wire [13:0] _GEN_3314 = 14'hcf2 == index ? 14'h19 : _GEN_3313;
  wire [13:0] _GEN_3315 = 14'hcf3 == index ? 14'h19 : _GEN_3314;
  wire [13:0] _GEN_3316 = 14'hcf4 == index ? 14'h19 : _GEN_3315;
  wire [13:0] _GEN_3317 = 14'hcf5 == index ? 14'h19 : _GEN_3316;
  wire [13:0] _GEN_3318 = 14'hcf6 == index ? 14'h19 : _GEN_3317;
  wire [13:0] _GEN_3319 = 14'hcf7 == index ? 14'h19 : _GEN_3318;
  wire [13:0] _GEN_3320 = 14'hcf8 == index ? 14'h19 : _GEN_3319;
  wire [13:0] _GEN_3321 = 14'hcf9 == index ? 14'h19 : _GEN_3320;
  wire [13:0] _GEN_3322 = 14'hcfa == index ? 14'h19 : _GEN_3321;
  wire [13:0] _GEN_3323 = 14'hcfb == index ? 14'h19 : _GEN_3322;
  wire [13:0] _GEN_3324 = 14'hcfc == index ? 14'h19 : _GEN_3323;
  wire [13:0] _GEN_3325 = 14'hcfd == index ? 14'h19 : _GEN_3324;
  wire [13:0] _GEN_3326 = 14'hcfe == index ? 14'h19 : _GEN_3325;
  wire [13:0] _GEN_3327 = 14'hcff == index ? 14'h19 : _GEN_3326;
  wire [13:0] _GEN_3328 = 14'hd00 == index ? 14'h0 : _GEN_3327;
  wire [13:0] _GEN_3329 = 14'hd01 == index ? 14'hd00 : _GEN_3328;
  wire [13:0] _GEN_3330 = 14'hd02 == index ? 14'h680 : _GEN_3329;
  wire [13:0] _GEN_3331 = 14'hd03 == index ? 14'h402 : _GEN_3330;
  wire [13:0] _GEN_3332 = 14'hd04 == index ? 14'h302 : _GEN_3331;
  wire [13:0] _GEN_3333 = 14'hd05 == index ? 14'h281 : _GEN_3332;
  wire [13:0] _GEN_3334 = 14'hd06 == index ? 14'h202 : _GEN_3333;
  wire [13:0] _GEN_3335 = 14'hd07 == index ? 14'h185 : _GEN_3334;
  wire [13:0] _GEN_3336 = 14'hd08 == index ? 14'h182 : _GEN_3335;
  wire [13:0] _GEN_3337 = 14'hd09 == index ? 14'h108 : _GEN_3336;
  wire [13:0] _GEN_3338 = 14'hd0a == index ? 14'h106 : _GEN_3337;
  wire [13:0] _GEN_3339 = 14'hd0b == index ? 14'h104 : _GEN_3338;
  wire [13:0] _GEN_3340 = 14'hd0c == index ? 14'h102 : _GEN_3339;
  wire [13:0] _GEN_3341 = 14'hd0d == index ? 14'h100 : _GEN_3340;
  wire [13:0] _GEN_3342 = 14'hd0e == index ? 14'h8c : _GEN_3341;
  wire [13:0] _GEN_3343 = 14'hd0f == index ? 14'h8b : _GEN_3342;
  wire [13:0] _GEN_3344 = 14'hd10 == index ? 14'h8a : _GEN_3343;
  wire [13:0] _GEN_3345 = 14'hd11 == index ? 14'h89 : _GEN_3344;
  wire [13:0] _GEN_3346 = 14'hd12 == index ? 14'h88 : _GEN_3345;
  wire [13:0] _GEN_3347 = 14'hd13 == index ? 14'h87 : _GEN_3346;
  wire [13:0] _GEN_3348 = 14'hd14 == index ? 14'h86 : _GEN_3347;
  wire [13:0] _GEN_3349 = 14'hd15 == index ? 14'h85 : _GEN_3348;
  wire [13:0] _GEN_3350 = 14'hd16 == index ? 14'h84 : _GEN_3349;
  wire [13:0] _GEN_3351 = 14'hd17 == index ? 14'h83 : _GEN_3350;
  wire [13:0] _GEN_3352 = 14'hd18 == index ? 14'h82 : _GEN_3351;
  wire [13:0] _GEN_3353 = 14'hd19 == index ? 14'h81 : _GEN_3352;
  wire [13:0] _GEN_3354 = 14'hd1a == index ? 14'h80 : _GEN_3353;
  wire [13:0] _GEN_3355 = 14'hd1b == index ? 14'h1a : _GEN_3354;
  wire [13:0] _GEN_3356 = 14'hd1c == index ? 14'h1a : _GEN_3355;
  wire [13:0] _GEN_3357 = 14'hd1d == index ? 14'h1a : _GEN_3356;
  wire [13:0] _GEN_3358 = 14'hd1e == index ? 14'h1a : _GEN_3357;
  wire [13:0] _GEN_3359 = 14'hd1f == index ? 14'h1a : _GEN_3358;
  wire [13:0] _GEN_3360 = 14'hd20 == index ? 14'h1a : _GEN_3359;
  wire [13:0] _GEN_3361 = 14'hd21 == index ? 14'h1a : _GEN_3360;
  wire [13:0] _GEN_3362 = 14'hd22 == index ? 14'h1a : _GEN_3361;
  wire [13:0] _GEN_3363 = 14'hd23 == index ? 14'h1a : _GEN_3362;
  wire [13:0] _GEN_3364 = 14'hd24 == index ? 14'h1a : _GEN_3363;
  wire [13:0] _GEN_3365 = 14'hd25 == index ? 14'h1a : _GEN_3364;
  wire [13:0] _GEN_3366 = 14'hd26 == index ? 14'h1a : _GEN_3365;
  wire [13:0] _GEN_3367 = 14'hd27 == index ? 14'h1a : _GEN_3366;
  wire [13:0] _GEN_3368 = 14'hd28 == index ? 14'h1a : _GEN_3367;
  wire [13:0] _GEN_3369 = 14'hd29 == index ? 14'h1a : _GEN_3368;
  wire [13:0] _GEN_3370 = 14'hd2a == index ? 14'h1a : _GEN_3369;
  wire [13:0] _GEN_3371 = 14'hd2b == index ? 14'h1a : _GEN_3370;
  wire [13:0] _GEN_3372 = 14'hd2c == index ? 14'h1a : _GEN_3371;
  wire [13:0] _GEN_3373 = 14'hd2d == index ? 14'h1a : _GEN_3372;
  wire [13:0] _GEN_3374 = 14'hd2e == index ? 14'h1a : _GEN_3373;
  wire [13:0] _GEN_3375 = 14'hd2f == index ? 14'h1a : _GEN_3374;
  wire [13:0] _GEN_3376 = 14'hd30 == index ? 14'h1a : _GEN_3375;
  wire [13:0] _GEN_3377 = 14'hd31 == index ? 14'h1a : _GEN_3376;
  wire [13:0] _GEN_3378 = 14'hd32 == index ? 14'h1a : _GEN_3377;
  wire [13:0] _GEN_3379 = 14'hd33 == index ? 14'h1a : _GEN_3378;
  wire [13:0] _GEN_3380 = 14'hd34 == index ? 14'h1a : _GEN_3379;
  wire [13:0] _GEN_3381 = 14'hd35 == index ? 14'h1a : _GEN_3380;
  wire [13:0] _GEN_3382 = 14'hd36 == index ? 14'h1a : _GEN_3381;
  wire [13:0] _GEN_3383 = 14'hd37 == index ? 14'h1a : _GEN_3382;
  wire [13:0] _GEN_3384 = 14'hd38 == index ? 14'h1a : _GEN_3383;
  wire [13:0] _GEN_3385 = 14'hd39 == index ? 14'h1a : _GEN_3384;
  wire [13:0] _GEN_3386 = 14'hd3a == index ? 14'h1a : _GEN_3385;
  wire [13:0] _GEN_3387 = 14'hd3b == index ? 14'h1a : _GEN_3386;
  wire [13:0] _GEN_3388 = 14'hd3c == index ? 14'h1a : _GEN_3387;
  wire [13:0] _GEN_3389 = 14'hd3d == index ? 14'h1a : _GEN_3388;
  wire [13:0] _GEN_3390 = 14'hd3e == index ? 14'h1a : _GEN_3389;
  wire [13:0] _GEN_3391 = 14'hd3f == index ? 14'h1a : _GEN_3390;
  wire [13:0] _GEN_3392 = 14'hd40 == index ? 14'h1a : _GEN_3391;
  wire [13:0] _GEN_3393 = 14'hd41 == index ? 14'h1a : _GEN_3392;
  wire [13:0] _GEN_3394 = 14'hd42 == index ? 14'h1a : _GEN_3393;
  wire [13:0] _GEN_3395 = 14'hd43 == index ? 14'h1a : _GEN_3394;
  wire [13:0] _GEN_3396 = 14'hd44 == index ? 14'h1a : _GEN_3395;
  wire [13:0] _GEN_3397 = 14'hd45 == index ? 14'h1a : _GEN_3396;
  wire [13:0] _GEN_3398 = 14'hd46 == index ? 14'h1a : _GEN_3397;
  wire [13:0] _GEN_3399 = 14'hd47 == index ? 14'h1a : _GEN_3398;
  wire [13:0] _GEN_3400 = 14'hd48 == index ? 14'h1a : _GEN_3399;
  wire [13:0] _GEN_3401 = 14'hd49 == index ? 14'h1a : _GEN_3400;
  wire [13:0] _GEN_3402 = 14'hd4a == index ? 14'h1a : _GEN_3401;
  wire [13:0] _GEN_3403 = 14'hd4b == index ? 14'h1a : _GEN_3402;
  wire [13:0] _GEN_3404 = 14'hd4c == index ? 14'h1a : _GEN_3403;
  wire [13:0] _GEN_3405 = 14'hd4d == index ? 14'h1a : _GEN_3404;
  wire [13:0] _GEN_3406 = 14'hd4e == index ? 14'h1a : _GEN_3405;
  wire [13:0] _GEN_3407 = 14'hd4f == index ? 14'h1a : _GEN_3406;
  wire [13:0] _GEN_3408 = 14'hd50 == index ? 14'h1a : _GEN_3407;
  wire [13:0] _GEN_3409 = 14'hd51 == index ? 14'h1a : _GEN_3408;
  wire [13:0] _GEN_3410 = 14'hd52 == index ? 14'h1a : _GEN_3409;
  wire [13:0] _GEN_3411 = 14'hd53 == index ? 14'h1a : _GEN_3410;
  wire [13:0] _GEN_3412 = 14'hd54 == index ? 14'h1a : _GEN_3411;
  wire [13:0] _GEN_3413 = 14'hd55 == index ? 14'h1a : _GEN_3412;
  wire [13:0] _GEN_3414 = 14'hd56 == index ? 14'h1a : _GEN_3413;
  wire [13:0] _GEN_3415 = 14'hd57 == index ? 14'h1a : _GEN_3414;
  wire [13:0] _GEN_3416 = 14'hd58 == index ? 14'h1a : _GEN_3415;
  wire [13:0] _GEN_3417 = 14'hd59 == index ? 14'h1a : _GEN_3416;
  wire [13:0] _GEN_3418 = 14'hd5a == index ? 14'h1a : _GEN_3417;
  wire [13:0] _GEN_3419 = 14'hd5b == index ? 14'h1a : _GEN_3418;
  wire [13:0] _GEN_3420 = 14'hd5c == index ? 14'h1a : _GEN_3419;
  wire [13:0] _GEN_3421 = 14'hd5d == index ? 14'h1a : _GEN_3420;
  wire [13:0] _GEN_3422 = 14'hd5e == index ? 14'h1a : _GEN_3421;
  wire [13:0] _GEN_3423 = 14'hd5f == index ? 14'h1a : _GEN_3422;
  wire [13:0] _GEN_3424 = 14'hd60 == index ? 14'h1a : _GEN_3423;
  wire [13:0] _GEN_3425 = 14'hd61 == index ? 14'h1a : _GEN_3424;
  wire [13:0] _GEN_3426 = 14'hd62 == index ? 14'h1a : _GEN_3425;
  wire [13:0] _GEN_3427 = 14'hd63 == index ? 14'h1a : _GEN_3426;
  wire [13:0] _GEN_3428 = 14'hd64 == index ? 14'h1a : _GEN_3427;
  wire [13:0] _GEN_3429 = 14'hd65 == index ? 14'h1a : _GEN_3428;
  wire [13:0] _GEN_3430 = 14'hd66 == index ? 14'h1a : _GEN_3429;
  wire [13:0] _GEN_3431 = 14'hd67 == index ? 14'h1a : _GEN_3430;
  wire [13:0] _GEN_3432 = 14'hd68 == index ? 14'h1a : _GEN_3431;
  wire [13:0] _GEN_3433 = 14'hd69 == index ? 14'h1a : _GEN_3432;
  wire [13:0] _GEN_3434 = 14'hd6a == index ? 14'h1a : _GEN_3433;
  wire [13:0] _GEN_3435 = 14'hd6b == index ? 14'h1a : _GEN_3434;
  wire [13:0] _GEN_3436 = 14'hd6c == index ? 14'h1a : _GEN_3435;
  wire [13:0] _GEN_3437 = 14'hd6d == index ? 14'h1a : _GEN_3436;
  wire [13:0] _GEN_3438 = 14'hd6e == index ? 14'h1a : _GEN_3437;
  wire [13:0] _GEN_3439 = 14'hd6f == index ? 14'h1a : _GEN_3438;
  wire [13:0] _GEN_3440 = 14'hd70 == index ? 14'h1a : _GEN_3439;
  wire [13:0] _GEN_3441 = 14'hd71 == index ? 14'h1a : _GEN_3440;
  wire [13:0] _GEN_3442 = 14'hd72 == index ? 14'h1a : _GEN_3441;
  wire [13:0] _GEN_3443 = 14'hd73 == index ? 14'h1a : _GEN_3442;
  wire [13:0] _GEN_3444 = 14'hd74 == index ? 14'h1a : _GEN_3443;
  wire [13:0] _GEN_3445 = 14'hd75 == index ? 14'h1a : _GEN_3444;
  wire [13:0] _GEN_3446 = 14'hd76 == index ? 14'h1a : _GEN_3445;
  wire [13:0] _GEN_3447 = 14'hd77 == index ? 14'h1a : _GEN_3446;
  wire [13:0] _GEN_3448 = 14'hd78 == index ? 14'h1a : _GEN_3447;
  wire [13:0] _GEN_3449 = 14'hd79 == index ? 14'h1a : _GEN_3448;
  wire [13:0] _GEN_3450 = 14'hd7a == index ? 14'h1a : _GEN_3449;
  wire [13:0] _GEN_3451 = 14'hd7b == index ? 14'h1a : _GEN_3450;
  wire [13:0] _GEN_3452 = 14'hd7c == index ? 14'h1a : _GEN_3451;
  wire [13:0] _GEN_3453 = 14'hd7d == index ? 14'h1a : _GEN_3452;
  wire [13:0] _GEN_3454 = 14'hd7e == index ? 14'h1a : _GEN_3453;
  wire [13:0] _GEN_3455 = 14'hd7f == index ? 14'h1a : _GEN_3454;
  wire [13:0] _GEN_3456 = 14'hd80 == index ? 14'h0 : _GEN_3455;
  wire [13:0] _GEN_3457 = 14'hd81 == index ? 14'hd80 : _GEN_3456;
  wire [13:0] _GEN_3458 = 14'hd82 == index ? 14'h681 : _GEN_3457;
  wire [13:0] _GEN_3459 = 14'hd83 == index ? 14'h480 : _GEN_3458;
  wire [13:0] _GEN_3460 = 14'hd84 == index ? 14'h303 : _GEN_3459;
  wire [13:0] _GEN_3461 = 14'hd85 == index ? 14'h282 : _GEN_3460;
  wire [13:0] _GEN_3462 = 14'hd86 == index ? 14'h203 : _GEN_3461;
  wire [13:0] _GEN_3463 = 14'hd87 == index ? 14'h186 : _GEN_3462;
  wire [13:0] _GEN_3464 = 14'hd88 == index ? 14'h183 : _GEN_3463;
  wire [13:0] _GEN_3465 = 14'hd89 == index ? 14'h180 : _GEN_3464;
  wire [13:0] _GEN_3466 = 14'hd8a == index ? 14'h107 : _GEN_3465;
  wire [13:0] _GEN_3467 = 14'hd8b == index ? 14'h105 : _GEN_3466;
  wire [13:0] _GEN_3468 = 14'hd8c == index ? 14'h103 : _GEN_3467;
  wire [13:0] _GEN_3469 = 14'hd8d == index ? 14'h101 : _GEN_3468;
  wire [13:0] _GEN_3470 = 14'hd8e == index ? 14'h8d : _GEN_3469;
  wire [13:0] _GEN_3471 = 14'hd8f == index ? 14'h8c : _GEN_3470;
  wire [13:0] _GEN_3472 = 14'hd90 == index ? 14'h8b : _GEN_3471;
  wire [13:0] _GEN_3473 = 14'hd91 == index ? 14'h8a : _GEN_3472;
  wire [13:0] _GEN_3474 = 14'hd92 == index ? 14'h89 : _GEN_3473;
  wire [13:0] _GEN_3475 = 14'hd93 == index ? 14'h88 : _GEN_3474;
  wire [13:0] _GEN_3476 = 14'hd94 == index ? 14'h87 : _GEN_3475;
  wire [13:0] _GEN_3477 = 14'hd95 == index ? 14'h86 : _GEN_3476;
  wire [13:0] _GEN_3478 = 14'hd96 == index ? 14'h85 : _GEN_3477;
  wire [13:0] _GEN_3479 = 14'hd97 == index ? 14'h84 : _GEN_3478;
  wire [13:0] _GEN_3480 = 14'hd98 == index ? 14'h83 : _GEN_3479;
  wire [13:0] _GEN_3481 = 14'hd99 == index ? 14'h82 : _GEN_3480;
  wire [13:0] _GEN_3482 = 14'hd9a == index ? 14'h81 : _GEN_3481;
  wire [13:0] _GEN_3483 = 14'hd9b == index ? 14'h80 : _GEN_3482;
  wire [13:0] _GEN_3484 = 14'hd9c == index ? 14'h1b : _GEN_3483;
  wire [13:0] _GEN_3485 = 14'hd9d == index ? 14'h1b : _GEN_3484;
  wire [13:0] _GEN_3486 = 14'hd9e == index ? 14'h1b : _GEN_3485;
  wire [13:0] _GEN_3487 = 14'hd9f == index ? 14'h1b : _GEN_3486;
  wire [13:0] _GEN_3488 = 14'hda0 == index ? 14'h1b : _GEN_3487;
  wire [13:0] _GEN_3489 = 14'hda1 == index ? 14'h1b : _GEN_3488;
  wire [13:0] _GEN_3490 = 14'hda2 == index ? 14'h1b : _GEN_3489;
  wire [13:0] _GEN_3491 = 14'hda3 == index ? 14'h1b : _GEN_3490;
  wire [13:0] _GEN_3492 = 14'hda4 == index ? 14'h1b : _GEN_3491;
  wire [13:0] _GEN_3493 = 14'hda5 == index ? 14'h1b : _GEN_3492;
  wire [13:0] _GEN_3494 = 14'hda6 == index ? 14'h1b : _GEN_3493;
  wire [13:0] _GEN_3495 = 14'hda7 == index ? 14'h1b : _GEN_3494;
  wire [13:0] _GEN_3496 = 14'hda8 == index ? 14'h1b : _GEN_3495;
  wire [13:0] _GEN_3497 = 14'hda9 == index ? 14'h1b : _GEN_3496;
  wire [13:0] _GEN_3498 = 14'hdaa == index ? 14'h1b : _GEN_3497;
  wire [13:0] _GEN_3499 = 14'hdab == index ? 14'h1b : _GEN_3498;
  wire [13:0] _GEN_3500 = 14'hdac == index ? 14'h1b : _GEN_3499;
  wire [13:0] _GEN_3501 = 14'hdad == index ? 14'h1b : _GEN_3500;
  wire [13:0] _GEN_3502 = 14'hdae == index ? 14'h1b : _GEN_3501;
  wire [13:0] _GEN_3503 = 14'hdaf == index ? 14'h1b : _GEN_3502;
  wire [13:0] _GEN_3504 = 14'hdb0 == index ? 14'h1b : _GEN_3503;
  wire [13:0] _GEN_3505 = 14'hdb1 == index ? 14'h1b : _GEN_3504;
  wire [13:0] _GEN_3506 = 14'hdb2 == index ? 14'h1b : _GEN_3505;
  wire [13:0] _GEN_3507 = 14'hdb3 == index ? 14'h1b : _GEN_3506;
  wire [13:0] _GEN_3508 = 14'hdb4 == index ? 14'h1b : _GEN_3507;
  wire [13:0] _GEN_3509 = 14'hdb5 == index ? 14'h1b : _GEN_3508;
  wire [13:0] _GEN_3510 = 14'hdb6 == index ? 14'h1b : _GEN_3509;
  wire [13:0] _GEN_3511 = 14'hdb7 == index ? 14'h1b : _GEN_3510;
  wire [13:0] _GEN_3512 = 14'hdb8 == index ? 14'h1b : _GEN_3511;
  wire [13:0] _GEN_3513 = 14'hdb9 == index ? 14'h1b : _GEN_3512;
  wire [13:0] _GEN_3514 = 14'hdba == index ? 14'h1b : _GEN_3513;
  wire [13:0] _GEN_3515 = 14'hdbb == index ? 14'h1b : _GEN_3514;
  wire [13:0] _GEN_3516 = 14'hdbc == index ? 14'h1b : _GEN_3515;
  wire [13:0] _GEN_3517 = 14'hdbd == index ? 14'h1b : _GEN_3516;
  wire [13:0] _GEN_3518 = 14'hdbe == index ? 14'h1b : _GEN_3517;
  wire [13:0] _GEN_3519 = 14'hdbf == index ? 14'h1b : _GEN_3518;
  wire [13:0] _GEN_3520 = 14'hdc0 == index ? 14'h1b : _GEN_3519;
  wire [13:0] _GEN_3521 = 14'hdc1 == index ? 14'h1b : _GEN_3520;
  wire [13:0] _GEN_3522 = 14'hdc2 == index ? 14'h1b : _GEN_3521;
  wire [13:0] _GEN_3523 = 14'hdc3 == index ? 14'h1b : _GEN_3522;
  wire [13:0] _GEN_3524 = 14'hdc4 == index ? 14'h1b : _GEN_3523;
  wire [13:0] _GEN_3525 = 14'hdc5 == index ? 14'h1b : _GEN_3524;
  wire [13:0] _GEN_3526 = 14'hdc6 == index ? 14'h1b : _GEN_3525;
  wire [13:0] _GEN_3527 = 14'hdc7 == index ? 14'h1b : _GEN_3526;
  wire [13:0] _GEN_3528 = 14'hdc8 == index ? 14'h1b : _GEN_3527;
  wire [13:0] _GEN_3529 = 14'hdc9 == index ? 14'h1b : _GEN_3528;
  wire [13:0] _GEN_3530 = 14'hdca == index ? 14'h1b : _GEN_3529;
  wire [13:0] _GEN_3531 = 14'hdcb == index ? 14'h1b : _GEN_3530;
  wire [13:0] _GEN_3532 = 14'hdcc == index ? 14'h1b : _GEN_3531;
  wire [13:0] _GEN_3533 = 14'hdcd == index ? 14'h1b : _GEN_3532;
  wire [13:0] _GEN_3534 = 14'hdce == index ? 14'h1b : _GEN_3533;
  wire [13:0] _GEN_3535 = 14'hdcf == index ? 14'h1b : _GEN_3534;
  wire [13:0] _GEN_3536 = 14'hdd0 == index ? 14'h1b : _GEN_3535;
  wire [13:0] _GEN_3537 = 14'hdd1 == index ? 14'h1b : _GEN_3536;
  wire [13:0] _GEN_3538 = 14'hdd2 == index ? 14'h1b : _GEN_3537;
  wire [13:0] _GEN_3539 = 14'hdd3 == index ? 14'h1b : _GEN_3538;
  wire [13:0] _GEN_3540 = 14'hdd4 == index ? 14'h1b : _GEN_3539;
  wire [13:0] _GEN_3541 = 14'hdd5 == index ? 14'h1b : _GEN_3540;
  wire [13:0] _GEN_3542 = 14'hdd6 == index ? 14'h1b : _GEN_3541;
  wire [13:0] _GEN_3543 = 14'hdd7 == index ? 14'h1b : _GEN_3542;
  wire [13:0] _GEN_3544 = 14'hdd8 == index ? 14'h1b : _GEN_3543;
  wire [13:0] _GEN_3545 = 14'hdd9 == index ? 14'h1b : _GEN_3544;
  wire [13:0] _GEN_3546 = 14'hdda == index ? 14'h1b : _GEN_3545;
  wire [13:0] _GEN_3547 = 14'hddb == index ? 14'h1b : _GEN_3546;
  wire [13:0] _GEN_3548 = 14'hddc == index ? 14'h1b : _GEN_3547;
  wire [13:0] _GEN_3549 = 14'hddd == index ? 14'h1b : _GEN_3548;
  wire [13:0] _GEN_3550 = 14'hdde == index ? 14'h1b : _GEN_3549;
  wire [13:0] _GEN_3551 = 14'hddf == index ? 14'h1b : _GEN_3550;
  wire [13:0] _GEN_3552 = 14'hde0 == index ? 14'h1b : _GEN_3551;
  wire [13:0] _GEN_3553 = 14'hde1 == index ? 14'h1b : _GEN_3552;
  wire [13:0] _GEN_3554 = 14'hde2 == index ? 14'h1b : _GEN_3553;
  wire [13:0] _GEN_3555 = 14'hde3 == index ? 14'h1b : _GEN_3554;
  wire [13:0] _GEN_3556 = 14'hde4 == index ? 14'h1b : _GEN_3555;
  wire [13:0] _GEN_3557 = 14'hde5 == index ? 14'h1b : _GEN_3556;
  wire [13:0] _GEN_3558 = 14'hde6 == index ? 14'h1b : _GEN_3557;
  wire [13:0] _GEN_3559 = 14'hde7 == index ? 14'h1b : _GEN_3558;
  wire [13:0] _GEN_3560 = 14'hde8 == index ? 14'h1b : _GEN_3559;
  wire [13:0] _GEN_3561 = 14'hde9 == index ? 14'h1b : _GEN_3560;
  wire [13:0] _GEN_3562 = 14'hdea == index ? 14'h1b : _GEN_3561;
  wire [13:0] _GEN_3563 = 14'hdeb == index ? 14'h1b : _GEN_3562;
  wire [13:0] _GEN_3564 = 14'hdec == index ? 14'h1b : _GEN_3563;
  wire [13:0] _GEN_3565 = 14'hded == index ? 14'h1b : _GEN_3564;
  wire [13:0] _GEN_3566 = 14'hdee == index ? 14'h1b : _GEN_3565;
  wire [13:0] _GEN_3567 = 14'hdef == index ? 14'h1b : _GEN_3566;
  wire [13:0] _GEN_3568 = 14'hdf0 == index ? 14'h1b : _GEN_3567;
  wire [13:0] _GEN_3569 = 14'hdf1 == index ? 14'h1b : _GEN_3568;
  wire [13:0] _GEN_3570 = 14'hdf2 == index ? 14'h1b : _GEN_3569;
  wire [13:0] _GEN_3571 = 14'hdf3 == index ? 14'h1b : _GEN_3570;
  wire [13:0] _GEN_3572 = 14'hdf4 == index ? 14'h1b : _GEN_3571;
  wire [13:0] _GEN_3573 = 14'hdf5 == index ? 14'h1b : _GEN_3572;
  wire [13:0] _GEN_3574 = 14'hdf6 == index ? 14'h1b : _GEN_3573;
  wire [13:0] _GEN_3575 = 14'hdf7 == index ? 14'h1b : _GEN_3574;
  wire [13:0] _GEN_3576 = 14'hdf8 == index ? 14'h1b : _GEN_3575;
  wire [13:0] _GEN_3577 = 14'hdf9 == index ? 14'h1b : _GEN_3576;
  wire [13:0] _GEN_3578 = 14'hdfa == index ? 14'h1b : _GEN_3577;
  wire [13:0] _GEN_3579 = 14'hdfb == index ? 14'h1b : _GEN_3578;
  wire [13:0] _GEN_3580 = 14'hdfc == index ? 14'h1b : _GEN_3579;
  wire [13:0] _GEN_3581 = 14'hdfd == index ? 14'h1b : _GEN_3580;
  wire [13:0] _GEN_3582 = 14'hdfe == index ? 14'h1b : _GEN_3581;
  wire [13:0] _GEN_3583 = 14'hdff == index ? 14'h1b : _GEN_3582;
  wire [13:0] _GEN_3584 = 14'he00 == index ? 14'h0 : _GEN_3583;
  wire [13:0] _GEN_3585 = 14'he01 == index ? 14'he00 : _GEN_3584;
  wire [13:0] _GEN_3586 = 14'he02 == index ? 14'h700 : _GEN_3585;
  wire [13:0] _GEN_3587 = 14'he03 == index ? 14'h481 : _GEN_3586;
  wire [13:0] _GEN_3588 = 14'he04 == index ? 14'h380 : _GEN_3587;
  wire [13:0] _GEN_3589 = 14'he05 == index ? 14'h283 : _GEN_3588;
  wire [13:0] _GEN_3590 = 14'he06 == index ? 14'h204 : _GEN_3589;
  wire [13:0] _GEN_3591 = 14'he07 == index ? 14'h200 : _GEN_3590;
  wire [13:0] _GEN_3592 = 14'he08 == index ? 14'h184 : _GEN_3591;
  wire [13:0] _GEN_3593 = 14'he09 == index ? 14'h181 : _GEN_3592;
  wire [13:0] _GEN_3594 = 14'he0a == index ? 14'h108 : _GEN_3593;
  wire [13:0] _GEN_3595 = 14'he0b == index ? 14'h106 : _GEN_3594;
  wire [13:0] _GEN_3596 = 14'he0c == index ? 14'h104 : _GEN_3595;
  wire [13:0] _GEN_3597 = 14'he0d == index ? 14'h102 : _GEN_3596;
  wire [13:0] _GEN_3598 = 14'he0e == index ? 14'h100 : _GEN_3597;
  wire [13:0] _GEN_3599 = 14'he0f == index ? 14'h8d : _GEN_3598;
  wire [13:0] _GEN_3600 = 14'he10 == index ? 14'h8c : _GEN_3599;
  wire [13:0] _GEN_3601 = 14'he11 == index ? 14'h8b : _GEN_3600;
  wire [13:0] _GEN_3602 = 14'he12 == index ? 14'h8a : _GEN_3601;
  wire [13:0] _GEN_3603 = 14'he13 == index ? 14'h89 : _GEN_3602;
  wire [13:0] _GEN_3604 = 14'he14 == index ? 14'h88 : _GEN_3603;
  wire [13:0] _GEN_3605 = 14'he15 == index ? 14'h87 : _GEN_3604;
  wire [13:0] _GEN_3606 = 14'he16 == index ? 14'h86 : _GEN_3605;
  wire [13:0] _GEN_3607 = 14'he17 == index ? 14'h85 : _GEN_3606;
  wire [13:0] _GEN_3608 = 14'he18 == index ? 14'h84 : _GEN_3607;
  wire [13:0] _GEN_3609 = 14'he19 == index ? 14'h83 : _GEN_3608;
  wire [13:0] _GEN_3610 = 14'he1a == index ? 14'h82 : _GEN_3609;
  wire [13:0] _GEN_3611 = 14'he1b == index ? 14'h81 : _GEN_3610;
  wire [13:0] _GEN_3612 = 14'he1c == index ? 14'h80 : _GEN_3611;
  wire [13:0] _GEN_3613 = 14'he1d == index ? 14'h1c : _GEN_3612;
  wire [13:0] _GEN_3614 = 14'he1e == index ? 14'h1c : _GEN_3613;
  wire [13:0] _GEN_3615 = 14'he1f == index ? 14'h1c : _GEN_3614;
  wire [13:0] _GEN_3616 = 14'he20 == index ? 14'h1c : _GEN_3615;
  wire [13:0] _GEN_3617 = 14'he21 == index ? 14'h1c : _GEN_3616;
  wire [13:0] _GEN_3618 = 14'he22 == index ? 14'h1c : _GEN_3617;
  wire [13:0] _GEN_3619 = 14'he23 == index ? 14'h1c : _GEN_3618;
  wire [13:0] _GEN_3620 = 14'he24 == index ? 14'h1c : _GEN_3619;
  wire [13:0] _GEN_3621 = 14'he25 == index ? 14'h1c : _GEN_3620;
  wire [13:0] _GEN_3622 = 14'he26 == index ? 14'h1c : _GEN_3621;
  wire [13:0] _GEN_3623 = 14'he27 == index ? 14'h1c : _GEN_3622;
  wire [13:0] _GEN_3624 = 14'he28 == index ? 14'h1c : _GEN_3623;
  wire [13:0] _GEN_3625 = 14'he29 == index ? 14'h1c : _GEN_3624;
  wire [13:0] _GEN_3626 = 14'he2a == index ? 14'h1c : _GEN_3625;
  wire [13:0] _GEN_3627 = 14'he2b == index ? 14'h1c : _GEN_3626;
  wire [13:0] _GEN_3628 = 14'he2c == index ? 14'h1c : _GEN_3627;
  wire [13:0] _GEN_3629 = 14'he2d == index ? 14'h1c : _GEN_3628;
  wire [13:0] _GEN_3630 = 14'he2e == index ? 14'h1c : _GEN_3629;
  wire [13:0] _GEN_3631 = 14'he2f == index ? 14'h1c : _GEN_3630;
  wire [13:0] _GEN_3632 = 14'he30 == index ? 14'h1c : _GEN_3631;
  wire [13:0] _GEN_3633 = 14'he31 == index ? 14'h1c : _GEN_3632;
  wire [13:0] _GEN_3634 = 14'he32 == index ? 14'h1c : _GEN_3633;
  wire [13:0] _GEN_3635 = 14'he33 == index ? 14'h1c : _GEN_3634;
  wire [13:0] _GEN_3636 = 14'he34 == index ? 14'h1c : _GEN_3635;
  wire [13:0] _GEN_3637 = 14'he35 == index ? 14'h1c : _GEN_3636;
  wire [13:0] _GEN_3638 = 14'he36 == index ? 14'h1c : _GEN_3637;
  wire [13:0] _GEN_3639 = 14'he37 == index ? 14'h1c : _GEN_3638;
  wire [13:0] _GEN_3640 = 14'he38 == index ? 14'h1c : _GEN_3639;
  wire [13:0] _GEN_3641 = 14'he39 == index ? 14'h1c : _GEN_3640;
  wire [13:0] _GEN_3642 = 14'he3a == index ? 14'h1c : _GEN_3641;
  wire [13:0] _GEN_3643 = 14'he3b == index ? 14'h1c : _GEN_3642;
  wire [13:0] _GEN_3644 = 14'he3c == index ? 14'h1c : _GEN_3643;
  wire [13:0] _GEN_3645 = 14'he3d == index ? 14'h1c : _GEN_3644;
  wire [13:0] _GEN_3646 = 14'he3e == index ? 14'h1c : _GEN_3645;
  wire [13:0] _GEN_3647 = 14'he3f == index ? 14'h1c : _GEN_3646;
  wire [13:0] _GEN_3648 = 14'he40 == index ? 14'h1c : _GEN_3647;
  wire [13:0] _GEN_3649 = 14'he41 == index ? 14'h1c : _GEN_3648;
  wire [13:0] _GEN_3650 = 14'he42 == index ? 14'h1c : _GEN_3649;
  wire [13:0] _GEN_3651 = 14'he43 == index ? 14'h1c : _GEN_3650;
  wire [13:0] _GEN_3652 = 14'he44 == index ? 14'h1c : _GEN_3651;
  wire [13:0] _GEN_3653 = 14'he45 == index ? 14'h1c : _GEN_3652;
  wire [13:0] _GEN_3654 = 14'he46 == index ? 14'h1c : _GEN_3653;
  wire [13:0] _GEN_3655 = 14'he47 == index ? 14'h1c : _GEN_3654;
  wire [13:0] _GEN_3656 = 14'he48 == index ? 14'h1c : _GEN_3655;
  wire [13:0] _GEN_3657 = 14'he49 == index ? 14'h1c : _GEN_3656;
  wire [13:0] _GEN_3658 = 14'he4a == index ? 14'h1c : _GEN_3657;
  wire [13:0] _GEN_3659 = 14'he4b == index ? 14'h1c : _GEN_3658;
  wire [13:0] _GEN_3660 = 14'he4c == index ? 14'h1c : _GEN_3659;
  wire [13:0] _GEN_3661 = 14'he4d == index ? 14'h1c : _GEN_3660;
  wire [13:0] _GEN_3662 = 14'he4e == index ? 14'h1c : _GEN_3661;
  wire [13:0] _GEN_3663 = 14'he4f == index ? 14'h1c : _GEN_3662;
  wire [13:0] _GEN_3664 = 14'he50 == index ? 14'h1c : _GEN_3663;
  wire [13:0] _GEN_3665 = 14'he51 == index ? 14'h1c : _GEN_3664;
  wire [13:0] _GEN_3666 = 14'he52 == index ? 14'h1c : _GEN_3665;
  wire [13:0] _GEN_3667 = 14'he53 == index ? 14'h1c : _GEN_3666;
  wire [13:0] _GEN_3668 = 14'he54 == index ? 14'h1c : _GEN_3667;
  wire [13:0] _GEN_3669 = 14'he55 == index ? 14'h1c : _GEN_3668;
  wire [13:0] _GEN_3670 = 14'he56 == index ? 14'h1c : _GEN_3669;
  wire [13:0] _GEN_3671 = 14'he57 == index ? 14'h1c : _GEN_3670;
  wire [13:0] _GEN_3672 = 14'he58 == index ? 14'h1c : _GEN_3671;
  wire [13:0] _GEN_3673 = 14'he59 == index ? 14'h1c : _GEN_3672;
  wire [13:0] _GEN_3674 = 14'he5a == index ? 14'h1c : _GEN_3673;
  wire [13:0] _GEN_3675 = 14'he5b == index ? 14'h1c : _GEN_3674;
  wire [13:0] _GEN_3676 = 14'he5c == index ? 14'h1c : _GEN_3675;
  wire [13:0] _GEN_3677 = 14'he5d == index ? 14'h1c : _GEN_3676;
  wire [13:0] _GEN_3678 = 14'he5e == index ? 14'h1c : _GEN_3677;
  wire [13:0] _GEN_3679 = 14'he5f == index ? 14'h1c : _GEN_3678;
  wire [13:0] _GEN_3680 = 14'he60 == index ? 14'h1c : _GEN_3679;
  wire [13:0] _GEN_3681 = 14'he61 == index ? 14'h1c : _GEN_3680;
  wire [13:0] _GEN_3682 = 14'he62 == index ? 14'h1c : _GEN_3681;
  wire [13:0] _GEN_3683 = 14'he63 == index ? 14'h1c : _GEN_3682;
  wire [13:0] _GEN_3684 = 14'he64 == index ? 14'h1c : _GEN_3683;
  wire [13:0] _GEN_3685 = 14'he65 == index ? 14'h1c : _GEN_3684;
  wire [13:0] _GEN_3686 = 14'he66 == index ? 14'h1c : _GEN_3685;
  wire [13:0] _GEN_3687 = 14'he67 == index ? 14'h1c : _GEN_3686;
  wire [13:0] _GEN_3688 = 14'he68 == index ? 14'h1c : _GEN_3687;
  wire [13:0] _GEN_3689 = 14'he69 == index ? 14'h1c : _GEN_3688;
  wire [13:0] _GEN_3690 = 14'he6a == index ? 14'h1c : _GEN_3689;
  wire [13:0] _GEN_3691 = 14'he6b == index ? 14'h1c : _GEN_3690;
  wire [13:0] _GEN_3692 = 14'he6c == index ? 14'h1c : _GEN_3691;
  wire [13:0] _GEN_3693 = 14'he6d == index ? 14'h1c : _GEN_3692;
  wire [13:0] _GEN_3694 = 14'he6e == index ? 14'h1c : _GEN_3693;
  wire [13:0] _GEN_3695 = 14'he6f == index ? 14'h1c : _GEN_3694;
  wire [13:0] _GEN_3696 = 14'he70 == index ? 14'h1c : _GEN_3695;
  wire [13:0] _GEN_3697 = 14'he71 == index ? 14'h1c : _GEN_3696;
  wire [13:0] _GEN_3698 = 14'he72 == index ? 14'h1c : _GEN_3697;
  wire [13:0] _GEN_3699 = 14'he73 == index ? 14'h1c : _GEN_3698;
  wire [13:0] _GEN_3700 = 14'he74 == index ? 14'h1c : _GEN_3699;
  wire [13:0] _GEN_3701 = 14'he75 == index ? 14'h1c : _GEN_3700;
  wire [13:0] _GEN_3702 = 14'he76 == index ? 14'h1c : _GEN_3701;
  wire [13:0] _GEN_3703 = 14'he77 == index ? 14'h1c : _GEN_3702;
  wire [13:0] _GEN_3704 = 14'he78 == index ? 14'h1c : _GEN_3703;
  wire [13:0] _GEN_3705 = 14'he79 == index ? 14'h1c : _GEN_3704;
  wire [13:0] _GEN_3706 = 14'he7a == index ? 14'h1c : _GEN_3705;
  wire [13:0] _GEN_3707 = 14'he7b == index ? 14'h1c : _GEN_3706;
  wire [13:0] _GEN_3708 = 14'he7c == index ? 14'h1c : _GEN_3707;
  wire [13:0] _GEN_3709 = 14'he7d == index ? 14'h1c : _GEN_3708;
  wire [13:0] _GEN_3710 = 14'he7e == index ? 14'h1c : _GEN_3709;
  wire [13:0] _GEN_3711 = 14'he7f == index ? 14'h1c : _GEN_3710;
  wire [13:0] _GEN_3712 = 14'he80 == index ? 14'h0 : _GEN_3711;
  wire [13:0] _GEN_3713 = 14'he81 == index ? 14'he80 : _GEN_3712;
  wire [13:0] _GEN_3714 = 14'he82 == index ? 14'h701 : _GEN_3713;
  wire [13:0] _GEN_3715 = 14'he83 == index ? 14'h482 : _GEN_3714;
  wire [13:0] _GEN_3716 = 14'he84 == index ? 14'h381 : _GEN_3715;
  wire [13:0] _GEN_3717 = 14'he85 == index ? 14'h284 : _GEN_3716;
  wire [13:0] _GEN_3718 = 14'he86 == index ? 14'h205 : _GEN_3717;
  wire [13:0] _GEN_3719 = 14'he87 == index ? 14'h201 : _GEN_3718;
  wire [13:0] _GEN_3720 = 14'he88 == index ? 14'h185 : _GEN_3719;
  wire [13:0] _GEN_3721 = 14'he89 == index ? 14'h182 : _GEN_3720;
  wire [13:0] _GEN_3722 = 14'he8a == index ? 14'h109 : _GEN_3721;
  wire [13:0] _GEN_3723 = 14'he8b == index ? 14'h107 : _GEN_3722;
  wire [13:0] _GEN_3724 = 14'he8c == index ? 14'h105 : _GEN_3723;
  wire [13:0] _GEN_3725 = 14'he8d == index ? 14'h103 : _GEN_3724;
  wire [13:0] _GEN_3726 = 14'he8e == index ? 14'h101 : _GEN_3725;
  wire [13:0] _GEN_3727 = 14'he8f == index ? 14'h8e : _GEN_3726;
  wire [13:0] _GEN_3728 = 14'he90 == index ? 14'h8d : _GEN_3727;
  wire [13:0] _GEN_3729 = 14'he91 == index ? 14'h8c : _GEN_3728;
  wire [13:0] _GEN_3730 = 14'he92 == index ? 14'h8b : _GEN_3729;
  wire [13:0] _GEN_3731 = 14'he93 == index ? 14'h8a : _GEN_3730;
  wire [13:0] _GEN_3732 = 14'he94 == index ? 14'h89 : _GEN_3731;
  wire [13:0] _GEN_3733 = 14'he95 == index ? 14'h88 : _GEN_3732;
  wire [13:0] _GEN_3734 = 14'he96 == index ? 14'h87 : _GEN_3733;
  wire [13:0] _GEN_3735 = 14'he97 == index ? 14'h86 : _GEN_3734;
  wire [13:0] _GEN_3736 = 14'he98 == index ? 14'h85 : _GEN_3735;
  wire [13:0] _GEN_3737 = 14'he99 == index ? 14'h84 : _GEN_3736;
  wire [13:0] _GEN_3738 = 14'he9a == index ? 14'h83 : _GEN_3737;
  wire [13:0] _GEN_3739 = 14'he9b == index ? 14'h82 : _GEN_3738;
  wire [13:0] _GEN_3740 = 14'he9c == index ? 14'h81 : _GEN_3739;
  wire [13:0] _GEN_3741 = 14'he9d == index ? 14'h80 : _GEN_3740;
  wire [13:0] _GEN_3742 = 14'he9e == index ? 14'h1d : _GEN_3741;
  wire [13:0] _GEN_3743 = 14'he9f == index ? 14'h1d : _GEN_3742;
  wire [13:0] _GEN_3744 = 14'hea0 == index ? 14'h1d : _GEN_3743;
  wire [13:0] _GEN_3745 = 14'hea1 == index ? 14'h1d : _GEN_3744;
  wire [13:0] _GEN_3746 = 14'hea2 == index ? 14'h1d : _GEN_3745;
  wire [13:0] _GEN_3747 = 14'hea3 == index ? 14'h1d : _GEN_3746;
  wire [13:0] _GEN_3748 = 14'hea4 == index ? 14'h1d : _GEN_3747;
  wire [13:0] _GEN_3749 = 14'hea5 == index ? 14'h1d : _GEN_3748;
  wire [13:0] _GEN_3750 = 14'hea6 == index ? 14'h1d : _GEN_3749;
  wire [13:0] _GEN_3751 = 14'hea7 == index ? 14'h1d : _GEN_3750;
  wire [13:0] _GEN_3752 = 14'hea8 == index ? 14'h1d : _GEN_3751;
  wire [13:0] _GEN_3753 = 14'hea9 == index ? 14'h1d : _GEN_3752;
  wire [13:0] _GEN_3754 = 14'heaa == index ? 14'h1d : _GEN_3753;
  wire [13:0] _GEN_3755 = 14'heab == index ? 14'h1d : _GEN_3754;
  wire [13:0] _GEN_3756 = 14'heac == index ? 14'h1d : _GEN_3755;
  wire [13:0] _GEN_3757 = 14'head == index ? 14'h1d : _GEN_3756;
  wire [13:0] _GEN_3758 = 14'heae == index ? 14'h1d : _GEN_3757;
  wire [13:0] _GEN_3759 = 14'heaf == index ? 14'h1d : _GEN_3758;
  wire [13:0] _GEN_3760 = 14'heb0 == index ? 14'h1d : _GEN_3759;
  wire [13:0] _GEN_3761 = 14'heb1 == index ? 14'h1d : _GEN_3760;
  wire [13:0] _GEN_3762 = 14'heb2 == index ? 14'h1d : _GEN_3761;
  wire [13:0] _GEN_3763 = 14'heb3 == index ? 14'h1d : _GEN_3762;
  wire [13:0] _GEN_3764 = 14'heb4 == index ? 14'h1d : _GEN_3763;
  wire [13:0] _GEN_3765 = 14'heb5 == index ? 14'h1d : _GEN_3764;
  wire [13:0] _GEN_3766 = 14'heb6 == index ? 14'h1d : _GEN_3765;
  wire [13:0] _GEN_3767 = 14'heb7 == index ? 14'h1d : _GEN_3766;
  wire [13:0] _GEN_3768 = 14'heb8 == index ? 14'h1d : _GEN_3767;
  wire [13:0] _GEN_3769 = 14'heb9 == index ? 14'h1d : _GEN_3768;
  wire [13:0] _GEN_3770 = 14'heba == index ? 14'h1d : _GEN_3769;
  wire [13:0] _GEN_3771 = 14'hebb == index ? 14'h1d : _GEN_3770;
  wire [13:0] _GEN_3772 = 14'hebc == index ? 14'h1d : _GEN_3771;
  wire [13:0] _GEN_3773 = 14'hebd == index ? 14'h1d : _GEN_3772;
  wire [13:0] _GEN_3774 = 14'hebe == index ? 14'h1d : _GEN_3773;
  wire [13:0] _GEN_3775 = 14'hebf == index ? 14'h1d : _GEN_3774;
  wire [13:0] _GEN_3776 = 14'hec0 == index ? 14'h1d : _GEN_3775;
  wire [13:0] _GEN_3777 = 14'hec1 == index ? 14'h1d : _GEN_3776;
  wire [13:0] _GEN_3778 = 14'hec2 == index ? 14'h1d : _GEN_3777;
  wire [13:0] _GEN_3779 = 14'hec3 == index ? 14'h1d : _GEN_3778;
  wire [13:0] _GEN_3780 = 14'hec4 == index ? 14'h1d : _GEN_3779;
  wire [13:0] _GEN_3781 = 14'hec5 == index ? 14'h1d : _GEN_3780;
  wire [13:0] _GEN_3782 = 14'hec6 == index ? 14'h1d : _GEN_3781;
  wire [13:0] _GEN_3783 = 14'hec7 == index ? 14'h1d : _GEN_3782;
  wire [13:0] _GEN_3784 = 14'hec8 == index ? 14'h1d : _GEN_3783;
  wire [13:0] _GEN_3785 = 14'hec9 == index ? 14'h1d : _GEN_3784;
  wire [13:0] _GEN_3786 = 14'heca == index ? 14'h1d : _GEN_3785;
  wire [13:0] _GEN_3787 = 14'hecb == index ? 14'h1d : _GEN_3786;
  wire [13:0] _GEN_3788 = 14'hecc == index ? 14'h1d : _GEN_3787;
  wire [13:0] _GEN_3789 = 14'hecd == index ? 14'h1d : _GEN_3788;
  wire [13:0] _GEN_3790 = 14'hece == index ? 14'h1d : _GEN_3789;
  wire [13:0] _GEN_3791 = 14'hecf == index ? 14'h1d : _GEN_3790;
  wire [13:0] _GEN_3792 = 14'hed0 == index ? 14'h1d : _GEN_3791;
  wire [13:0] _GEN_3793 = 14'hed1 == index ? 14'h1d : _GEN_3792;
  wire [13:0] _GEN_3794 = 14'hed2 == index ? 14'h1d : _GEN_3793;
  wire [13:0] _GEN_3795 = 14'hed3 == index ? 14'h1d : _GEN_3794;
  wire [13:0] _GEN_3796 = 14'hed4 == index ? 14'h1d : _GEN_3795;
  wire [13:0] _GEN_3797 = 14'hed5 == index ? 14'h1d : _GEN_3796;
  wire [13:0] _GEN_3798 = 14'hed6 == index ? 14'h1d : _GEN_3797;
  wire [13:0] _GEN_3799 = 14'hed7 == index ? 14'h1d : _GEN_3798;
  wire [13:0] _GEN_3800 = 14'hed8 == index ? 14'h1d : _GEN_3799;
  wire [13:0] _GEN_3801 = 14'hed9 == index ? 14'h1d : _GEN_3800;
  wire [13:0] _GEN_3802 = 14'heda == index ? 14'h1d : _GEN_3801;
  wire [13:0] _GEN_3803 = 14'hedb == index ? 14'h1d : _GEN_3802;
  wire [13:0] _GEN_3804 = 14'hedc == index ? 14'h1d : _GEN_3803;
  wire [13:0] _GEN_3805 = 14'hedd == index ? 14'h1d : _GEN_3804;
  wire [13:0] _GEN_3806 = 14'hede == index ? 14'h1d : _GEN_3805;
  wire [13:0] _GEN_3807 = 14'hedf == index ? 14'h1d : _GEN_3806;
  wire [13:0] _GEN_3808 = 14'hee0 == index ? 14'h1d : _GEN_3807;
  wire [13:0] _GEN_3809 = 14'hee1 == index ? 14'h1d : _GEN_3808;
  wire [13:0] _GEN_3810 = 14'hee2 == index ? 14'h1d : _GEN_3809;
  wire [13:0] _GEN_3811 = 14'hee3 == index ? 14'h1d : _GEN_3810;
  wire [13:0] _GEN_3812 = 14'hee4 == index ? 14'h1d : _GEN_3811;
  wire [13:0] _GEN_3813 = 14'hee5 == index ? 14'h1d : _GEN_3812;
  wire [13:0] _GEN_3814 = 14'hee6 == index ? 14'h1d : _GEN_3813;
  wire [13:0] _GEN_3815 = 14'hee7 == index ? 14'h1d : _GEN_3814;
  wire [13:0] _GEN_3816 = 14'hee8 == index ? 14'h1d : _GEN_3815;
  wire [13:0] _GEN_3817 = 14'hee9 == index ? 14'h1d : _GEN_3816;
  wire [13:0] _GEN_3818 = 14'heea == index ? 14'h1d : _GEN_3817;
  wire [13:0] _GEN_3819 = 14'heeb == index ? 14'h1d : _GEN_3818;
  wire [13:0] _GEN_3820 = 14'heec == index ? 14'h1d : _GEN_3819;
  wire [13:0] _GEN_3821 = 14'heed == index ? 14'h1d : _GEN_3820;
  wire [13:0] _GEN_3822 = 14'heee == index ? 14'h1d : _GEN_3821;
  wire [13:0] _GEN_3823 = 14'heef == index ? 14'h1d : _GEN_3822;
  wire [13:0] _GEN_3824 = 14'hef0 == index ? 14'h1d : _GEN_3823;
  wire [13:0] _GEN_3825 = 14'hef1 == index ? 14'h1d : _GEN_3824;
  wire [13:0] _GEN_3826 = 14'hef2 == index ? 14'h1d : _GEN_3825;
  wire [13:0] _GEN_3827 = 14'hef3 == index ? 14'h1d : _GEN_3826;
  wire [13:0] _GEN_3828 = 14'hef4 == index ? 14'h1d : _GEN_3827;
  wire [13:0] _GEN_3829 = 14'hef5 == index ? 14'h1d : _GEN_3828;
  wire [13:0] _GEN_3830 = 14'hef6 == index ? 14'h1d : _GEN_3829;
  wire [13:0] _GEN_3831 = 14'hef7 == index ? 14'h1d : _GEN_3830;
  wire [13:0] _GEN_3832 = 14'hef8 == index ? 14'h1d : _GEN_3831;
  wire [13:0] _GEN_3833 = 14'hef9 == index ? 14'h1d : _GEN_3832;
  wire [13:0] _GEN_3834 = 14'hefa == index ? 14'h1d : _GEN_3833;
  wire [13:0] _GEN_3835 = 14'hefb == index ? 14'h1d : _GEN_3834;
  wire [13:0] _GEN_3836 = 14'hefc == index ? 14'h1d : _GEN_3835;
  wire [13:0] _GEN_3837 = 14'hefd == index ? 14'h1d : _GEN_3836;
  wire [13:0] _GEN_3838 = 14'hefe == index ? 14'h1d : _GEN_3837;
  wire [13:0] _GEN_3839 = 14'heff == index ? 14'h1d : _GEN_3838;
  wire [13:0] _GEN_3840 = 14'hf00 == index ? 14'h0 : _GEN_3839;
  wire [13:0] _GEN_3841 = 14'hf01 == index ? 14'hf00 : _GEN_3840;
  wire [13:0] _GEN_3842 = 14'hf02 == index ? 14'h780 : _GEN_3841;
  wire [13:0] _GEN_3843 = 14'hf03 == index ? 14'h500 : _GEN_3842;
  wire [13:0] _GEN_3844 = 14'hf04 == index ? 14'h382 : _GEN_3843;
  wire [13:0] _GEN_3845 = 14'hf05 == index ? 14'h300 : _GEN_3844;
  wire [13:0] _GEN_3846 = 14'hf06 == index ? 14'h280 : _GEN_3845;
  wire [13:0] _GEN_3847 = 14'hf07 == index ? 14'h202 : _GEN_3846;
  wire [13:0] _GEN_3848 = 14'hf08 == index ? 14'h186 : _GEN_3847;
  wire [13:0] _GEN_3849 = 14'hf09 == index ? 14'h183 : _GEN_3848;
  wire [13:0] _GEN_3850 = 14'hf0a == index ? 14'h180 : _GEN_3849;
  wire [13:0] _GEN_3851 = 14'hf0b == index ? 14'h108 : _GEN_3850;
  wire [13:0] _GEN_3852 = 14'hf0c == index ? 14'h106 : _GEN_3851;
  wire [13:0] _GEN_3853 = 14'hf0d == index ? 14'h104 : _GEN_3852;
  wire [13:0] _GEN_3854 = 14'hf0e == index ? 14'h102 : _GEN_3853;
  wire [13:0] _GEN_3855 = 14'hf0f == index ? 14'h100 : _GEN_3854;
  wire [13:0] _GEN_3856 = 14'hf10 == index ? 14'h8e : _GEN_3855;
  wire [13:0] _GEN_3857 = 14'hf11 == index ? 14'h8d : _GEN_3856;
  wire [13:0] _GEN_3858 = 14'hf12 == index ? 14'h8c : _GEN_3857;
  wire [13:0] _GEN_3859 = 14'hf13 == index ? 14'h8b : _GEN_3858;
  wire [13:0] _GEN_3860 = 14'hf14 == index ? 14'h8a : _GEN_3859;
  wire [13:0] _GEN_3861 = 14'hf15 == index ? 14'h89 : _GEN_3860;
  wire [13:0] _GEN_3862 = 14'hf16 == index ? 14'h88 : _GEN_3861;
  wire [13:0] _GEN_3863 = 14'hf17 == index ? 14'h87 : _GEN_3862;
  wire [13:0] _GEN_3864 = 14'hf18 == index ? 14'h86 : _GEN_3863;
  wire [13:0] _GEN_3865 = 14'hf19 == index ? 14'h85 : _GEN_3864;
  wire [13:0] _GEN_3866 = 14'hf1a == index ? 14'h84 : _GEN_3865;
  wire [13:0] _GEN_3867 = 14'hf1b == index ? 14'h83 : _GEN_3866;
  wire [13:0] _GEN_3868 = 14'hf1c == index ? 14'h82 : _GEN_3867;
  wire [13:0] _GEN_3869 = 14'hf1d == index ? 14'h81 : _GEN_3868;
  wire [13:0] _GEN_3870 = 14'hf1e == index ? 14'h80 : _GEN_3869;
  wire [13:0] _GEN_3871 = 14'hf1f == index ? 14'h1e : _GEN_3870;
  wire [13:0] _GEN_3872 = 14'hf20 == index ? 14'h1e : _GEN_3871;
  wire [13:0] _GEN_3873 = 14'hf21 == index ? 14'h1e : _GEN_3872;
  wire [13:0] _GEN_3874 = 14'hf22 == index ? 14'h1e : _GEN_3873;
  wire [13:0] _GEN_3875 = 14'hf23 == index ? 14'h1e : _GEN_3874;
  wire [13:0] _GEN_3876 = 14'hf24 == index ? 14'h1e : _GEN_3875;
  wire [13:0] _GEN_3877 = 14'hf25 == index ? 14'h1e : _GEN_3876;
  wire [13:0] _GEN_3878 = 14'hf26 == index ? 14'h1e : _GEN_3877;
  wire [13:0] _GEN_3879 = 14'hf27 == index ? 14'h1e : _GEN_3878;
  wire [13:0] _GEN_3880 = 14'hf28 == index ? 14'h1e : _GEN_3879;
  wire [13:0] _GEN_3881 = 14'hf29 == index ? 14'h1e : _GEN_3880;
  wire [13:0] _GEN_3882 = 14'hf2a == index ? 14'h1e : _GEN_3881;
  wire [13:0] _GEN_3883 = 14'hf2b == index ? 14'h1e : _GEN_3882;
  wire [13:0] _GEN_3884 = 14'hf2c == index ? 14'h1e : _GEN_3883;
  wire [13:0] _GEN_3885 = 14'hf2d == index ? 14'h1e : _GEN_3884;
  wire [13:0] _GEN_3886 = 14'hf2e == index ? 14'h1e : _GEN_3885;
  wire [13:0] _GEN_3887 = 14'hf2f == index ? 14'h1e : _GEN_3886;
  wire [13:0] _GEN_3888 = 14'hf30 == index ? 14'h1e : _GEN_3887;
  wire [13:0] _GEN_3889 = 14'hf31 == index ? 14'h1e : _GEN_3888;
  wire [13:0] _GEN_3890 = 14'hf32 == index ? 14'h1e : _GEN_3889;
  wire [13:0] _GEN_3891 = 14'hf33 == index ? 14'h1e : _GEN_3890;
  wire [13:0] _GEN_3892 = 14'hf34 == index ? 14'h1e : _GEN_3891;
  wire [13:0] _GEN_3893 = 14'hf35 == index ? 14'h1e : _GEN_3892;
  wire [13:0] _GEN_3894 = 14'hf36 == index ? 14'h1e : _GEN_3893;
  wire [13:0] _GEN_3895 = 14'hf37 == index ? 14'h1e : _GEN_3894;
  wire [13:0] _GEN_3896 = 14'hf38 == index ? 14'h1e : _GEN_3895;
  wire [13:0] _GEN_3897 = 14'hf39 == index ? 14'h1e : _GEN_3896;
  wire [13:0] _GEN_3898 = 14'hf3a == index ? 14'h1e : _GEN_3897;
  wire [13:0] _GEN_3899 = 14'hf3b == index ? 14'h1e : _GEN_3898;
  wire [13:0] _GEN_3900 = 14'hf3c == index ? 14'h1e : _GEN_3899;
  wire [13:0] _GEN_3901 = 14'hf3d == index ? 14'h1e : _GEN_3900;
  wire [13:0] _GEN_3902 = 14'hf3e == index ? 14'h1e : _GEN_3901;
  wire [13:0] _GEN_3903 = 14'hf3f == index ? 14'h1e : _GEN_3902;
  wire [13:0] _GEN_3904 = 14'hf40 == index ? 14'h1e : _GEN_3903;
  wire [13:0] _GEN_3905 = 14'hf41 == index ? 14'h1e : _GEN_3904;
  wire [13:0] _GEN_3906 = 14'hf42 == index ? 14'h1e : _GEN_3905;
  wire [13:0] _GEN_3907 = 14'hf43 == index ? 14'h1e : _GEN_3906;
  wire [13:0] _GEN_3908 = 14'hf44 == index ? 14'h1e : _GEN_3907;
  wire [13:0] _GEN_3909 = 14'hf45 == index ? 14'h1e : _GEN_3908;
  wire [13:0] _GEN_3910 = 14'hf46 == index ? 14'h1e : _GEN_3909;
  wire [13:0] _GEN_3911 = 14'hf47 == index ? 14'h1e : _GEN_3910;
  wire [13:0] _GEN_3912 = 14'hf48 == index ? 14'h1e : _GEN_3911;
  wire [13:0] _GEN_3913 = 14'hf49 == index ? 14'h1e : _GEN_3912;
  wire [13:0] _GEN_3914 = 14'hf4a == index ? 14'h1e : _GEN_3913;
  wire [13:0] _GEN_3915 = 14'hf4b == index ? 14'h1e : _GEN_3914;
  wire [13:0] _GEN_3916 = 14'hf4c == index ? 14'h1e : _GEN_3915;
  wire [13:0] _GEN_3917 = 14'hf4d == index ? 14'h1e : _GEN_3916;
  wire [13:0] _GEN_3918 = 14'hf4e == index ? 14'h1e : _GEN_3917;
  wire [13:0] _GEN_3919 = 14'hf4f == index ? 14'h1e : _GEN_3918;
  wire [13:0] _GEN_3920 = 14'hf50 == index ? 14'h1e : _GEN_3919;
  wire [13:0] _GEN_3921 = 14'hf51 == index ? 14'h1e : _GEN_3920;
  wire [13:0] _GEN_3922 = 14'hf52 == index ? 14'h1e : _GEN_3921;
  wire [13:0] _GEN_3923 = 14'hf53 == index ? 14'h1e : _GEN_3922;
  wire [13:0] _GEN_3924 = 14'hf54 == index ? 14'h1e : _GEN_3923;
  wire [13:0] _GEN_3925 = 14'hf55 == index ? 14'h1e : _GEN_3924;
  wire [13:0] _GEN_3926 = 14'hf56 == index ? 14'h1e : _GEN_3925;
  wire [13:0] _GEN_3927 = 14'hf57 == index ? 14'h1e : _GEN_3926;
  wire [13:0] _GEN_3928 = 14'hf58 == index ? 14'h1e : _GEN_3927;
  wire [13:0] _GEN_3929 = 14'hf59 == index ? 14'h1e : _GEN_3928;
  wire [13:0] _GEN_3930 = 14'hf5a == index ? 14'h1e : _GEN_3929;
  wire [13:0] _GEN_3931 = 14'hf5b == index ? 14'h1e : _GEN_3930;
  wire [13:0] _GEN_3932 = 14'hf5c == index ? 14'h1e : _GEN_3931;
  wire [13:0] _GEN_3933 = 14'hf5d == index ? 14'h1e : _GEN_3932;
  wire [13:0] _GEN_3934 = 14'hf5e == index ? 14'h1e : _GEN_3933;
  wire [13:0] _GEN_3935 = 14'hf5f == index ? 14'h1e : _GEN_3934;
  wire [13:0] _GEN_3936 = 14'hf60 == index ? 14'h1e : _GEN_3935;
  wire [13:0] _GEN_3937 = 14'hf61 == index ? 14'h1e : _GEN_3936;
  wire [13:0] _GEN_3938 = 14'hf62 == index ? 14'h1e : _GEN_3937;
  wire [13:0] _GEN_3939 = 14'hf63 == index ? 14'h1e : _GEN_3938;
  wire [13:0] _GEN_3940 = 14'hf64 == index ? 14'h1e : _GEN_3939;
  wire [13:0] _GEN_3941 = 14'hf65 == index ? 14'h1e : _GEN_3940;
  wire [13:0] _GEN_3942 = 14'hf66 == index ? 14'h1e : _GEN_3941;
  wire [13:0] _GEN_3943 = 14'hf67 == index ? 14'h1e : _GEN_3942;
  wire [13:0] _GEN_3944 = 14'hf68 == index ? 14'h1e : _GEN_3943;
  wire [13:0] _GEN_3945 = 14'hf69 == index ? 14'h1e : _GEN_3944;
  wire [13:0] _GEN_3946 = 14'hf6a == index ? 14'h1e : _GEN_3945;
  wire [13:0] _GEN_3947 = 14'hf6b == index ? 14'h1e : _GEN_3946;
  wire [13:0] _GEN_3948 = 14'hf6c == index ? 14'h1e : _GEN_3947;
  wire [13:0] _GEN_3949 = 14'hf6d == index ? 14'h1e : _GEN_3948;
  wire [13:0] _GEN_3950 = 14'hf6e == index ? 14'h1e : _GEN_3949;
  wire [13:0] _GEN_3951 = 14'hf6f == index ? 14'h1e : _GEN_3950;
  wire [13:0] _GEN_3952 = 14'hf70 == index ? 14'h1e : _GEN_3951;
  wire [13:0] _GEN_3953 = 14'hf71 == index ? 14'h1e : _GEN_3952;
  wire [13:0] _GEN_3954 = 14'hf72 == index ? 14'h1e : _GEN_3953;
  wire [13:0] _GEN_3955 = 14'hf73 == index ? 14'h1e : _GEN_3954;
  wire [13:0] _GEN_3956 = 14'hf74 == index ? 14'h1e : _GEN_3955;
  wire [13:0] _GEN_3957 = 14'hf75 == index ? 14'h1e : _GEN_3956;
  wire [13:0] _GEN_3958 = 14'hf76 == index ? 14'h1e : _GEN_3957;
  wire [13:0] _GEN_3959 = 14'hf77 == index ? 14'h1e : _GEN_3958;
  wire [13:0] _GEN_3960 = 14'hf78 == index ? 14'h1e : _GEN_3959;
  wire [13:0] _GEN_3961 = 14'hf79 == index ? 14'h1e : _GEN_3960;
  wire [13:0] _GEN_3962 = 14'hf7a == index ? 14'h1e : _GEN_3961;
  wire [13:0] _GEN_3963 = 14'hf7b == index ? 14'h1e : _GEN_3962;
  wire [13:0] _GEN_3964 = 14'hf7c == index ? 14'h1e : _GEN_3963;
  wire [13:0] _GEN_3965 = 14'hf7d == index ? 14'h1e : _GEN_3964;
  wire [13:0] _GEN_3966 = 14'hf7e == index ? 14'h1e : _GEN_3965;
  wire [13:0] _GEN_3967 = 14'hf7f == index ? 14'h1e : _GEN_3966;
  wire [13:0] _GEN_3968 = 14'hf80 == index ? 14'h0 : _GEN_3967;
  wire [13:0] _GEN_3969 = 14'hf81 == index ? 14'hf80 : _GEN_3968;
  wire [13:0] _GEN_3970 = 14'hf82 == index ? 14'h781 : _GEN_3969;
  wire [13:0] _GEN_3971 = 14'hf83 == index ? 14'h501 : _GEN_3970;
  wire [13:0] _GEN_3972 = 14'hf84 == index ? 14'h383 : _GEN_3971;
  wire [13:0] _GEN_3973 = 14'hf85 == index ? 14'h301 : _GEN_3972;
  wire [13:0] _GEN_3974 = 14'hf86 == index ? 14'h281 : _GEN_3973;
  wire [13:0] _GEN_3975 = 14'hf87 == index ? 14'h203 : _GEN_3974;
  wire [13:0] _GEN_3976 = 14'hf88 == index ? 14'h187 : _GEN_3975;
  wire [13:0] _GEN_3977 = 14'hf89 == index ? 14'h184 : _GEN_3976;
  wire [13:0] _GEN_3978 = 14'hf8a == index ? 14'h181 : _GEN_3977;
  wire [13:0] _GEN_3979 = 14'hf8b == index ? 14'h109 : _GEN_3978;
  wire [13:0] _GEN_3980 = 14'hf8c == index ? 14'h107 : _GEN_3979;
  wire [13:0] _GEN_3981 = 14'hf8d == index ? 14'h105 : _GEN_3980;
  wire [13:0] _GEN_3982 = 14'hf8e == index ? 14'h103 : _GEN_3981;
  wire [13:0] _GEN_3983 = 14'hf8f == index ? 14'h101 : _GEN_3982;
  wire [13:0] _GEN_3984 = 14'hf90 == index ? 14'h8f : _GEN_3983;
  wire [13:0] _GEN_3985 = 14'hf91 == index ? 14'h8e : _GEN_3984;
  wire [13:0] _GEN_3986 = 14'hf92 == index ? 14'h8d : _GEN_3985;
  wire [13:0] _GEN_3987 = 14'hf93 == index ? 14'h8c : _GEN_3986;
  wire [13:0] _GEN_3988 = 14'hf94 == index ? 14'h8b : _GEN_3987;
  wire [13:0] _GEN_3989 = 14'hf95 == index ? 14'h8a : _GEN_3988;
  wire [13:0] _GEN_3990 = 14'hf96 == index ? 14'h89 : _GEN_3989;
  wire [13:0] _GEN_3991 = 14'hf97 == index ? 14'h88 : _GEN_3990;
  wire [13:0] _GEN_3992 = 14'hf98 == index ? 14'h87 : _GEN_3991;
  wire [13:0] _GEN_3993 = 14'hf99 == index ? 14'h86 : _GEN_3992;
  wire [13:0] _GEN_3994 = 14'hf9a == index ? 14'h85 : _GEN_3993;
  wire [13:0] _GEN_3995 = 14'hf9b == index ? 14'h84 : _GEN_3994;
  wire [13:0] _GEN_3996 = 14'hf9c == index ? 14'h83 : _GEN_3995;
  wire [13:0] _GEN_3997 = 14'hf9d == index ? 14'h82 : _GEN_3996;
  wire [13:0] _GEN_3998 = 14'hf9e == index ? 14'h81 : _GEN_3997;
  wire [13:0] _GEN_3999 = 14'hf9f == index ? 14'h80 : _GEN_3998;
  wire [13:0] _GEN_4000 = 14'hfa0 == index ? 14'h1f : _GEN_3999;
  wire [13:0] _GEN_4001 = 14'hfa1 == index ? 14'h1f : _GEN_4000;
  wire [13:0] _GEN_4002 = 14'hfa2 == index ? 14'h1f : _GEN_4001;
  wire [13:0] _GEN_4003 = 14'hfa3 == index ? 14'h1f : _GEN_4002;
  wire [13:0] _GEN_4004 = 14'hfa4 == index ? 14'h1f : _GEN_4003;
  wire [13:0] _GEN_4005 = 14'hfa5 == index ? 14'h1f : _GEN_4004;
  wire [13:0] _GEN_4006 = 14'hfa6 == index ? 14'h1f : _GEN_4005;
  wire [13:0] _GEN_4007 = 14'hfa7 == index ? 14'h1f : _GEN_4006;
  wire [13:0] _GEN_4008 = 14'hfa8 == index ? 14'h1f : _GEN_4007;
  wire [13:0] _GEN_4009 = 14'hfa9 == index ? 14'h1f : _GEN_4008;
  wire [13:0] _GEN_4010 = 14'hfaa == index ? 14'h1f : _GEN_4009;
  wire [13:0] _GEN_4011 = 14'hfab == index ? 14'h1f : _GEN_4010;
  wire [13:0] _GEN_4012 = 14'hfac == index ? 14'h1f : _GEN_4011;
  wire [13:0] _GEN_4013 = 14'hfad == index ? 14'h1f : _GEN_4012;
  wire [13:0] _GEN_4014 = 14'hfae == index ? 14'h1f : _GEN_4013;
  wire [13:0] _GEN_4015 = 14'hfaf == index ? 14'h1f : _GEN_4014;
  wire [13:0] _GEN_4016 = 14'hfb0 == index ? 14'h1f : _GEN_4015;
  wire [13:0] _GEN_4017 = 14'hfb1 == index ? 14'h1f : _GEN_4016;
  wire [13:0] _GEN_4018 = 14'hfb2 == index ? 14'h1f : _GEN_4017;
  wire [13:0] _GEN_4019 = 14'hfb3 == index ? 14'h1f : _GEN_4018;
  wire [13:0] _GEN_4020 = 14'hfb4 == index ? 14'h1f : _GEN_4019;
  wire [13:0] _GEN_4021 = 14'hfb5 == index ? 14'h1f : _GEN_4020;
  wire [13:0] _GEN_4022 = 14'hfb6 == index ? 14'h1f : _GEN_4021;
  wire [13:0] _GEN_4023 = 14'hfb7 == index ? 14'h1f : _GEN_4022;
  wire [13:0] _GEN_4024 = 14'hfb8 == index ? 14'h1f : _GEN_4023;
  wire [13:0] _GEN_4025 = 14'hfb9 == index ? 14'h1f : _GEN_4024;
  wire [13:0] _GEN_4026 = 14'hfba == index ? 14'h1f : _GEN_4025;
  wire [13:0] _GEN_4027 = 14'hfbb == index ? 14'h1f : _GEN_4026;
  wire [13:0] _GEN_4028 = 14'hfbc == index ? 14'h1f : _GEN_4027;
  wire [13:0] _GEN_4029 = 14'hfbd == index ? 14'h1f : _GEN_4028;
  wire [13:0] _GEN_4030 = 14'hfbe == index ? 14'h1f : _GEN_4029;
  wire [13:0] _GEN_4031 = 14'hfbf == index ? 14'h1f : _GEN_4030;
  wire [13:0] _GEN_4032 = 14'hfc0 == index ? 14'h1f : _GEN_4031;
  wire [13:0] _GEN_4033 = 14'hfc1 == index ? 14'h1f : _GEN_4032;
  wire [13:0] _GEN_4034 = 14'hfc2 == index ? 14'h1f : _GEN_4033;
  wire [13:0] _GEN_4035 = 14'hfc3 == index ? 14'h1f : _GEN_4034;
  wire [13:0] _GEN_4036 = 14'hfc4 == index ? 14'h1f : _GEN_4035;
  wire [13:0] _GEN_4037 = 14'hfc5 == index ? 14'h1f : _GEN_4036;
  wire [13:0] _GEN_4038 = 14'hfc6 == index ? 14'h1f : _GEN_4037;
  wire [13:0] _GEN_4039 = 14'hfc7 == index ? 14'h1f : _GEN_4038;
  wire [13:0] _GEN_4040 = 14'hfc8 == index ? 14'h1f : _GEN_4039;
  wire [13:0] _GEN_4041 = 14'hfc9 == index ? 14'h1f : _GEN_4040;
  wire [13:0] _GEN_4042 = 14'hfca == index ? 14'h1f : _GEN_4041;
  wire [13:0] _GEN_4043 = 14'hfcb == index ? 14'h1f : _GEN_4042;
  wire [13:0] _GEN_4044 = 14'hfcc == index ? 14'h1f : _GEN_4043;
  wire [13:0] _GEN_4045 = 14'hfcd == index ? 14'h1f : _GEN_4044;
  wire [13:0] _GEN_4046 = 14'hfce == index ? 14'h1f : _GEN_4045;
  wire [13:0] _GEN_4047 = 14'hfcf == index ? 14'h1f : _GEN_4046;
  wire [13:0] _GEN_4048 = 14'hfd0 == index ? 14'h1f : _GEN_4047;
  wire [13:0] _GEN_4049 = 14'hfd1 == index ? 14'h1f : _GEN_4048;
  wire [13:0] _GEN_4050 = 14'hfd2 == index ? 14'h1f : _GEN_4049;
  wire [13:0] _GEN_4051 = 14'hfd3 == index ? 14'h1f : _GEN_4050;
  wire [13:0] _GEN_4052 = 14'hfd4 == index ? 14'h1f : _GEN_4051;
  wire [13:0] _GEN_4053 = 14'hfd5 == index ? 14'h1f : _GEN_4052;
  wire [13:0] _GEN_4054 = 14'hfd6 == index ? 14'h1f : _GEN_4053;
  wire [13:0] _GEN_4055 = 14'hfd7 == index ? 14'h1f : _GEN_4054;
  wire [13:0] _GEN_4056 = 14'hfd8 == index ? 14'h1f : _GEN_4055;
  wire [13:0] _GEN_4057 = 14'hfd9 == index ? 14'h1f : _GEN_4056;
  wire [13:0] _GEN_4058 = 14'hfda == index ? 14'h1f : _GEN_4057;
  wire [13:0] _GEN_4059 = 14'hfdb == index ? 14'h1f : _GEN_4058;
  wire [13:0] _GEN_4060 = 14'hfdc == index ? 14'h1f : _GEN_4059;
  wire [13:0] _GEN_4061 = 14'hfdd == index ? 14'h1f : _GEN_4060;
  wire [13:0] _GEN_4062 = 14'hfde == index ? 14'h1f : _GEN_4061;
  wire [13:0] _GEN_4063 = 14'hfdf == index ? 14'h1f : _GEN_4062;
  wire [13:0] _GEN_4064 = 14'hfe0 == index ? 14'h1f : _GEN_4063;
  wire [13:0] _GEN_4065 = 14'hfe1 == index ? 14'h1f : _GEN_4064;
  wire [13:0] _GEN_4066 = 14'hfe2 == index ? 14'h1f : _GEN_4065;
  wire [13:0] _GEN_4067 = 14'hfe3 == index ? 14'h1f : _GEN_4066;
  wire [13:0] _GEN_4068 = 14'hfe4 == index ? 14'h1f : _GEN_4067;
  wire [13:0] _GEN_4069 = 14'hfe5 == index ? 14'h1f : _GEN_4068;
  wire [13:0] _GEN_4070 = 14'hfe6 == index ? 14'h1f : _GEN_4069;
  wire [13:0] _GEN_4071 = 14'hfe7 == index ? 14'h1f : _GEN_4070;
  wire [13:0] _GEN_4072 = 14'hfe8 == index ? 14'h1f : _GEN_4071;
  wire [13:0] _GEN_4073 = 14'hfe9 == index ? 14'h1f : _GEN_4072;
  wire [13:0] _GEN_4074 = 14'hfea == index ? 14'h1f : _GEN_4073;
  wire [13:0] _GEN_4075 = 14'hfeb == index ? 14'h1f : _GEN_4074;
  wire [13:0] _GEN_4076 = 14'hfec == index ? 14'h1f : _GEN_4075;
  wire [13:0] _GEN_4077 = 14'hfed == index ? 14'h1f : _GEN_4076;
  wire [13:0] _GEN_4078 = 14'hfee == index ? 14'h1f : _GEN_4077;
  wire [13:0] _GEN_4079 = 14'hfef == index ? 14'h1f : _GEN_4078;
  wire [13:0] _GEN_4080 = 14'hff0 == index ? 14'h1f : _GEN_4079;
  wire [13:0] _GEN_4081 = 14'hff1 == index ? 14'h1f : _GEN_4080;
  wire [13:0] _GEN_4082 = 14'hff2 == index ? 14'h1f : _GEN_4081;
  wire [13:0] _GEN_4083 = 14'hff3 == index ? 14'h1f : _GEN_4082;
  wire [13:0] _GEN_4084 = 14'hff4 == index ? 14'h1f : _GEN_4083;
  wire [13:0] _GEN_4085 = 14'hff5 == index ? 14'h1f : _GEN_4084;
  wire [13:0] _GEN_4086 = 14'hff6 == index ? 14'h1f : _GEN_4085;
  wire [13:0] _GEN_4087 = 14'hff7 == index ? 14'h1f : _GEN_4086;
  wire [13:0] _GEN_4088 = 14'hff8 == index ? 14'h1f : _GEN_4087;
  wire [13:0] _GEN_4089 = 14'hff9 == index ? 14'h1f : _GEN_4088;
  wire [13:0] _GEN_4090 = 14'hffa == index ? 14'h1f : _GEN_4089;
  wire [13:0] _GEN_4091 = 14'hffb == index ? 14'h1f : _GEN_4090;
  wire [13:0] _GEN_4092 = 14'hffc == index ? 14'h1f : _GEN_4091;
  wire [13:0] _GEN_4093 = 14'hffd == index ? 14'h1f : _GEN_4092;
  wire [13:0] _GEN_4094 = 14'hffe == index ? 14'h1f : _GEN_4093;
  wire [13:0] _GEN_4095 = 14'hfff == index ? 14'h1f : _GEN_4094;
  wire [13:0] _GEN_4096 = 14'h1000 == index ? 14'h0 : _GEN_4095;
  wire [13:0] _GEN_4097 = 14'h1001 == index ? 14'h1000 : _GEN_4096;
  wire [13:0] _GEN_4098 = 14'h1002 == index ? 14'h800 : _GEN_4097;
  wire [13:0] _GEN_4099 = 14'h1003 == index ? 14'h502 : _GEN_4098;
  wire [13:0] _GEN_4100 = 14'h1004 == index ? 14'h400 : _GEN_4099;
  wire [13:0] _GEN_4101 = 14'h1005 == index ? 14'h302 : _GEN_4100;
  wire [13:0] _GEN_4102 = 14'h1006 == index ? 14'h282 : _GEN_4101;
  wire [13:0] _GEN_4103 = 14'h1007 == index ? 14'h204 : _GEN_4102;
  wire [13:0] _GEN_4104 = 14'h1008 == index ? 14'h200 : _GEN_4103;
  wire [13:0] _GEN_4105 = 14'h1009 == index ? 14'h185 : _GEN_4104;
  wire [13:0] _GEN_4106 = 14'h100a == index ? 14'h182 : _GEN_4105;
  wire [13:0] _GEN_4107 = 14'h100b == index ? 14'h10a : _GEN_4106;
  wire [13:0] _GEN_4108 = 14'h100c == index ? 14'h108 : _GEN_4107;
  wire [13:0] _GEN_4109 = 14'h100d == index ? 14'h106 : _GEN_4108;
  wire [13:0] _GEN_4110 = 14'h100e == index ? 14'h104 : _GEN_4109;
  wire [13:0] _GEN_4111 = 14'h100f == index ? 14'h102 : _GEN_4110;
  wire [13:0] _GEN_4112 = 14'h1010 == index ? 14'h100 : _GEN_4111;
  wire [13:0] _GEN_4113 = 14'h1011 == index ? 14'h8f : _GEN_4112;
  wire [13:0] _GEN_4114 = 14'h1012 == index ? 14'h8e : _GEN_4113;
  wire [13:0] _GEN_4115 = 14'h1013 == index ? 14'h8d : _GEN_4114;
  wire [13:0] _GEN_4116 = 14'h1014 == index ? 14'h8c : _GEN_4115;
  wire [13:0] _GEN_4117 = 14'h1015 == index ? 14'h8b : _GEN_4116;
  wire [13:0] _GEN_4118 = 14'h1016 == index ? 14'h8a : _GEN_4117;
  wire [13:0] _GEN_4119 = 14'h1017 == index ? 14'h89 : _GEN_4118;
  wire [13:0] _GEN_4120 = 14'h1018 == index ? 14'h88 : _GEN_4119;
  wire [13:0] _GEN_4121 = 14'h1019 == index ? 14'h87 : _GEN_4120;
  wire [13:0] _GEN_4122 = 14'h101a == index ? 14'h86 : _GEN_4121;
  wire [13:0] _GEN_4123 = 14'h101b == index ? 14'h85 : _GEN_4122;
  wire [13:0] _GEN_4124 = 14'h101c == index ? 14'h84 : _GEN_4123;
  wire [13:0] _GEN_4125 = 14'h101d == index ? 14'h83 : _GEN_4124;
  wire [13:0] _GEN_4126 = 14'h101e == index ? 14'h82 : _GEN_4125;
  wire [13:0] _GEN_4127 = 14'h101f == index ? 14'h81 : _GEN_4126;
  wire [13:0] _GEN_4128 = 14'h1020 == index ? 14'h80 : _GEN_4127;
  wire [13:0] _GEN_4129 = 14'h1021 == index ? 14'h20 : _GEN_4128;
  wire [13:0] _GEN_4130 = 14'h1022 == index ? 14'h20 : _GEN_4129;
  wire [13:0] _GEN_4131 = 14'h1023 == index ? 14'h20 : _GEN_4130;
  wire [13:0] _GEN_4132 = 14'h1024 == index ? 14'h20 : _GEN_4131;
  wire [13:0] _GEN_4133 = 14'h1025 == index ? 14'h20 : _GEN_4132;
  wire [13:0] _GEN_4134 = 14'h1026 == index ? 14'h20 : _GEN_4133;
  wire [13:0] _GEN_4135 = 14'h1027 == index ? 14'h20 : _GEN_4134;
  wire [13:0] _GEN_4136 = 14'h1028 == index ? 14'h20 : _GEN_4135;
  wire [13:0] _GEN_4137 = 14'h1029 == index ? 14'h20 : _GEN_4136;
  wire [13:0] _GEN_4138 = 14'h102a == index ? 14'h20 : _GEN_4137;
  wire [13:0] _GEN_4139 = 14'h102b == index ? 14'h20 : _GEN_4138;
  wire [13:0] _GEN_4140 = 14'h102c == index ? 14'h20 : _GEN_4139;
  wire [13:0] _GEN_4141 = 14'h102d == index ? 14'h20 : _GEN_4140;
  wire [13:0] _GEN_4142 = 14'h102e == index ? 14'h20 : _GEN_4141;
  wire [13:0] _GEN_4143 = 14'h102f == index ? 14'h20 : _GEN_4142;
  wire [13:0] _GEN_4144 = 14'h1030 == index ? 14'h20 : _GEN_4143;
  wire [13:0] _GEN_4145 = 14'h1031 == index ? 14'h20 : _GEN_4144;
  wire [13:0] _GEN_4146 = 14'h1032 == index ? 14'h20 : _GEN_4145;
  wire [13:0] _GEN_4147 = 14'h1033 == index ? 14'h20 : _GEN_4146;
  wire [13:0] _GEN_4148 = 14'h1034 == index ? 14'h20 : _GEN_4147;
  wire [13:0] _GEN_4149 = 14'h1035 == index ? 14'h20 : _GEN_4148;
  wire [13:0] _GEN_4150 = 14'h1036 == index ? 14'h20 : _GEN_4149;
  wire [13:0] _GEN_4151 = 14'h1037 == index ? 14'h20 : _GEN_4150;
  wire [13:0] _GEN_4152 = 14'h1038 == index ? 14'h20 : _GEN_4151;
  wire [13:0] _GEN_4153 = 14'h1039 == index ? 14'h20 : _GEN_4152;
  wire [13:0] _GEN_4154 = 14'h103a == index ? 14'h20 : _GEN_4153;
  wire [13:0] _GEN_4155 = 14'h103b == index ? 14'h20 : _GEN_4154;
  wire [13:0] _GEN_4156 = 14'h103c == index ? 14'h20 : _GEN_4155;
  wire [13:0] _GEN_4157 = 14'h103d == index ? 14'h20 : _GEN_4156;
  wire [13:0] _GEN_4158 = 14'h103e == index ? 14'h20 : _GEN_4157;
  wire [13:0] _GEN_4159 = 14'h103f == index ? 14'h20 : _GEN_4158;
  wire [13:0] _GEN_4160 = 14'h1040 == index ? 14'h20 : _GEN_4159;
  wire [13:0] _GEN_4161 = 14'h1041 == index ? 14'h20 : _GEN_4160;
  wire [13:0] _GEN_4162 = 14'h1042 == index ? 14'h20 : _GEN_4161;
  wire [13:0] _GEN_4163 = 14'h1043 == index ? 14'h20 : _GEN_4162;
  wire [13:0] _GEN_4164 = 14'h1044 == index ? 14'h20 : _GEN_4163;
  wire [13:0] _GEN_4165 = 14'h1045 == index ? 14'h20 : _GEN_4164;
  wire [13:0] _GEN_4166 = 14'h1046 == index ? 14'h20 : _GEN_4165;
  wire [13:0] _GEN_4167 = 14'h1047 == index ? 14'h20 : _GEN_4166;
  wire [13:0] _GEN_4168 = 14'h1048 == index ? 14'h20 : _GEN_4167;
  wire [13:0] _GEN_4169 = 14'h1049 == index ? 14'h20 : _GEN_4168;
  wire [13:0] _GEN_4170 = 14'h104a == index ? 14'h20 : _GEN_4169;
  wire [13:0] _GEN_4171 = 14'h104b == index ? 14'h20 : _GEN_4170;
  wire [13:0] _GEN_4172 = 14'h104c == index ? 14'h20 : _GEN_4171;
  wire [13:0] _GEN_4173 = 14'h104d == index ? 14'h20 : _GEN_4172;
  wire [13:0] _GEN_4174 = 14'h104e == index ? 14'h20 : _GEN_4173;
  wire [13:0] _GEN_4175 = 14'h104f == index ? 14'h20 : _GEN_4174;
  wire [13:0] _GEN_4176 = 14'h1050 == index ? 14'h20 : _GEN_4175;
  wire [13:0] _GEN_4177 = 14'h1051 == index ? 14'h20 : _GEN_4176;
  wire [13:0] _GEN_4178 = 14'h1052 == index ? 14'h20 : _GEN_4177;
  wire [13:0] _GEN_4179 = 14'h1053 == index ? 14'h20 : _GEN_4178;
  wire [13:0] _GEN_4180 = 14'h1054 == index ? 14'h20 : _GEN_4179;
  wire [13:0] _GEN_4181 = 14'h1055 == index ? 14'h20 : _GEN_4180;
  wire [13:0] _GEN_4182 = 14'h1056 == index ? 14'h20 : _GEN_4181;
  wire [13:0] _GEN_4183 = 14'h1057 == index ? 14'h20 : _GEN_4182;
  wire [13:0] _GEN_4184 = 14'h1058 == index ? 14'h20 : _GEN_4183;
  wire [13:0] _GEN_4185 = 14'h1059 == index ? 14'h20 : _GEN_4184;
  wire [13:0] _GEN_4186 = 14'h105a == index ? 14'h20 : _GEN_4185;
  wire [13:0] _GEN_4187 = 14'h105b == index ? 14'h20 : _GEN_4186;
  wire [13:0] _GEN_4188 = 14'h105c == index ? 14'h20 : _GEN_4187;
  wire [13:0] _GEN_4189 = 14'h105d == index ? 14'h20 : _GEN_4188;
  wire [13:0] _GEN_4190 = 14'h105e == index ? 14'h20 : _GEN_4189;
  wire [13:0] _GEN_4191 = 14'h105f == index ? 14'h20 : _GEN_4190;
  wire [13:0] _GEN_4192 = 14'h1060 == index ? 14'h20 : _GEN_4191;
  wire [13:0] _GEN_4193 = 14'h1061 == index ? 14'h20 : _GEN_4192;
  wire [13:0] _GEN_4194 = 14'h1062 == index ? 14'h20 : _GEN_4193;
  wire [13:0] _GEN_4195 = 14'h1063 == index ? 14'h20 : _GEN_4194;
  wire [13:0] _GEN_4196 = 14'h1064 == index ? 14'h20 : _GEN_4195;
  wire [13:0] _GEN_4197 = 14'h1065 == index ? 14'h20 : _GEN_4196;
  wire [13:0] _GEN_4198 = 14'h1066 == index ? 14'h20 : _GEN_4197;
  wire [13:0] _GEN_4199 = 14'h1067 == index ? 14'h20 : _GEN_4198;
  wire [13:0] _GEN_4200 = 14'h1068 == index ? 14'h20 : _GEN_4199;
  wire [13:0] _GEN_4201 = 14'h1069 == index ? 14'h20 : _GEN_4200;
  wire [13:0] _GEN_4202 = 14'h106a == index ? 14'h20 : _GEN_4201;
  wire [13:0] _GEN_4203 = 14'h106b == index ? 14'h20 : _GEN_4202;
  wire [13:0] _GEN_4204 = 14'h106c == index ? 14'h20 : _GEN_4203;
  wire [13:0] _GEN_4205 = 14'h106d == index ? 14'h20 : _GEN_4204;
  wire [13:0] _GEN_4206 = 14'h106e == index ? 14'h20 : _GEN_4205;
  wire [13:0] _GEN_4207 = 14'h106f == index ? 14'h20 : _GEN_4206;
  wire [13:0] _GEN_4208 = 14'h1070 == index ? 14'h20 : _GEN_4207;
  wire [13:0] _GEN_4209 = 14'h1071 == index ? 14'h20 : _GEN_4208;
  wire [13:0] _GEN_4210 = 14'h1072 == index ? 14'h20 : _GEN_4209;
  wire [13:0] _GEN_4211 = 14'h1073 == index ? 14'h20 : _GEN_4210;
  wire [13:0] _GEN_4212 = 14'h1074 == index ? 14'h20 : _GEN_4211;
  wire [13:0] _GEN_4213 = 14'h1075 == index ? 14'h20 : _GEN_4212;
  wire [13:0] _GEN_4214 = 14'h1076 == index ? 14'h20 : _GEN_4213;
  wire [13:0] _GEN_4215 = 14'h1077 == index ? 14'h20 : _GEN_4214;
  wire [13:0] _GEN_4216 = 14'h1078 == index ? 14'h20 : _GEN_4215;
  wire [13:0] _GEN_4217 = 14'h1079 == index ? 14'h20 : _GEN_4216;
  wire [13:0] _GEN_4218 = 14'h107a == index ? 14'h20 : _GEN_4217;
  wire [13:0] _GEN_4219 = 14'h107b == index ? 14'h20 : _GEN_4218;
  wire [13:0] _GEN_4220 = 14'h107c == index ? 14'h20 : _GEN_4219;
  wire [13:0] _GEN_4221 = 14'h107d == index ? 14'h20 : _GEN_4220;
  wire [13:0] _GEN_4222 = 14'h107e == index ? 14'h20 : _GEN_4221;
  wire [13:0] _GEN_4223 = 14'h107f == index ? 14'h20 : _GEN_4222;
  wire [13:0] _GEN_4224 = 14'h1080 == index ? 14'h0 : _GEN_4223;
  wire [13:0] _GEN_4225 = 14'h1081 == index ? 14'h1080 : _GEN_4224;
  wire [13:0] _GEN_4226 = 14'h1082 == index ? 14'h801 : _GEN_4225;
  wire [13:0] _GEN_4227 = 14'h1083 == index ? 14'h580 : _GEN_4226;
  wire [13:0] _GEN_4228 = 14'h1084 == index ? 14'h401 : _GEN_4227;
  wire [13:0] _GEN_4229 = 14'h1085 == index ? 14'h303 : _GEN_4228;
  wire [13:0] _GEN_4230 = 14'h1086 == index ? 14'h283 : _GEN_4229;
  wire [13:0] _GEN_4231 = 14'h1087 == index ? 14'h205 : _GEN_4230;
  wire [13:0] _GEN_4232 = 14'h1088 == index ? 14'h201 : _GEN_4231;
  wire [13:0] _GEN_4233 = 14'h1089 == index ? 14'h186 : _GEN_4232;
  wire [13:0] _GEN_4234 = 14'h108a == index ? 14'h183 : _GEN_4233;
  wire [13:0] _GEN_4235 = 14'h108b == index ? 14'h180 : _GEN_4234;
  wire [13:0] _GEN_4236 = 14'h108c == index ? 14'h109 : _GEN_4235;
  wire [13:0] _GEN_4237 = 14'h108d == index ? 14'h107 : _GEN_4236;
  wire [13:0] _GEN_4238 = 14'h108e == index ? 14'h105 : _GEN_4237;
  wire [13:0] _GEN_4239 = 14'h108f == index ? 14'h103 : _GEN_4238;
  wire [13:0] _GEN_4240 = 14'h1090 == index ? 14'h101 : _GEN_4239;
  wire [13:0] _GEN_4241 = 14'h1091 == index ? 14'h90 : _GEN_4240;
  wire [13:0] _GEN_4242 = 14'h1092 == index ? 14'h8f : _GEN_4241;
  wire [13:0] _GEN_4243 = 14'h1093 == index ? 14'h8e : _GEN_4242;
  wire [13:0] _GEN_4244 = 14'h1094 == index ? 14'h8d : _GEN_4243;
  wire [13:0] _GEN_4245 = 14'h1095 == index ? 14'h8c : _GEN_4244;
  wire [13:0] _GEN_4246 = 14'h1096 == index ? 14'h8b : _GEN_4245;
  wire [13:0] _GEN_4247 = 14'h1097 == index ? 14'h8a : _GEN_4246;
  wire [13:0] _GEN_4248 = 14'h1098 == index ? 14'h89 : _GEN_4247;
  wire [13:0] _GEN_4249 = 14'h1099 == index ? 14'h88 : _GEN_4248;
  wire [13:0] _GEN_4250 = 14'h109a == index ? 14'h87 : _GEN_4249;
  wire [13:0] _GEN_4251 = 14'h109b == index ? 14'h86 : _GEN_4250;
  wire [13:0] _GEN_4252 = 14'h109c == index ? 14'h85 : _GEN_4251;
  wire [13:0] _GEN_4253 = 14'h109d == index ? 14'h84 : _GEN_4252;
  wire [13:0] _GEN_4254 = 14'h109e == index ? 14'h83 : _GEN_4253;
  wire [13:0] _GEN_4255 = 14'h109f == index ? 14'h82 : _GEN_4254;
  wire [13:0] _GEN_4256 = 14'h10a0 == index ? 14'h81 : _GEN_4255;
  wire [13:0] _GEN_4257 = 14'h10a1 == index ? 14'h80 : _GEN_4256;
  wire [13:0] _GEN_4258 = 14'h10a2 == index ? 14'h21 : _GEN_4257;
  wire [13:0] _GEN_4259 = 14'h10a3 == index ? 14'h21 : _GEN_4258;
  wire [13:0] _GEN_4260 = 14'h10a4 == index ? 14'h21 : _GEN_4259;
  wire [13:0] _GEN_4261 = 14'h10a5 == index ? 14'h21 : _GEN_4260;
  wire [13:0] _GEN_4262 = 14'h10a6 == index ? 14'h21 : _GEN_4261;
  wire [13:0] _GEN_4263 = 14'h10a7 == index ? 14'h21 : _GEN_4262;
  wire [13:0] _GEN_4264 = 14'h10a8 == index ? 14'h21 : _GEN_4263;
  wire [13:0] _GEN_4265 = 14'h10a9 == index ? 14'h21 : _GEN_4264;
  wire [13:0] _GEN_4266 = 14'h10aa == index ? 14'h21 : _GEN_4265;
  wire [13:0] _GEN_4267 = 14'h10ab == index ? 14'h21 : _GEN_4266;
  wire [13:0] _GEN_4268 = 14'h10ac == index ? 14'h21 : _GEN_4267;
  wire [13:0] _GEN_4269 = 14'h10ad == index ? 14'h21 : _GEN_4268;
  wire [13:0] _GEN_4270 = 14'h10ae == index ? 14'h21 : _GEN_4269;
  wire [13:0] _GEN_4271 = 14'h10af == index ? 14'h21 : _GEN_4270;
  wire [13:0] _GEN_4272 = 14'h10b0 == index ? 14'h21 : _GEN_4271;
  wire [13:0] _GEN_4273 = 14'h10b1 == index ? 14'h21 : _GEN_4272;
  wire [13:0] _GEN_4274 = 14'h10b2 == index ? 14'h21 : _GEN_4273;
  wire [13:0] _GEN_4275 = 14'h10b3 == index ? 14'h21 : _GEN_4274;
  wire [13:0] _GEN_4276 = 14'h10b4 == index ? 14'h21 : _GEN_4275;
  wire [13:0] _GEN_4277 = 14'h10b5 == index ? 14'h21 : _GEN_4276;
  wire [13:0] _GEN_4278 = 14'h10b6 == index ? 14'h21 : _GEN_4277;
  wire [13:0] _GEN_4279 = 14'h10b7 == index ? 14'h21 : _GEN_4278;
  wire [13:0] _GEN_4280 = 14'h10b8 == index ? 14'h21 : _GEN_4279;
  wire [13:0] _GEN_4281 = 14'h10b9 == index ? 14'h21 : _GEN_4280;
  wire [13:0] _GEN_4282 = 14'h10ba == index ? 14'h21 : _GEN_4281;
  wire [13:0] _GEN_4283 = 14'h10bb == index ? 14'h21 : _GEN_4282;
  wire [13:0] _GEN_4284 = 14'h10bc == index ? 14'h21 : _GEN_4283;
  wire [13:0] _GEN_4285 = 14'h10bd == index ? 14'h21 : _GEN_4284;
  wire [13:0] _GEN_4286 = 14'h10be == index ? 14'h21 : _GEN_4285;
  wire [13:0] _GEN_4287 = 14'h10bf == index ? 14'h21 : _GEN_4286;
  wire [13:0] _GEN_4288 = 14'h10c0 == index ? 14'h21 : _GEN_4287;
  wire [13:0] _GEN_4289 = 14'h10c1 == index ? 14'h21 : _GEN_4288;
  wire [13:0] _GEN_4290 = 14'h10c2 == index ? 14'h21 : _GEN_4289;
  wire [13:0] _GEN_4291 = 14'h10c3 == index ? 14'h21 : _GEN_4290;
  wire [13:0] _GEN_4292 = 14'h10c4 == index ? 14'h21 : _GEN_4291;
  wire [13:0] _GEN_4293 = 14'h10c5 == index ? 14'h21 : _GEN_4292;
  wire [13:0] _GEN_4294 = 14'h10c6 == index ? 14'h21 : _GEN_4293;
  wire [13:0] _GEN_4295 = 14'h10c7 == index ? 14'h21 : _GEN_4294;
  wire [13:0] _GEN_4296 = 14'h10c8 == index ? 14'h21 : _GEN_4295;
  wire [13:0] _GEN_4297 = 14'h10c9 == index ? 14'h21 : _GEN_4296;
  wire [13:0] _GEN_4298 = 14'h10ca == index ? 14'h21 : _GEN_4297;
  wire [13:0] _GEN_4299 = 14'h10cb == index ? 14'h21 : _GEN_4298;
  wire [13:0] _GEN_4300 = 14'h10cc == index ? 14'h21 : _GEN_4299;
  wire [13:0] _GEN_4301 = 14'h10cd == index ? 14'h21 : _GEN_4300;
  wire [13:0] _GEN_4302 = 14'h10ce == index ? 14'h21 : _GEN_4301;
  wire [13:0] _GEN_4303 = 14'h10cf == index ? 14'h21 : _GEN_4302;
  wire [13:0] _GEN_4304 = 14'h10d0 == index ? 14'h21 : _GEN_4303;
  wire [13:0] _GEN_4305 = 14'h10d1 == index ? 14'h21 : _GEN_4304;
  wire [13:0] _GEN_4306 = 14'h10d2 == index ? 14'h21 : _GEN_4305;
  wire [13:0] _GEN_4307 = 14'h10d3 == index ? 14'h21 : _GEN_4306;
  wire [13:0] _GEN_4308 = 14'h10d4 == index ? 14'h21 : _GEN_4307;
  wire [13:0] _GEN_4309 = 14'h10d5 == index ? 14'h21 : _GEN_4308;
  wire [13:0] _GEN_4310 = 14'h10d6 == index ? 14'h21 : _GEN_4309;
  wire [13:0] _GEN_4311 = 14'h10d7 == index ? 14'h21 : _GEN_4310;
  wire [13:0] _GEN_4312 = 14'h10d8 == index ? 14'h21 : _GEN_4311;
  wire [13:0] _GEN_4313 = 14'h10d9 == index ? 14'h21 : _GEN_4312;
  wire [13:0] _GEN_4314 = 14'h10da == index ? 14'h21 : _GEN_4313;
  wire [13:0] _GEN_4315 = 14'h10db == index ? 14'h21 : _GEN_4314;
  wire [13:0] _GEN_4316 = 14'h10dc == index ? 14'h21 : _GEN_4315;
  wire [13:0] _GEN_4317 = 14'h10dd == index ? 14'h21 : _GEN_4316;
  wire [13:0] _GEN_4318 = 14'h10de == index ? 14'h21 : _GEN_4317;
  wire [13:0] _GEN_4319 = 14'h10df == index ? 14'h21 : _GEN_4318;
  wire [13:0] _GEN_4320 = 14'h10e0 == index ? 14'h21 : _GEN_4319;
  wire [13:0] _GEN_4321 = 14'h10e1 == index ? 14'h21 : _GEN_4320;
  wire [13:0] _GEN_4322 = 14'h10e2 == index ? 14'h21 : _GEN_4321;
  wire [13:0] _GEN_4323 = 14'h10e3 == index ? 14'h21 : _GEN_4322;
  wire [13:0] _GEN_4324 = 14'h10e4 == index ? 14'h21 : _GEN_4323;
  wire [13:0] _GEN_4325 = 14'h10e5 == index ? 14'h21 : _GEN_4324;
  wire [13:0] _GEN_4326 = 14'h10e6 == index ? 14'h21 : _GEN_4325;
  wire [13:0] _GEN_4327 = 14'h10e7 == index ? 14'h21 : _GEN_4326;
  wire [13:0] _GEN_4328 = 14'h10e8 == index ? 14'h21 : _GEN_4327;
  wire [13:0] _GEN_4329 = 14'h10e9 == index ? 14'h21 : _GEN_4328;
  wire [13:0] _GEN_4330 = 14'h10ea == index ? 14'h21 : _GEN_4329;
  wire [13:0] _GEN_4331 = 14'h10eb == index ? 14'h21 : _GEN_4330;
  wire [13:0] _GEN_4332 = 14'h10ec == index ? 14'h21 : _GEN_4331;
  wire [13:0] _GEN_4333 = 14'h10ed == index ? 14'h21 : _GEN_4332;
  wire [13:0] _GEN_4334 = 14'h10ee == index ? 14'h21 : _GEN_4333;
  wire [13:0] _GEN_4335 = 14'h10ef == index ? 14'h21 : _GEN_4334;
  wire [13:0] _GEN_4336 = 14'h10f0 == index ? 14'h21 : _GEN_4335;
  wire [13:0] _GEN_4337 = 14'h10f1 == index ? 14'h21 : _GEN_4336;
  wire [13:0] _GEN_4338 = 14'h10f2 == index ? 14'h21 : _GEN_4337;
  wire [13:0] _GEN_4339 = 14'h10f3 == index ? 14'h21 : _GEN_4338;
  wire [13:0] _GEN_4340 = 14'h10f4 == index ? 14'h21 : _GEN_4339;
  wire [13:0] _GEN_4341 = 14'h10f5 == index ? 14'h21 : _GEN_4340;
  wire [13:0] _GEN_4342 = 14'h10f6 == index ? 14'h21 : _GEN_4341;
  wire [13:0] _GEN_4343 = 14'h10f7 == index ? 14'h21 : _GEN_4342;
  wire [13:0] _GEN_4344 = 14'h10f8 == index ? 14'h21 : _GEN_4343;
  wire [13:0] _GEN_4345 = 14'h10f9 == index ? 14'h21 : _GEN_4344;
  wire [13:0] _GEN_4346 = 14'h10fa == index ? 14'h21 : _GEN_4345;
  wire [13:0] _GEN_4347 = 14'h10fb == index ? 14'h21 : _GEN_4346;
  wire [13:0] _GEN_4348 = 14'h10fc == index ? 14'h21 : _GEN_4347;
  wire [13:0] _GEN_4349 = 14'h10fd == index ? 14'h21 : _GEN_4348;
  wire [13:0] _GEN_4350 = 14'h10fe == index ? 14'h21 : _GEN_4349;
  wire [13:0] _GEN_4351 = 14'h10ff == index ? 14'h21 : _GEN_4350;
  wire [13:0] _GEN_4352 = 14'h1100 == index ? 14'h0 : _GEN_4351;
  wire [13:0] _GEN_4353 = 14'h1101 == index ? 14'h1100 : _GEN_4352;
  wire [13:0] _GEN_4354 = 14'h1102 == index ? 14'h880 : _GEN_4353;
  wire [13:0] _GEN_4355 = 14'h1103 == index ? 14'h581 : _GEN_4354;
  wire [13:0] _GEN_4356 = 14'h1104 == index ? 14'h402 : _GEN_4355;
  wire [13:0] _GEN_4357 = 14'h1105 == index ? 14'h304 : _GEN_4356;
  wire [13:0] _GEN_4358 = 14'h1106 == index ? 14'h284 : _GEN_4357;
  wire [13:0] _GEN_4359 = 14'h1107 == index ? 14'h206 : _GEN_4358;
  wire [13:0] _GEN_4360 = 14'h1108 == index ? 14'h202 : _GEN_4359;
  wire [13:0] _GEN_4361 = 14'h1109 == index ? 14'h187 : _GEN_4360;
  wire [13:0] _GEN_4362 = 14'h110a == index ? 14'h184 : _GEN_4361;
  wire [13:0] _GEN_4363 = 14'h110b == index ? 14'h181 : _GEN_4362;
  wire [13:0] _GEN_4364 = 14'h110c == index ? 14'h10a : _GEN_4363;
  wire [13:0] _GEN_4365 = 14'h110d == index ? 14'h108 : _GEN_4364;
  wire [13:0] _GEN_4366 = 14'h110e == index ? 14'h106 : _GEN_4365;
  wire [13:0] _GEN_4367 = 14'h110f == index ? 14'h104 : _GEN_4366;
  wire [13:0] _GEN_4368 = 14'h1110 == index ? 14'h102 : _GEN_4367;
  wire [13:0] _GEN_4369 = 14'h1111 == index ? 14'h100 : _GEN_4368;
  wire [13:0] _GEN_4370 = 14'h1112 == index ? 14'h90 : _GEN_4369;
  wire [13:0] _GEN_4371 = 14'h1113 == index ? 14'h8f : _GEN_4370;
  wire [13:0] _GEN_4372 = 14'h1114 == index ? 14'h8e : _GEN_4371;
  wire [13:0] _GEN_4373 = 14'h1115 == index ? 14'h8d : _GEN_4372;
  wire [13:0] _GEN_4374 = 14'h1116 == index ? 14'h8c : _GEN_4373;
  wire [13:0] _GEN_4375 = 14'h1117 == index ? 14'h8b : _GEN_4374;
  wire [13:0] _GEN_4376 = 14'h1118 == index ? 14'h8a : _GEN_4375;
  wire [13:0] _GEN_4377 = 14'h1119 == index ? 14'h89 : _GEN_4376;
  wire [13:0] _GEN_4378 = 14'h111a == index ? 14'h88 : _GEN_4377;
  wire [13:0] _GEN_4379 = 14'h111b == index ? 14'h87 : _GEN_4378;
  wire [13:0] _GEN_4380 = 14'h111c == index ? 14'h86 : _GEN_4379;
  wire [13:0] _GEN_4381 = 14'h111d == index ? 14'h85 : _GEN_4380;
  wire [13:0] _GEN_4382 = 14'h111e == index ? 14'h84 : _GEN_4381;
  wire [13:0] _GEN_4383 = 14'h111f == index ? 14'h83 : _GEN_4382;
  wire [13:0] _GEN_4384 = 14'h1120 == index ? 14'h82 : _GEN_4383;
  wire [13:0] _GEN_4385 = 14'h1121 == index ? 14'h81 : _GEN_4384;
  wire [13:0] _GEN_4386 = 14'h1122 == index ? 14'h80 : _GEN_4385;
  wire [13:0] _GEN_4387 = 14'h1123 == index ? 14'h22 : _GEN_4386;
  wire [13:0] _GEN_4388 = 14'h1124 == index ? 14'h22 : _GEN_4387;
  wire [13:0] _GEN_4389 = 14'h1125 == index ? 14'h22 : _GEN_4388;
  wire [13:0] _GEN_4390 = 14'h1126 == index ? 14'h22 : _GEN_4389;
  wire [13:0] _GEN_4391 = 14'h1127 == index ? 14'h22 : _GEN_4390;
  wire [13:0] _GEN_4392 = 14'h1128 == index ? 14'h22 : _GEN_4391;
  wire [13:0] _GEN_4393 = 14'h1129 == index ? 14'h22 : _GEN_4392;
  wire [13:0] _GEN_4394 = 14'h112a == index ? 14'h22 : _GEN_4393;
  wire [13:0] _GEN_4395 = 14'h112b == index ? 14'h22 : _GEN_4394;
  wire [13:0] _GEN_4396 = 14'h112c == index ? 14'h22 : _GEN_4395;
  wire [13:0] _GEN_4397 = 14'h112d == index ? 14'h22 : _GEN_4396;
  wire [13:0] _GEN_4398 = 14'h112e == index ? 14'h22 : _GEN_4397;
  wire [13:0] _GEN_4399 = 14'h112f == index ? 14'h22 : _GEN_4398;
  wire [13:0] _GEN_4400 = 14'h1130 == index ? 14'h22 : _GEN_4399;
  wire [13:0] _GEN_4401 = 14'h1131 == index ? 14'h22 : _GEN_4400;
  wire [13:0] _GEN_4402 = 14'h1132 == index ? 14'h22 : _GEN_4401;
  wire [13:0] _GEN_4403 = 14'h1133 == index ? 14'h22 : _GEN_4402;
  wire [13:0] _GEN_4404 = 14'h1134 == index ? 14'h22 : _GEN_4403;
  wire [13:0] _GEN_4405 = 14'h1135 == index ? 14'h22 : _GEN_4404;
  wire [13:0] _GEN_4406 = 14'h1136 == index ? 14'h22 : _GEN_4405;
  wire [13:0] _GEN_4407 = 14'h1137 == index ? 14'h22 : _GEN_4406;
  wire [13:0] _GEN_4408 = 14'h1138 == index ? 14'h22 : _GEN_4407;
  wire [13:0] _GEN_4409 = 14'h1139 == index ? 14'h22 : _GEN_4408;
  wire [13:0] _GEN_4410 = 14'h113a == index ? 14'h22 : _GEN_4409;
  wire [13:0] _GEN_4411 = 14'h113b == index ? 14'h22 : _GEN_4410;
  wire [13:0] _GEN_4412 = 14'h113c == index ? 14'h22 : _GEN_4411;
  wire [13:0] _GEN_4413 = 14'h113d == index ? 14'h22 : _GEN_4412;
  wire [13:0] _GEN_4414 = 14'h113e == index ? 14'h22 : _GEN_4413;
  wire [13:0] _GEN_4415 = 14'h113f == index ? 14'h22 : _GEN_4414;
  wire [13:0] _GEN_4416 = 14'h1140 == index ? 14'h22 : _GEN_4415;
  wire [13:0] _GEN_4417 = 14'h1141 == index ? 14'h22 : _GEN_4416;
  wire [13:0] _GEN_4418 = 14'h1142 == index ? 14'h22 : _GEN_4417;
  wire [13:0] _GEN_4419 = 14'h1143 == index ? 14'h22 : _GEN_4418;
  wire [13:0] _GEN_4420 = 14'h1144 == index ? 14'h22 : _GEN_4419;
  wire [13:0] _GEN_4421 = 14'h1145 == index ? 14'h22 : _GEN_4420;
  wire [13:0] _GEN_4422 = 14'h1146 == index ? 14'h22 : _GEN_4421;
  wire [13:0] _GEN_4423 = 14'h1147 == index ? 14'h22 : _GEN_4422;
  wire [13:0] _GEN_4424 = 14'h1148 == index ? 14'h22 : _GEN_4423;
  wire [13:0] _GEN_4425 = 14'h1149 == index ? 14'h22 : _GEN_4424;
  wire [13:0] _GEN_4426 = 14'h114a == index ? 14'h22 : _GEN_4425;
  wire [13:0] _GEN_4427 = 14'h114b == index ? 14'h22 : _GEN_4426;
  wire [13:0] _GEN_4428 = 14'h114c == index ? 14'h22 : _GEN_4427;
  wire [13:0] _GEN_4429 = 14'h114d == index ? 14'h22 : _GEN_4428;
  wire [13:0] _GEN_4430 = 14'h114e == index ? 14'h22 : _GEN_4429;
  wire [13:0] _GEN_4431 = 14'h114f == index ? 14'h22 : _GEN_4430;
  wire [13:0] _GEN_4432 = 14'h1150 == index ? 14'h22 : _GEN_4431;
  wire [13:0] _GEN_4433 = 14'h1151 == index ? 14'h22 : _GEN_4432;
  wire [13:0] _GEN_4434 = 14'h1152 == index ? 14'h22 : _GEN_4433;
  wire [13:0] _GEN_4435 = 14'h1153 == index ? 14'h22 : _GEN_4434;
  wire [13:0] _GEN_4436 = 14'h1154 == index ? 14'h22 : _GEN_4435;
  wire [13:0] _GEN_4437 = 14'h1155 == index ? 14'h22 : _GEN_4436;
  wire [13:0] _GEN_4438 = 14'h1156 == index ? 14'h22 : _GEN_4437;
  wire [13:0] _GEN_4439 = 14'h1157 == index ? 14'h22 : _GEN_4438;
  wire [13:0] _GEN_4440 = 14'h1158 == index ? 14'h22 : _GEN_4439;
  wire [13:0] _GEN_4441 = 14'h1159 == index ? 14'h22 : _GEN_4440;
  wire [13:0] _GEN_4442 = 14'h115a == index ? 14'h22 : _GEN_4441;
  wire [13:0] _GEN_4443 = 14'h115b == index ? 14'h22 : _GEN_4442;
  wire [13:0] _GEN_4444 = 14'h115c == index ? 14'h22 : _GEN_4443;
  wire [13:0] _GEN_4445 = 14'h115d == index ? 14'h22 : _GEN_4444;
  wire [13:0] _GEN_4446 = 14'h115e == index ? 14'h22 : _GEN_4445;
  wire [13:0] _GEN_4447 = 14'h115f == index ? 14'h22 : _GEN_4446;
  wire [13:0] _GEN_4448 = 14'h1160 == index ? 14'h22 : _GEN_4447;
  wire [13:0] _GEN_4449 = 14'h1161 == index ? 14'h22 : _GEN_4448;
  wire [13:0] _GEN_4450 = 14'h1162 == index ? 14'h22 : _GEN_4449;
  wire [13:0] _GEN_4451 = 14'h1163 == index ? 14'h22 : _GEN_4450;
  wire [13:0] _GEN_4452 = 14'h1164 == index ? 14'h22 : _GEN_4451;
  wire [13:0] _GEN_4453 = 14'h1165 == index ? 14'h22 : _GEN_4452;
  wire [13:0] _GEN_4454 = 14'h1166 == index ? 14'h22 : _GEN_4453;
  wire [13:0] _GEN_4455 = 14'h1167 == index ? 14'h22 : _GEN_4454;
  wire [13:0] _GEN_4456 = 14'h1168 == index ? 14'h22 : _GEN_4455;
  wire [13:0] _GEN_4457 = 14'h1169 == index ? 14'h22 : _GEN_4456;
  wire [13:0] _GEN_4458 = 14'h116a == index ? 14'h22 : _GEN_4457;
  wire [13:0] _GEN_4459 = 14'h116b == index ? 14'h22 : _GEN_4458;
  wire [13:0] _GEN_4460 = 14'h116c == index ? 14'h22 : _GEN_4459;
  wire [13:0] _GEN_4461 = 14'h116d == index ? 14'h22 : _GEN_4460;
  wire [13:0] _GEN_4462 = 14'h116e == index ? 14'h22 : _GEN_4461;
  wire [13:0] _GEN_4463 = 14'h116f == index ? 14'h22 : _GEN_4462;
  wire [13:0] _GEN_4464 = 14'h1170 == index ? 14'h22 : _GEN_4463;
  wire [13:0] _GEN_4465 = 14'h1171 == index ? 14'h22 : _GEN_4464;
  wire [13:0] _GEN_4466 = 14'h1172 == index ? 14'h22 : _GEN_4465;
  wire [13:0] _GEN_4467 = 14'h1173 == index ? 14'h22 : _GEN_4466;
  wire [13:0] _GEN_4468 = 14'h1174 == index ? 14'h22 : _GEN_4467;
  wire [13:0] _GEN_4469 = 14'h1175 == index ? 14'h22 : _GEN_4468;
  wire [13:0] _GEN_4470 = 14'h1176 == index ? 14'h22 : _GEN_4469;
  wire [13:0] _GEN_4471 = 14'h1177 == index ? 14'h22 : _GEN_4470;
  wire [13:0] _GEN_4472 = 14'h1178 == index ? 14'h22 : _GEN_4471;
  wire [13:0] _GEN_4473 = 14'h1179 == index ? 14'h22 : _GEN_4472;
  wire [13:0] _GEN_4474 = 14'h117a == index ? 14'h22 : _GEN_4473;
  wire [13:0] _GEN_4475 = 14'h117b == index ? 14'h22 : _GEN_4474;
  wire [13:0] _GEN_4476 = 14'h117c == index ? 14'h22 : _GEN_4475;
  wire [13:0] _GEN_4477 = 14'h117d == index ? 14'h22 : _GEN_4476;
  wire [13:0] _GEN_4478 = 14'h117e == index ? 14'h22 : _GEN_4477;
  wire [13:0] _GEN_4479 = 14'h117f == index ? 14'h22 : _GEN_4478;
  wire [13:0] _GEN_4480 = 14'h1180 == index ? 14'h0 : _GEN_4479;
  wire [13:0] _GEN_4481 = 14'h1181 == index ? 14'h1180 : _GEN_4480;
  wire [13:0] _GEN_4482 = 14'h1182 == index ? 14'h881 : _GEN_4481;
  wire [13:0] _GEN_4483 = 14'h1183 == index ? 14'h582 : _GEN_4482;
  wire [13:0] _GEN_4484 = 14'h1184 == index ? 14'h403 : _GEN_4483;
  wire [13:0] _GEN_4485 = 14'h1185 == index ? 14'h380 : _GEN_4484;
  wire [13:0] _GEN_4486 = 14'h1186 == index ? 14'h285 : _GEN_4485;
  wire [13:0] _GEN_4487 = 14'h1187 == index ? 14'h280 : _GEN_4486;
  wire [13:0] _GEN_4488 = 14'h1188 == index ? 14'h203 : _GEN_4487;
  wire [13:0] _GEN_4489 = 14'h1189 == index ? 14'h188 : _GEN_4488;
  wire [13:0] _GEN_4490 = 14'h118a == index ? 14'h185 : _GEN_4489;
  wire [13:0] _GEN_4491 = 14'h118b == index ? 14'h182 : _GEN_4490;
  wire [13:0] _GEN_4492 = 14'h118c == index ? 14'h10b : _GEN_4491;
  wire [13:0] _GEN_4493 = 14'h118d == index ? 14'h109 : _GEN_4492;
  wire [13:0] _GEN_4494 = 14'h118e == index ? 14'h107 : _GEN_4493;
  wire [13:0] _GEN_4495 = 14'h118f == index ? 14'h105 : _GEN_4494;
  wire [13:0] _GEN_4496 = 14'h1190 == index ? 14'h103 : _GEN_4495;
  wire [13:0] _GEN_4497 = 14'h1191 == index ? 14'h101 : _GEN_4496;
  wire [13:0] _GEN_4498 = 14'h1192 == index ? 14'h91 : _GEN_4497;
  wire [13:0] _GEN_4499 = 14'h1193 == index ? 14'h90 : _GEN_4498;
  wire [13:0] _GEN_4500 = 14'h1194 == index ? 14'h8f : _GEN_4499;
  wire [13:0] _GEN_4501 = 14'h1195 == index ? 14'h8e : _GEN_4500;
  wire [13:0] _GEN_4502 = 14'h1196 == index ? 14'h8d : _GEN_4501;
  wire [13:0] _GEN_4503 = 14'h1197 == index ? 14'h8c : _GEN_4502;
  wire [13:0] _GEN_4504 = 14'h1198 == index ? 14'h8b : _GEN_4503;
  wire [13:0] _GEN_4505 = 14'h1199 == index ? 14'h8a : _GEN_4504;
  wire [13:0] _GEN_4506 = 14'h119a == index ? 14'h89 : _GEN_4505;
  wire [13:0] _GEN_4507 = 14'h119b == index ? 14'h88 : _GEN_4506;
  wire [13:0] _GEN_4508 = 14'h119c == index ? 14'h87 : _GEN_4507;
  wire [13:0] _GEN_4509 = 14'h119d == index ? 14'h86 : _GEN_4508;
  wire [13:0] _GEN_4510 = 14'h119e == index ? 14'h85 : _GEN_4509;
  wire [13:0] _GEN_4511 = 14'h119f == index ? 14'h84 : _GEN_4510;
  wire [13:0] _GEN_4512 = 14'h11a0 == index ? 14'h83 : _GEN_4511;
  wire [13:0] _GEN_4513 = 14'h11a1 == index ? 14'h82 : _GEN_4512;
  wire [13:0] _GEN_4514 = 14'h11a2 == index ? 14'h81 : _GEN_4513;
  wire [13:0] _GEN_4515 = 14'h11a3 == index ? 14'h80 : _GEN_4514;
  wire [13:0] _GEN_4516 = 14'h11a4 == index ? 14'h23 : _GEN_4515;
  wire [13:0] _GEN_4517 = 14'h11a5 == index ? 14'h23 : _GEN_4516;
  wire [13:0] _GEN_4518 = 14'h11a6 == index ? 14'h23 : _GEN_4517;
  wire [13:0] _GEN_4519 = 14'h11a7 == index ? 14'h23 : _GEN_4518;
  wire [13:0] _GEN_4520 = 14'h11a8 == index ? 14'h23 : _GEN_4519;
  wire [13:0] _GEN_4521 = 14'h11a9 == index ? 14'h23 : _GEN_4520;
  wire [13:0] _GEN_4522 = 14'h11aa == index ? 14'h23 : _GEN_4521;
  wire [13:0] _GEN_4523 = 14'h11ab == index ? 14'h23 : _GEN_4522;
  wire [13:0] _GEN_4524 = 14'h11ac == index ? 14'h23 : _GEN_4523;
  wire [13:0] _GEN_4525 = 14'h11ad == index ? 14'h23 : _GEN_4524;
  wire [13:0] _GEN_4526 = 14'h11ae == index ? 14'h23 : _GEN_4525;
  wire [13:0] _GEN_4527 = 14'h11af == index ? 14'h23 : _GEN_4526;
  wire [13:0] _GEN_4528 = 14'h11b0 == index ? 14'h23 : _GEN_4527;
  wire [13:0] _GEN_4529 = 14'h11b1 == index ? 14'h23 : _GEN_4528;
  wire [13:0] _GEN_4530 = 14'h11b2 == index ? 14'h23 : _GEN_4529;
  wire [13:0] _GEN_4531 = 14'h11b3 == index ? 14'h23 : _GEN_4530;
  wire [13:0] _GEN_4532 = 14'h11b4 == index ? 14'h23 : _GEN_4531;
  wire [13:0] _GEN_4533 = 14'h11b5 == index ? 14'h23 : _GEN_4532;
  wire [13:0] _GEN_4534 = 14'h11b6 == index ? 14'h23 : _GEN_4533;
  wire [13:0] _GEN_4535 = 14'h11b7 == index ? 14'h23 : _GEN_4534;
  wire [13:0] _GEN_4536 = 14'h11b8 == index ? 14'h23 : _GEN_4535;
  wire [13:0] _GEN_4537 = 14'h11b9 == index ? 14'h23 : _GEN_4536;
  wire [13:0] _GEN_4538 = 14'h11ba == index ? 14'h23 : _GEN_4537;
  wire [13:0] _GEN_4539 = 14'h11bb == index ? 14'h23 : _GEN_4538;
  wire [13:0] _GEN_4540 = 14'h11bc == index ? 14'h23 : _GEN_4539;
  wire [13:0] _GEN_4541 = 14'h11bd == index ? 14'h23 : _GEN_4540;
  wire [13:0] _GEN_4542 = 14'h11be == index ? 14'h23 : _GEN_4541;
  wire [13:0] _GEN_4543 = 14'h11bf == index ? 14'h23 : _GEN_4542;
  wire [13:0] _GEN_4544 = 14'h11c0 == index ? 14'h23 : _GEN_4543;
  wire [13:0] _GEN_4545 = 14'h11c1 == index ? 14'h23 : _GEN_4544;
  wire [13:0] _GEN_4546 = 14'h11c2 == index ? 14'h23 : _GEN_4545;
  wire [13:0] _GEN_4547 = 14'h11c3 == index ? 14'h23 : _GEN_4546;
  wire [13:0] _GEN_4548 = 14'h11c4 == index ? 14'h23 : _GEN_4547;
  wire [13:0] _GEN_4549 = 14'h11c5 == index ? 14'h23 : _GEN_4548;
  wire [13:0] _GEN_4550 = 14'h11c6 == index ? 14'h23 : _GEN_4549;
  wire [13:0] _GEN_4551 = 14'h11c7 == index ? 14'h23 : _GEN_4550;
  wire [13:0] _GEN_4552 = 14'h11c8 == index ? 14'h23 : _GEN_4551;
  wire [13:0] _GEN_4553 = 14'h11c9 == index ? 14'h23 : _GEN_4552;
  wire [13:0] _GEN_4554 = 14'h11ca == index ? 14'h23 : _GEN_4553;
  wire [13:0] _GEN_4555 = 14'h11cb == index ? 14'h23 : _GEN_4554;
  wire [13:0] _GEN_4556 = 14'h11cc == index ? 14'h23 : _GEN_4555;
  wire [13:0] _GEN_4557 = 14'h11cd == index ? 14'h23 : _GEN_4556;
  wire [13:0] _GEN_4558 = 14'h11ce == index ? 14'h23 : _GEN_4557;
  wire [13:0] _GEN_4559 = 14'h11cf == index ? 14'h23 : _GEN_4558;
  wire [13:0] _GEN_4560 = 14'h11d0 == index ? 14'h23 : _GEN_4559;
  wire [13:0] _GEN_4561 = 14'h11d1 == index ? 14'h23 : _GEN_4560;
  wire [13:0] _GEN_4562 = 14'h11d2 == index ? 14'h23 : _GEN_4561;
  wire [13:0] _GEN_4563 = 14'h11d3 == index ? 14'h23 : _GEN_4562;
  wire [13:0] _GEN_4564 = 14'h11d4 == index ? 14'h23 : _GEN_4563;
  wire [13:0] _GEN_4565 = 14'h11d5 == index ? 14'h23 : _GEN_4564;
  wire [13:0] _GEN_4566 = 14'h11d6 == index ? 14'h23 : _GEN_4565;
  wire [13:0] _GEN_4567 = 14'h11d7 == index ? 14'h23 : _GEN_4566;
  wire [13:0] _GEN_4568 = 14'h11d8 == index ? 14'h23 : _GEN_4567;
  wire [13:0] _GEN_4569 = 14'h11d9 == index ? 14'h23 : _GEN_4568;
  wire [13:0] _GEN_4570 = 14'h11da == index ? 14'h23 : _GEN_4569;
  wire [13:0] _GEN_4571 = 14'h11db == index ? 14'h23 : _GEN_4570;
  wire [13:0] _GEN_4572 = 14'h11dc == index ? 14'h23 : _GEN_4571;
  wire [13:0] _GEN_4573 = 14'h11dd == index ? 14'h23 : _GEN_4572;
  wire [13:0] _GEN_4574 = 14'h11de == index ? 14'h23 : _GEN_4573;
  wire [13:0] _GEN_4575 = 14'h11df == index ? 14'h23 : _GEN_4574;
  wire [13:0] _GEN_4576 = 14'h11e0 == index ? 14'h23 : _GEN_4575;
  wire [13:0] _GEN_4577 = 14'h11e1 == index ? 14'h23 : _GEN_4576;
  wire [13:0] _GEN_4578 = 14'h11e2 == index ? 14'h23 : _GEN_4577;
  wire [13:0] _GEN_4579 = 14'h11e3 == index ? 14'h23 : _GEN_4578;
  wire [13:0] _GEN_4580 = 14'h11e4 == index ? 14'h23 : _GEN_4579;
  wire [13:0] _GEN_4581 = 14'h11e5 == index ? 14'h23 : _GEN_4580;
  wire [13:0] _GEN_4582 = 14'h11e6 == index ? 14'h23 : _GEN_4581;
  wire [13:0] _GEN_4583 = 14'h11e7 == index ? 14'h23 : _GEN_4582;
  wire [13:0] _GEN_4584 = 14'h11e8 == index ? 14'h23 : _GEN_4583;
  wire [13:0] _GEN_4585 = 14'h11e9 == index ? 14'h23 : _GEN_4584;
  wire [13:0] _GEN_4586 = 14'h11ea == index ? 14'h23 : _GEN_4585;
  wire [13:0] _GEN_4587 = 14'h11eb == index ? 14'h23 : _GEN_4586;
  wire [13:0] _GEN_4588 = 14'h11ec == index ? 14'h23 : _GEN_4587;
  wire [13:0] _GEN_4589 = 14'h11ed == index ? 14'h23 : _GEN_4588;
  wire [13:0] _GEN_4590 = 14'h11ee == index ? 14'h23 : _GEN_4589;
  wire [13:0] _GEN_4591 = 14'h11ef == index ? 14'h23 : _GEN_4590;
  wire [13:0] _GEN_4592 = 14'h11f0 == index ? 14'h23 : _GEN_4591;
  wire [13:0] _GEN_4593 = 14'h11f1 == index ? 14'h23 : _GEN_4592;
  wire [13:0] _GEN_4594 = 14'h11f2 == index ? 14'h23 : _GEN_4593;
  wire [13:0] _GEN_4595 = 14'h11f3 == index ? 14'h23 : _GEN_4594;
  wire [13:0] _GEN_4596 = 14'h11f4 == index ? 14'h23 : _GEN_4595;
  wire [13:0] _GEN_4597 = 14'h11f5 == index ? 14'h23 : _GEN_4596;
  wire [13:0] _GEN_4598 = 14'h11f6 == index ? 14'h23 : _GEN_4597;
  wire [13:0] _GEN_4599 = 14'h11f7 == index ? 14'h23 : _GEN_4598;
  wire [13:0] _GEN_4600 = 14'h11f8 == index ? 14'h23 : _GEN_4599;
  wire [13:0] _GEN_4601 = 14'h11f9 == index ? 14'h23 : _GEN_4600;
  wire [13:0] _GEN_4602 = 14'h11fa == index ? 14'h23 : _GEN_4601;
  wire [13:0] _GEN_4603 = 14'h11fb == index ? 14'h23 : _GEN_4602;
  wire [13:0] _GEN_4604 = 14'h11fc == index ? 14'h23 : _GEN_4603;
  wire [13:0] _GEN_4605 = 14'h11fd == index ? 14'h23 : _GEN_4604;
  wire [13:0] _GEN_4606 = 14'h11fe == index ? 14'h23 : _GEN_4605;
  wire [13:0] _GEN_4607 = 14'h11ff == index ? 14'h23 : _GEN_4606;
  wire [13:0] _GEN_4608 = 14'h1200 == index ? 14'h0 : _GEN_4607;
  wire [13:0] _GEN_4609 = 14'h1201 == index ? 14'h1200 : _GEN_4608;
  wire [13:0] _GEN_4610 = 14'h1202 == index ? 14'h900 : _GEN_4609;
  wire [13:0] _GEN_4611 = 14'h1203 == index ? 14'h600 : _GEN_4610;
  wire [13:0] _GEN_4612 = 14'h1204 == index ? 14'h480 : _GEN_4611;
  wire [13:0] _GEN_4613 = 14'h1205 == index ? 14'h381 : _GEN_4612;
  wire [13:0] _GEN_4614 = 14'h1206 == index ? 14'h300 : _GEN_4613;
  wire [13:0] _GEN_4615 = 14'h1207 == index ? 14'h281 : _GEN_4614;
  wire [13:0] _GEN_4616 = 14'h1208 == index ? 14'h204 : _GEN_4615;
  wire [13:0] _GEN_4617 = 14'h1209 == index ? 14'h200 : _GEN_4616;
  wire [13:0] _GEN_4618 = 14'h120a == index ? 14'h186 : _GEN_4617;
  wire [13:0] _GEN_4619 = 14'h120b == index ? 14'h183 : _GEN_4618;
  wire [13:0] _GEN_4620 = 14'h120c == index ? 14'h180 : _GEN_4619;
  wire [13:0] _GEN_4621 = 14'h120d == index ? 14'h10a : _GEN_4620;
  wire [13:0] _GEN_4622 = 14'h120e == index ? 14'h108 : _GEN_4621;
  wire [13:0] _GEN_4623 = 14'h120f == index ? 14'h106 : _GEN_4622;
  wire [13:0] _GEN_4624 = 14'h1210 == index ? 14'h104 : _GEN_4623;
  wire [13:0] _GEN_4625 = 14'h1211 == index ? 14'h102 : _GEN_4624;
  wire [13:0] _GEN_4626 = 14'h1212 == index ? 14'h100 : _GEN_4625;
  wire [13:0] _GEN_4627 = 14'h1213 == index ? 14'h91 : _GEN_4626;
  wire [13:0] _GEN_4628 = 14'h1214 == index ? 14'h90 : _GEN_4627;
  wire [13:0] _GEN_4629 = 14'h1215 == index ? 14'h8f : _GEN_4628;
  wire [13:0] _GEN_4630 = 14'h1216 == index ? 14'h8e : _GEN_4629;
  wire [13:0] _GEN_4631 = 14'h1217 == index ? 14'h8d : _GEN_4630;
  wire [13:0] _GEN_4632 = 14'h1218 == index ? 14'h8c : _GEN_4631;
  wire [13:0] _GEN_4633 = 14'h1219 == index ? 14'h8b : _GEN_4632;
  wire [13:0] _GEN_4634 = 14'h121a == index ? 14'h8a : _GEN_4633;
  wire [13:0] _GEN_4635 = 14'h121b == index ? 14'h89 : _GEN_4634;
  wire [13:0] _GEN_4636 = 14'h121c == index ? 14'h88 : _GEN_4635;
  wire [13:0] _GEN_4637 = 14'h121d == index ? 14'h87 : _GEN_4636;
  wire [13:0] _GEN_4638 = 14'h121e == index ? 14'h86 : _GEN_4637;
  wire [13:0] _GEN_4639 = 14'h121f == index ? 14'h85 : _GEN_4638;
  wire [13:0] _GEN_4640 = 14'h1220 == index ? 14'h84 : _GEN_4639;
  wire [13:0] _GEN_4641 = 14'h1221 == index ? 14'h83 : _GEN_4640;
  wire [13:0] _GEN_4642 = 14'h1222 == index ? 14'h82 : _GEN_4641;
  wire [13:0] _GEN_4643 = 14'h1223 == index ? 14'h81 : _GEN_4642;
  wire [13:0] _GEN_4644 = 14'h1224 == index ? 14'h80 : _GEN_4643;
  wire [13:0] _GEN_4645 = 14'h1225 == index ? 14'h24 : _GEN_4644;
  wire [13:0] _GEN_4646 = 14'h1226 == index ? 14'h24 : _GEN_4645;
  wire [13:0] _GEN_4647 = 14'h1227 == index ? 14'h24 : _GEN_4646;
  wire [13:0] _GEN_4648 = 14'h1228 == index ? 14'h24 : _GEN_4647;
  wire [13:0] _GEN_4649 = 14'h1229 == index ? 14'h24 : _GEN_4648;
  wire [13:0] _GEN_4650 = 14'h122a == index ? 14'h24 : _GEN_4649;
  wire [13:0] _GEN_4651 = 14'h122b == index ? 14'h24 : _GEN_4650;
  wire [13:0] _GEN_4652 = 14'h122c == index ? 14'h24 : _GEN_4651;
  wire [13:0] _GEN_4653 = 14'h122d == index ? 14'h24 : _GEN_4652;
  wire [13:0] _GEN_4654 = 14'h122e == index ? 14'h24 : _GEN_4653;
  wire [13:0] _GEN_4655 = 14'h122f == index ? 14'h24 : _GEN_4654;
  wire [13:0] _GEN_4656 = 14'h1230 == index ? 14'h24 : _GEN_4655;
  wire [13:0] _GEN_4657 = 14'h1231 == index ? 14'h24 : _GEN_4656;
  wire [13:0] _GEN_4658 = 14'h1232 == index ? 14'h24 : _GEN_4657;
  wire [13:0] _GEN_4659 = 14'h1233 == index ? 14'h24 : _GEN_4658;
  wire [13:0] _GEN_4660 = 14'h1234 == index ? 14'h24 : _GEN_4659;
  wire [13:0] _GEN_4661 = 14'h1235 == index ? 14'h24 : _GEN_4660;
  wire [13:0] _GEN_4662 = 14'h1236 == index ? 14'h24 : _GEN_4661;
  wire [13:0] _GEN_4663 = 14'h1237 == index ? 14'h24 : _GEN_4662;
  wire [13:0] _GEN_4664 = 14'h1238 == index ? 14'h24 : _GEN_4663;
  wire [13:0] _GEN_4665 = 14'h1239 == index ? 14'h24 : _GEN_4664;
  wire [13:0] _GEN_4666 = 14'h123a == index ? 14'h24 : _GEN_4665;
  wire [13:0] _GEN_4667 = 14'h123b == index ? 14'h24 : _GEN_4666;
  wire [13:0] _GEN_4668 = 14'h123c == index ? 14'h24 : _GEN_4667;
  wire [13:0] _GEN_4669 = 14'h123d == index ? 14'h24 : _GEN_4668;
  wire [13:0] _GEN_4670 = 14'h123e == index ? 14'h24 : _GEN_4669;
  wire [13:0] _GEN_4671 = 14'h123f == index ? 14'h24 : _GEN_4670;
  wire [13:0] _GEN_4672 = 14'h1240 == index ? 14'h24 : _GEN_4671;
  wire [13:0] _GEN_4673 = 14'h1241 == index ? 14'h24 : _GEN_4672;
  wire [13:0] _GEN_4674 = 14'h1242 == index ? 14'h24 : _GEN_4673;
  wire [13:0] _GEN_4675 = 14'h1243 == index ? 14'h24 : _GEN_4674;
  wire [13:0] _GEN_4676 = 14'h1244 == index ? 14'h24 : _GEN_4675;
  wire [13:0] _GEN_4677 = 14'h1245 == index ? 14'h24 : _GEN_4676;
  wire [13:0] _GEN_4678 = 14'h1246 == index ? 14'h24 : _GEN_4677;
  wire [13:0] _GEN_4679 = 14'h1247 == index ? 14'h24 : _GEN_4678;
  wire [13:0] _GEN_4680 = 14'h1248 == index ? 14'h24 : _GEN_4679;
  wire [13:0] _GEN_4681 = 14'h1249 == index ? 14'h24 : _GEN_4680;
  wire [13:0] _GEN_4682 = 14'h124a == index ? 14'h24 : _GEN_4681;
  wire [13:0] _GEN_4683 = 14'h124b == index ? 14'h24 : _GEN_4682;
  wire [13:0] _GEN_4684 = 14'h124c == index ? 14'h24 : _GEN_4683;
  wire [13:0] _GEN_4685 = 14'h124d == index ? 14'h24 : _GEN_4684;
  wire [13:0] _GEN_4686 = 14'h124e == index ? 14'h24 : _GEN_4685;
  wire [13:0] _GEN_4687 = 14'h124f == index ? 14'h24 : _GEN_4686;
  wire [13:0] _GEN_4688 = 14'h1250 == index ? 14'h24 : _GEN_4687;
  wire [13:0] _GEN_4689 = 14'h1251 == index ? 14'h24 : _GEN_4688;
  wire [13:0] _GEN_4690 = 14'h1252 == index ? 14'h24 : _GEN_4689;
  wire [13:0] _GEN_4691 = 14'h1253 == index ? 14'h24 : _GEN_4690;
  wire [13:0] _GEN_4692 = 14'h1254 == index ? 14'h24 : _GEN_4691;
  wire [13:0] _GEN_4693 = 14'h1255 == index ? 14'h24 : _GEN_4692;
  wire [13:0] _GEN_4694 = 14'h1256 == index ? 14'h24 : _GEN_4693;
  wire [13:0] _GEN_4695 = 14'h1257 == index ? 14'h24 : _GEN_4694;
  wire [13:0] _GEN_4696 = 14'h1258 == index ? 14'h24 : _GEN_4695;
  wire [13:0] _GEN_4697 = 14'h1259 == index ? 14'h24 : _GEN_4696;
  wire [13:0] _GEN_4698 = 14'h125a == index ? 14'h24 : _GEN_4697;
  wire [13:0] _GEN_4699 = 14'h125b == index ? 14'h24 : _GEN_4698;
  wire [13:0] _GEN_4700 = 14'h125c == index ? 14'h24 : _GEN_4699;
  wire [13:0] _GEN_4701 = 14'h125d == index ? 14'h24 : _GEN_4700;
  wire [13:0] _GEN_4702 = 14'h125e == index ? 14'h24 : _GEN_4701;
  wire [13:0] _GEN_4703 = 14'h125f == index ? 14'h24 : _GEN_4702;
  wire [13:0] _GEN_4704 = 14'h1260 == index ? 14'h24 : _GEN_4703;
  wire [13:0] _GEN_4705 = 14'h1261 == index ? 14'h24 : _GEN_4704;
  wire [13:0] _GEN_4706 = 14'h1262 == index ? 14'h24 : _GEN_4705;
  wire [13:0] _GEN_4707 = 14'h1263 == index ? 14'h24 : _GEN_4706;
  wire [13:0] _GEN_4708 = 14'h1264 == index ? 14'h24 : _GEN_4707;
  wire [13:0] _GEN_4709 = 14'h1265 == index ? 14'h24 : _GEN_4708;
  wire [13:0] _GEN_4710 = 14'h1266 == index ? 14'h24 : _GEN_4709;
  wire [13:0] _GEN_4711 = 14'h1267 == index ? 14'h24 : _GEN_4710;
  wire [13:0] _GEN_4712 = 14'h1268 == index ? 14'h24 : _GEN_4711;
  wire [13:0] _GEN_4713 = 14'h1269 == index ? 14'h24 : _GEN_4712;
  wire [13:0] _GEN_4714 = 14'h126a == index ? 14'h24 : _GEN_4713;
  wire [13:0] _GEN_4715 = 14'h126b == index ? 14'h24 : _GEN_4714;
  wire [13:0] _GEN_4716 = 14'h126c == index ? 14'h24 : _GEN_4715;
  wire [13:0] _GEN_4717 = 14'h126d == index ? 14'h24 : _GEN_4716;
  wire [13:0] _GEN_4718 = 14'h126e == index ? 14'h24 : _GEN_4717;
  wire [13:0] _GEN_4719 = 14'h126f == index ? 14'h24 : _GEN_4718;
  wire [13:0] _GEN_4720 = 14'h1270 == index ? 14'h24 : _GEN_4719;
  wire [13:0] _GEN_4721 = 14'h1271 == index ? 14'h24 : _GEN_4720;
  wire [13:0] _GEN_4722 = 14'h1272 == index ? 14'h24 : _GEN_4721;
  wire [13:0] _GEN_4723 = 14'h1273 == index ? 14'h24 : _GEN_4722;
  wire [13:0] _GEN_4724 = 14'h1274 == index ? 14'h24 : _GEN_4723;
  wire [13:0] _GEN_4725 = 14'h1275 == index ? 14'h24 : _GEN_4724;
  wire [13:0] _GEN_4726 = 14'h1276 == index ? 14'h24 : _GEN_4725;
  wire [13:0] _GEN_4727 = 14'h1277 == index ? 14'h24 : _GEN_4726;
  wire [13:0] _GEN_4728 = 14'h1278 == index ? 14'h24 : _GEN_4727;
  wire [13:0] _GEN_4729 = 14'h1279 == index ? 14'h24 : _GEN_4728;
  wire [13:0] _GEN_4730 = 14'h127a == index ? 14'h24 : _GEN_4729;
  wire [13:0] _GEN_4731 = 14'h127b == index ? 14'h24 : _GEN_4730;
  wire [13:0] _GEN_4732 = 14'h127c == index ? 14'h24 : _GEN_4731;
  wire [13:0] _GEN_4733 = 14'h127d == index ? 14'h24 : _GEN_4732;
  wire [13:0] _GEN_4734 = 14'h127e == index ? 14'h24 : _GEN_4733;
  wire [13:0] _GEN_4735 = 14'h127f == index ? 14'h24 : _GEN_4734;
  wire [13:0] _GEN_4736 = 14'h1280 == index ? 14'h0 : _GEN_4735;
  wire [13:0] _GEN_4737 = 14'h1281 == index ? 14'h1280 : _GEN_4736;
  wire [13:0] _GEN_4738 = 14'h1282 == index ? 14'h901 : _GEN_4737;
  wire [13:0] _GEN_4739 = 14'h1283 == index ? 14'h601 : _GEN_4738;
  wire [13:0] _GEN_4740 = 14'h1284 == index ? 14'h481 : _GEN_4739;
  wire [13:0] _GEN_4741 = 14'h1285 == index ? 14'h382 : _GEN_4740;
  wire [13:0] _GEN_4742 = 14'h1286 == index ? 14'h301 : _GEN_4741;
  wire [13:0] _GEN_4743 = 14'h1287 == index ? 14'h282 : _GEN_4742;
  wire [13:0] _GEN_4744 = 14'h1288 == index ? 14'h205 : _GEN_4743;
  wire [13:0] _GEN_4745 = 14'h1289 == index ? 14'h201 : _GEN_4744;
  wire [13:0] _GEN_4746 = 14'h128a == index ? 14'h187 : _GEN_4745;
  wire [13:0] _GEN_4747 = 14'h128b == index ? 14'h184 : _GEN_4746;
  wire [13:0] _GEN_4748 = 14'h128c == index ? 14'h181 : _GEN_4747;
  wire [13:0] _GEN_4749 = 14'h128d == index ? 14'h10b : _GEN_4748;
  wire [13:0] _GEN_4750 = 14'h128e == index ? 14'h109 : _GEN_4749;
  wire [13:0] _GEN_4751 = 14'h128f == index ? 14'h107 : _GEN_4750;
  wire [13:0] _GEN_4752 = 14'h1290 == index ? 14'h105 : _GEN_4751;
  wire [13:0] _GEN_4753 = 14'h1291 == index ? 14'h103 : _GEN_4752;
  wire [13:0] _GEN_4754 = 14'h1292 == index ? 14'h101 : _GEN_4753;
  wire [13:0] _GEN_4755 = 14'h1293 == index ? 14'h92 : _GEN_4754;
  wire [13:0] _GEN_4756 = 14'h1294 == index ? 14'h91 : _GEN_4755;
  wire [13:0] _GEN_4757 = 14'h1295 == index ? 14'h90 : _GEN_4756;
  wire [13:0] _GEN_4758 = 14'h1296 == index ? 14'h8f : _GEN_4757;
  wire [13:0] _GEN_4759 = 14'h1297 == index ? 14'h8e : _GEN_4758;
  wire [13:0] _GEN_4760 = 14'h1298 == index ? 14'h8d : _GEN_4759;
  wire [13:0] _GEN_4761 = 14'h1299 == index ? 14'h8c : _GEN_4760;
  wire [13:0] _GEN_4762 = 14'h129a == index ? 14'h8b : _GEN_4761;
  wire [13:0] _GEN_4763 = 14'h129b == index ? 14'h8a : _GEN_4762;
  wire [13:0] _GEN_4764 = 14'h129c == index ? 14'h89 : _GEN_4763;
  wire [13:0] _GEN_4765 = 14'h129d == index ? 14'h88 : _GEN_4764;
  wire [13:0] _GEN_4766 = 14'h129e == index ? 14'h87 : _GEN_4765;
  wire [13:0] _GEN_4767 = 14'h129f == index ? 14'h86 : _GEN_4766;
  wire [13:0] _GEN_4768 = 14'h12a0 == index ? 14'h85 : _GEN_4767;
  wire [13:0] _GEN_4769 = 14'h12a1 == index ? 14'h84 : _GEN_4768;
  wire [13:0] _GEN_4770 = 14'h12a2 == index ? 14'h83 : _GEN_4769;
  wire [13:0] _GEN_4771 = 14'h12a3 == index ? 14'h82 : _GEN_4770;
  wire [13:0] _GEN_4772 = 14'h12a4 == index ? 14'h81 : _GEN_4771;
  wire [13:0] _GEN_4773 = 14'h12a5 == index ? 14'h80 : _GEN_4772;
  wire [13:0] _GEN_4774 = 14'h12a6 == index ? 14'h25 : _GEN_4773;
  wire [13:0] _GEN_4775 = 14'h12a7 == index ? 14'h25 : _GEN_4774;
  wire [13:0] _GEN_4776 = 14'h12a8 == index ? 14'h25 : _GEN_4775;
  wire [13:0] _GEN_4777 = 14'h12a9 == index ? 14'h25 : _GEN_4776;
  wire [13:0] _GEN_4778 = 14'h12aa == index ? 14'h25 : _GEN_4777;
  wire [13:0] _GEN_4779 = 14'h12ab == index ? 14'h25 : _GEN_4778;
  wire [13:0] _GEN_4780 = 14'h12ac == index ? 14'h25 : _GEN_4779;
  wire [13:0] _GEN_4781 = 14'h12ad == index ? 14'h25 : _GEN_4780;
  wire [13:0] _GEN_4782 = 14'h12ae == index ? 14'h25 : _GEN_4781;
  wire [13:0] _GEN_4783 = 14'h12af == index ? 14'h25 : _GEN_4782;
  wire [13:0] _GEN_4784 = 14'h12b0 == index ? 14'h25 : _GEN_4783;
  wire [13:0] _GEN_4785 = 14'h12b1 == index ? 14'h25 : _GEN_4784;
  wire [13:0] _GEN_4786 = 14'h12b2 == index ? 14'h25 : _GEN_4785;
  wire [13:0] _GEN_4787 = 14'h12b3 == index ? 14'h25 : _GEN_4786;
  wire [13:0] _GEN_4788 = 14'h12b4 == index ? 14'h25 : _GEN_4787;
  wire [13:0] _GEN_4789 = 14'h12b5 == index ? 14'h25 : _GEN_4788;
  wire [13:0] _GEN_4790 = 14'h12b6 == index ? 14'h25 : _GEN_4789;
  wire [13:0] _GEN_4791 = 14'h12b7 == index ? 14'h25 : _GEN_4790;
  wire [13:0] _GEN_4792 = 14'h12b8 == index ? 14'h25 : _GEN_4791;
  wire [13:0] _GEN_4793 = 14'h12b9 == index ? 14'h25 : _GEN_4792;
  wire [13:0] _GEN_4794 = 14'h12ba == index ? 14'h25 : _GEN_4793;
  wire [13:0] _GEN_4795 = 14'h12bb == index ? 14'h25 : _GEN_4794;
  wire [13:0] _GEN_4796 = 14'h12bc == index ? 14'h25 : _GEN_4795;
  wire [13:0] _GEN_4797 = 14'h12bd == index ? 14'h25 : _GEN_4796;
  wire [13:0] _GEN_4798 = 14'h12be == index ? 14'h25 : _GEN_4797;
  wire [13:0] _GEN_4799 = 14'h12bf == index ? 14'h25 : _GEN_4798;
  wire [13:0] _GEN_4800 = 14'h12c0 == index ? 14'h25 : _GEN_4799;
  wire [13:0] _GEN_4801 = 14'h12c1 == index ? 14'h25 : _GEN_4800;
  wire [13:0] _GEN_4802 = 14'h12c2 == index ? 14'h25 : _GEN_4801;
  wire [13:0] _GEN_4803 = 14'h12c3 == index ? 14'h25 : _GEN_4802;
  wire [13:0] _GEN_4804 = 14'h12c4 == index ? 14'h25 : _GEN_4803;
  wire [13:0] _GEN_4805 = 14'h12c5 == index ? 14'h25 : _GEN_4804;
  wire [13:0] _GEN_4806 = 14'h12c6 == index ? 14'h25 : _GEN_4805;
  wire [13:0] _GEN_4807 = 14'h12c7 == index ? 14'h25 : _GEN_4806;
  wire [13:0] _GEN_4808 = 14'h12c8 == index ? 14'h25 : _GEN_4807;
  wire [13:0] _GEN_4809 = 14'h12c9 == index ? 14'h25 : _GEN_4808;
  wire [13:0] _GEN_4810 = 14'h12ca == index ? 14'h25 : _GEN_4809;
  wire [13:0] _GEN_4811 = 14'h12cb == index ? 14'h25 : _GEN_4810;
  wire [13:0] _GEN_4812 = 14'h12cc == index ? 14'h25 : _GEN_4811;
  wire [13:0] _GEN_4813 = 14'h12cd == index ? 14'h25 : _GEN_4812;
  wire [13:0] _GEN_4814 = 14'h12ce == index ? 14'h25 : _GEN_4813;
  wire [13:0] _GEN_4815 = 14'h12cf == index ? 14'h25 : _GEN_4814;
  wire [13:0] _GEN_4816 = 14'h12d0 == index ? 14'h25 : _GEN_4815;
  wire [13:0] _GEN_4817 = 14'h12d1 == index ? 14'h25 : _GEN_4816;
  wire [13:0] _GEN_4818 = 14'h12d2 == index ? 14'h25 : _GEN_4817;
  wire [13:0] _GEN_4819 = 14'h12d3 == index ? 14'h25 : _GEN_4818;
  wire [13:0] _GEN_4820 = 14'h12d4 == index ? 14'h25 : _GEN_4819;
  wire [13:0] _GEN_4821 = 14'h12d5 == index ? 14'h25 : _GEN_4820;
  wire [13:0] _GEN_4822 = 14'h12d6 == index ? 14'h25 : _GEN_4821;
  wire [13:0] _GEN_4823 = 14'h12d7 == index ? 14'h25 : _GEN_4822;
  wire [13:0] _GEN_4824 = 14'h12d8 == index ? 14'h25 : _GEN_4823;
  wire [13:0] _GEN_4825 = 14'h12d9 == index ? 14'h25 : _GEN_4824;
  wire [13:0] _GEN_4826 = 14'h12da == index ? 14'h25 : _GEN_4825;
  wire [13:0] _GEN_4827 = 14'h12db == index ? 14'h25 : _GEN_4826;
  wire [13:0] _GEN_4828 = 14'h12dc == index ? 14'h25 : _GEN_4827;
  wire [13:0] _GEN_4829 = 14'h12dd == index ? 14'h25 : _GEN_4828;
  wire [13:0] _GEN_4830 = 14'h12de == index ? 14'h25 : _GEN_4829;
  wire [13:0] _GEN_4831 = 14'h12df == index ? 14'h25 : _GEN_4830;
  wire [13:0] _GEN_4832 = 14'h12e0 == index ? 14'h25 : _GEN_4831;
  wire [13:0] _GEN_4833 = 14'h12e1 == index ? 14'h25 : _GEN_4832;
  wire [13:0] _GEN_4834 = 14'h12e2 == index ? 14'h25 : _GEN_4833;
  wire [13:0] _GEN_4835 = 14'h12e3 == index ? 14'h25 : _GEN_4834;
  wire [13:0] _GEN_4836 = 14'h12e4 == index ? 14'h25 : _GEN_4835;
  wire [13:0] _GEN_4837 = 14'h12e5 == index ? 14'h25 : _GEN_4836;
  wire [13:0] _GEN_4838 = 14'h12e6 == index ? 14'h25 : _GEN_4837;
  wire [13:0] _GEN_4839 = 14'h12e7 == index ? 14'h25 : _GEN_4838;
  wire [13:0] _GEN_4840 = 14'h12e8 == index ? 14'h25 : _GEN_4839;
  wire [13:0] _GEN_4841 = 14'h12e9 == index ? 14'h25 : _GEN_4840;
  wire [13:0] _GEN_4842 = 14'h12ea == index ? 14'h25 : _GEN_4841;
  wire [13:0] _GEN_4843 = 14'h12eb == index ? 14'h25 : _GEN_4842;
  wire [13:0] _GEN_4844 = 14'h12ec == index ? 14'h25 : _GEN_4843;
  wire [13:0] _GEN_4845 = 14'h12ed == index ? 14'h25 : _GEN_4844;
  wire [13:0] _GEN_4846 = 14'h12ee == index ? 14'h25 : _GEN_4845;
  wire [13:0] _GEN_4847 = 14'h12ef == index ? 14'h25 : _GEN_4846;
  wire [13:0] _GEN_4848 = 14'h12f0 == index ? 14'h25 : _GEN_4847;
  wire [13:0] _GEN_4849 = 14'h12f1 == index ? 14'h25 : _GEN_4848;
  wire [13:0] _GEN_4850 = 14'h12f2 == index ? 14'h25 : _GEN_4849;
  wire [13:0] _GEN_4851 = 14'h12f3 == index ? 14'h25 : _GEN_4850;
  wire [13:0] _GEN_4852 = 14'h12f4 == index ? 14'h25 : _GEN_4851;
  wire [13:0] _GEN_4853 = 14'h12f5 == index ? 14'h25 : _GEN_4852;
  wire [13:0] _GEN_4854 = 14'h12f6 == index ? 14'h25 : _GEN_4853;
  wire [13:0] _GEN_4855 = 14'h12f7 == index ? 14'h25 : _GEN_4854;
  wire [13:0] _GEN_4856 = 14'h12f8 == index ? 14'h25 : _GEN_4855;
  wire [13:0] _GEN_4857 = 14'h12f9 == index ? 14'h25 : _GEN_4856;
  wire [13:0] _GEN_4858 = 14'h12fa == index ? 14'h25 : _GEN_4857;
  wire [13:0] _GEN_4859 = 14'h12fb == index ? 14'h25 : _GEN_4858;
  wire [13:0] _GEN_4860 = 14'h12fc == index ? 14'h25 : _GEN_4859;
  wire [13:0] _GEN_4861 = 14'h12fd == index ? 14'h25 : _GEN_4860;
  wire [13:0] _GEN_4862 = 14'h12fe == index ? 14'h25 : _GEN_4861;
  wire [13:0] _GEN_4863 = 14'h12ff == index ? 14'h25 : _GEN_4862;
  wire [13:0] _GEN_4864 = 14'h1300 == index ? 14'h0 : _GEN_4863;
  wire [13:0] _GEN_4865 = 14'h1301 == index ? 14'h1300 : _GEN_4864;
  wire [13:0] _GEN_4866 = 14'h1302 == index ? 14'h980 : _GEN_4865;
  wire [13:0] _GEN_4867 = 14'h1303 == index ? 14'h602 : _GEN_4866;
  wire [13:0] _GEN_4868 = 14'h1304 == index ? 14'h482 : _GEN_4867;
  wire [13:0] _GEN_4869 = 14'h1305 == index ? 14'h383 : _GEN_4868;
  wire [13:0] _GEN_4870 = 14'h1306 == index ? 14'h302 : _GEN_4869;
  wire [13:0] _GEN_4871 = 14'h1307 == index ? 14'h283 : _GEN_4870;
  wire [13:0] _GEN_4872 = 14'h1308 == index ? 14'h206 : _GEN_4871;
  wire [13:0] _GEN_4873 = 14'h1309 == index ? 14'h202 : _GEN_4872;
  wire [13:0] _GEN_4874 = 14'h130a == index ? 14'h188 : _GEN_4873;
  wire [13:0] _GEN_4875 = 14'h130b == index ? 14'h185 : _GEN_4874;
  wire [13:0] _GEN_4876 = 14'h130c == index ? 14'h182 : _GEN_4875;
  wire [13:0] _GEN_4877 = 14'h130d == index ? 14'h10c : _GEN_4876;
  wire [13:0] _GEN_4878 = 14'h130e == index ? 14'h10a : _GEN_4877;
  wire [13:0] _GEN_4879 = 14'h130f == index ? 14'h108 : _GEN_4878;
  wire [13:0] _GEN_4880 = 14'h1310 == index ? 14'h106 : _GEN_4879;
  wire [13:0] _GEN_4881 = 14'h1311 == index ? 14'h104 : _GEN_4880;
  wire [13:0] _GEN_4882 = 14'h1312 == index ? 14'h102 : _GEN_4881;
  wire [13:0] _GEN_4883 = 14'h1313 == index ? 14'h100 : _GEN_4882;
  wire [13:0] _GEN_4884 = 14'h1314 == index ? 14'h92 : _GEN_4883;
  wire [13:0] _GEN_4885 = 14'h1315 == index ? 14'h91 : _GEN_4884;
  wire [13:0] _GEN_4886 = 14'h1316 == index ? 14'h90 : _GEN_4885;
  wire [13:0] _GEN_4887 = 14'h1317 == index ? 14'h8f : _GEN_4886;
  wire [13:0] _GEN_4888 = 14'h1318 == index ? 14'h8e : _GEN_4887;
  wire [13:0] _GEN_4889 = 14'h1319 == index ? 14'h8d : _GEN_4888;
  wire [13:0] _GEN_4890 = 14'h131a == index ? 14'h8c : _GEN_4889;
  wire [13:0] _GEN_4891 = 14'h131b == index ? 14'h8b : _GEN_4890;
  wire [13:0] _GEN_4892 = 14'h131c == index ? 14'h8a : _GEN_4891;
  wire [13:0] _GEN_4893 = 14'h131d == index ? 14'h89 : _GEN_4892;
  wire [13:0] _GEN_4894 = 14'h131e == index ? 14'h88 : _GEN_4893;
  wire [13:0] _GEN_4895 = 14'h131f == index ? 14'h87 : _GEN_4894;
  wire [13:0] _GEN_4896 = 14'h1320 == index ? 14'h86 : _GEN_4895;
  wire [13:0] _GEN_4897 = 14'h1321 == index ? 14'h85 : _GEN_4896;
  wire [13:0] _GEN_4898 = 14'h1322 == index ? 14'h84 : _GEN_4897;
  wire [13:0] _GEN_4899 = 14'h1323 == index ? 14'h83 : _GEN_4898;
  wire [13:0] _GEN_4900 = 14'h1324 == index ? 14'h82 : _GEN_4899;
  wire [13:0] _GEN_4901 = 14'h1325 == index ? 14'h81 : _GEN_4900;
  wire [13:0] _GEN_4902 = 14'h1326 == index ? 14'h80 : _GEN_4901;
  wire [13:0] _GEN_4903 = 14'h1327 == index ? 14'h26 : _GEN_4902;
  wire [13:0] _GEN_4904 = 14'h1328 == index ? 14'h26 : _GEN_4903;
  wire [13:0] _GEN_4905 = 14'h1329 == index ? 14'h26 : _GEN_4904;
  wire [13:0] _GEN_4906 = 14'h132a == index ? 14'h26 : _GEN_4905;
  wire [13:0] _GEN_4907 = 14'h132b == index ? 14'h26 : _GEN_4906;
  wire [13:0] _GEN_4908 = 14'h132c == index ? 14'h26 : _GEN_4907;
  wire [13:0] _GEN_4909 = 14'h132d == index ? 14'h26 : _GEN_4908;
  wire [13:0] _GEN_4910 = 14'h132e == index ? 14'h26 : _GEN_4909;
  wire [13:0] _GEN_4911 = 14'h132f == index ? 14'h26 : _GEN_4910;
  wire [13:0] _GEN_4912 = 14'h1330 == index ? 14'h26 : _GEN_4911;
  wire [13:0] _GEN_4913 = 14'h1331 == index ? 14'h26 : _GEN_4912;
  wire [13:0] _GEN_4914 = 14'h1332 == index ? 14'h26 : _GEN_4913;
  wire [13:0] _GEN_4915 = 14'h1333 == index ? 14'h26 : _GEN_4914;
  wire [13:0] _GEN_4916 = 14'h1334 == index ? 14'h26 : _GEN_4915;
  wire [13:0] _GEN_4917 = 14'h1335 == index ? 14'h26 : _GEN_4916;
  wire [13:0] _GEN_4918 = 14'h1336 == index ? 14'h26 : _GEN_4917;
  wire [13:0] _GEN_4919 = 14'h1337 == index ? 14'h26 : _GEN_4918;
  wire [13:0] _GEN_4920 = 14'h1338 == index ? 14'h26 : _GEN_4919;
  wire [13:0] _GEN_4921 = 14'h1339 == index ? 14'h26 : _GEN_4920;
  wire [13:0] _GEN_4922 = 14'h133a == index ? 14'h26 : _GEN_4921;
  wire [13:0] _GEN_4923 = 14'h133b == index ? 14'h26 : _GEN_4922;
  wire [13:0] _GEN_4924 = 14'h133c == index ? 14'h26 : _GEN_4923;
  wire [13:0] _GEN_4925 = 14'h133d == index ? 14'h26 : _GEN_4924;
  wire [13:0] _GEN_4926 = 14'h133e == index ? 14'h26 : _GEN_4925;
  wire [13:0] _GEN_4927 = 14'h133f == index ? 14'h26 : _GEN_4926;
  wire [13:0] _GEN_4928 = 14'h1340 == index ? 14'h26 : _GEN_4927;
  wire [13:0] _GEN_4929 = 14'h1341 == index ? 14'h26 : _GEN_4928;
  wire [13:0] _GEN_4930 = 14'h1342 == index ? 14'h26 : _GEN_4929;
  wire [13:0] _GEN_4931 = 14'h1343 == index ? 14'h26 : _GEN_4930;
  wire [13:0] _GEN_4932 = 14'h1344 == index ? 14'h26 : _GEN_4931;
  wire [13:0] _GEN_4933 = 14'h1345 == index ? 14'h26 : _GEN_4932;
  wire [13:0] _GEN_4934 = 14'h1346 == index ? 14'h26 : _GEN_4933;
  wire [13:0] _GEN_4935 = 14'h1347 == index ? 14'h26 : _GEN_4934;
  wire [13:0] _GEN_4936 = 14'h1348 == index ? 14'h26 : _GEN_4935;
  wire [13:0] _GEN_4937 = 14'h1349 == index ? 14'h26 : _GEN_4936;
  wire [13:0] _GEN_4938 = 14'h134a == index ? 14'h26 : _GEN_4937;
  wire [13:0] _GEN_4939 = 14'h134b == index ? 14'h26 : _GEN_4938;
  wire [13:0] _GEN_4940 = 14'h134c == index ? 14'h26 : _GEN_4939;
  wire [13:0] _GEN_4941 = 14'h134d == index ? 14'h26 : _GEN_4940;
  wire [13:0] _GEN_4942 = 14'h134e == index ? 14'h26 : _GEN_4941;
  wire [13:0] _GEN_4943 = 14'h134f == index ? 14'h26 : _GEN_4942;
  wire [13:0] _GEN_4944 = 14'h1350 == index ? 14'h26 : _GEN_4943;
  wire [13:0] _GEN_4945 = 14'h1351 == index ? 14'h26 : _GEN_4944;
  wire [13:0] _GEN_4946 = 14'h1352 == index ? 14'h26 : _GEN_4945;
  wire [13:0] _GEN_4947 = 14'h1353 == index ? 14'h26 : _GEN_4946;
  wire [13:0] _GEN_4948 = 14'h1354 == index ? 14'h26 : _GEN_4947;
  wire [13:0] _GEN_4949 = 14'h1355 == index ? 14'h26 : _GEN_4948;
  wire [13:0] _GEN_4950 = 14'h1356 == index ? 14'h26 : _GEN_4949;
  wire [13:0] _GEN_4951 = 14'h1357 == index ? 14'h26 : _GEN_4950;
  wire [13:0] _GEN_4952 = 14'h1358 == index ? 14'h26 : _GEN_4951;
  wire [13:0] _GEN_4953 = 14'h1359 == index ? 14'h26 : _GEN_4952;
  wire [13:0] _GEN_4954 = 14'h135a == index ? 14'h26 : _GEN_4953;
  wire [13:0] _GEN_4955 = 14'h135b == index ? 14'h26 : _GEN_4954;
  wire [13:0] _GEN_4956 = 14'h135c == index ? 14'h26 : _GEN_4955;
  wire [13:0] _GEN_4957 = 14'h135d == index ? 14'h26 : _GEN_4956;
  wire [13:0] _GEN_4958 = 14'h135e == index ? 14'h26 : _GEN_4957;
  wire [13:0] _GEN_4959 = 14'h135f == index ? 14'h26 : _GEN_4958;
  wire [13:0] _GEN_4960 = 14'h1360 == index ? 14'h26 : _GEN_4959;
  wire [13:0] _GEN_4961 = 14'h1361 == index ? 14'h26 : _GEN_4960;
  wire [13:0] _GEN_4962 = 14'h1362 == index ? 14'h26 : _GEN_4961;
  wire [13:0] _GEN_4963 = 14'h1363 == index ? 14'h26 : _GEN_4962;
  wire [13:0] _GEN_4964 = 14'h1364 == index ? 14'h26 : _GEN_4963;
  wire [13:0] _GEN_4965 = 14'h1365 == index ? 14'h26 : _GEN_4964;
  wire [13:0] _GEN_4966 = 14'h1366 == index ? 14'h26 : _GEN_4965;
  wire [13:0] _GEN_4967 = 14'h1367 == index ? 14'h26 : _GEN_4966;
  wire [13:0] _GEN_4968 = 14'h1368 == index ? 14'h26 : _GEN_4967;
  wire [13:0] _GEN_4969 = 14'h1369 == index ? 14'h26 : _GEN_4968;
  wire [13:0] _GEN_4970 = 14'h136a == index ? 14'h26 : _GEN_4969;
  wire [13:0] _GEN_4971 = 14'h136b == index ? 14'h26 : _GEN_4970;
  wire [13:0] _GEN_4972 = 14'h136c == index ? 14'h26 : _GEN_4971;
  wire [13:0] _GEN_4973 = 14'h136d == index ? 14'h26 : _GEN_4972;
  wire [13:0] _GEN_4974 = 14'h136e == index ? 14'h26 : _GEN_4973;
  wire [13:0] _GEN_4975 = 14'h136f == index ? 14'h26 : _GEN_4974;
  wire [13:0] _GEN_4976 = 14'h1370 == index ? 14'h26 : _GEN_4975;
  wire [13:0] _GEN_4977 = 14'h1371 == index ? 14'h26 : _GEN_4976;
  wire [13:0] _GEN_4978 = 14'h1372 == index ? 14'h26 : _GEN_4977;
  wire [13:0] _GEN_4979 = 14'h1373 == index ? 14'h26 : _GEN_4978;
  wire [13:0] _GEN_4980 = 14'h1374 == index ? 14'h26 : _GEN_4979;
  wire [13:0] _GEN_4981 = 14'h1375 == index ? 14'h26 : _GEN_4980;
  wire [13:0] _GEN_4982 = 14'h1376 == index ? 14'h26 : _GEN_4981;
  wire [13:0] _GEN_4983 = 14'h1377 == index ? 14'h26 : _GEN_4982;
  wire [13:0] _GEN_4984 = 14'h1378 == index ? 14'h26 : _GEN_4983;
  wire [13:0] _GEN_4985 = 14'h1379 == index ? 14'h26 : _GEN_4984;
  wire [13:0] _GEN_4986 = 14'h137a == index ? 14'h26 : _GEN_4985;
  wire [13:0] _GEN_4987 = 14'h137b == index ? 14'h26 : _GEN_4986;
  wire [13:0] _GEN_4988 = 14'h137c == index ? 14'h26 : _GEN_4987;
  wire [13:0] _GEN_4989 = 14'h137d == index ? 14'h26 : _GEN_4988;
  wire [13:0] _GEN_4990 = 14'h137e == index ? 14'h26 : _GEN_4989;
  wire [13:0] _GEN_4991 = 14'h137f == index ? 14'h26 : _GEN_4990;
  wire [13:0] _GEN_4992 = 14'h1380 == index ? 14'h0 : _GEN_4991;
  wire [13:0] _GEN_4993 = 14'h1381 == index ? 14'h1380 : _GEN_4992;
  wire [13:0] _GEN_4994 = 14'h1382 == index ? 14'h981 : _GEN_4993;
  wire [13:0] _GEN_4995 = 14'h1383 == index ? 14'h680 : _GEN_4994;
  wire [13:0] _GEN_4996 = 14'h1384 == index ? 14'h483 : _GEN_4995;
  wire [13:0] _GEN_4997 = 14'h1385 == index ? 14'h384 : _GEN_4996;
  wire [13:0] _GEN_4998 = 14'h1386 == index ? 14'h303 : _GEN_4997;
  wire [13:0] _GEN_4999 = 14'h1387 == index ? 14'h284 : _GEN_4998;
  wire [13:0] _GEN_5000 = 14'h1388 == index ? 14'h207 : _GEN_4999;
  wire [13:0] _GEN_5001 = 14'h1389 == index ? 14'h203 : _GEN_5000;
  wire [13:0] _GEN_5002 = 14'h138a == index ? 14'h189 : _GEN_5001;
  wire [13:0] _GEN_5003 = 14'h138b == index ? 14'h186 : _GEN_5002;
  wire [13:0] _GEN_5004 = 14'h138c == index ? 14'h183 : _GEN_5003;
  wire [13:0] _GEN_5005 = 14'h138d == index ? 14'h180 : _GEN_5004;
  wire [13:0] _GEN_5006 = 14'h138e == index ? 14'h10b : _GEN_5005;
  wire [13:0] _GEN_5007 = 14'h138f == index ? 14'h109 : _GEN_5006;
  wire [13:0] _GEN_5008 = 14'h1390 == index ? 14'h107 : _GEN_5007;
  wire [13:0] _GEN_5009 = 14'h1391 == index ? 14'h105 : _GEN_5008;
  wire [13:0] _GEN_5010 = 14'h1392 == index ? 14'h103 : _GEN_5009;
  wire [13:0] _GEN_5011 = 14'h1393 == index ? 14'h101 : _GEN_5010;
  wire [13:0] _GEN_5012 = 14'h1394 == index ? 14'h93 : _GEN_5011;
  wire [13:0] _GEN_5013 = 14'h1395 == index ? 14'h92 : _GEN_5012;
  wire [13:0] _GEN_5014 = 14'h1396 == index ? 14'h91 : _GEN_5013;
  wire [13:0] _GEN_5015 = 14'h1397 == index ? 14'h90 : _GEN_5014;
  wire [13:0] _GEN_5016 = 14'h1398 == index ? 14'h8f : _GEN_5015;
  wire [13:0] _GEN_5017 = 14'h1399 == index ? 14'h8e : _GEN_5016;
  wire [13:0] _GEN_5018 = 14'h139a == index ? 14'h8d : _GEN_5017;
  wire [13:0] _GEN_5019 = 14'h139b == index ? 14'h8c : _GEN_5018;
  wire [13:0] _GEN_5020 = 14'h139c == index ? 14'h8b : _GEN_5019;
  wire [13:0] _GEN_5021 = 14'h139d == index ? 14'h8a : _GEN_5020;
  wire [13:0] _GEN_5022 = 14'h139e == index ? 14'h89 : _GEN_5021;
  wire [13:0] _GEN_5023 = 14'h139f == index ? 14'h88 : _GEN_5022;
  wire [13:0] _GEN_5024 = 14'h13a0 == index ? 14'h87 : _GEN_5023;
  wire [13:0] _GEN_5025 = 14'h13a1 == index ? 14'h86 : _GEN_5024;
  wire [13:0] _GEN_5026 = 14'h13a2 == index ? 14'h85 : _GEN_5025;
  wire [13:0] _GEN_5027 = 14'h13a3 == index ? 14'h84 : _GEN_5026;
  wire [13:0] _GEN_5028 = 14'h13a4 == index ? 14'h83 : _GEN_5027;
  wire [13:0] _GEN_5029 = 14'h13a5 == index ? 14'h82 : _GEN_5028;
  wire [13:0] _GEN_5030 = 14'h13a6 == index ? 14'h81 : _GEN_5029;
  wire [13:0] _GEN_5031 = 14'h13a7 == index ? 14'h80 : _GEN_5030;
  wire [13:0] _GEN_5032 = 14'h13a8 == index ? 14'h27 : _GEN_5031;
  wire [13:0] _GEN_5033 = 14'h13a9 == index ? 14'h27 : _GEN_5032;
  wire [13:0] _GEN_5034 = 14'h13aa == index ? 14'h27 : _GEN_5033;
  wire [13:0] _GEN_5035 = 14'h13ab == index ? 14'h27 : _GEN_5034;
  wire [13:0] _GEN_5036 = 14'h13ac == index ? 14'h27 : _GEN_5035;
  wire [13:0] _GEN_5037 = 14'h13ad == index ? 14'h27 : _GEN_5036;
  wire [13:0] _GEN_5038 = 14'h13ae == index ? 14'h27 : _GEN_5037;
  wire [13:0] _GEN_5039 = 14'h13af == index ? 14'h27 : _GEN_5038;
  wire [13:0] _GEN_5040 = 14'h13b0 == index ? 14'h27 : _GEN_5039;
  wire [13:0] _GEN_5041 = 14'h13b1 == index ? 14'h27 : _GEN_5040;
  wire [13:0] _GEN_5042 = 14'h13b2 == index ? 14'h27 : _GEN_5041;
  wire [13:0] _GEN_5043 = 14'h13b3 == index ? 14'h27 : _GEN_5042;
  wire [13:0] _GEN_5044 = 14'h13b4 == index ? 14'h27 : _GEN_5043;
  wire [13:0] _GEN_5045 = 14'h13b5 == index ? 14'h27 : _GEN_5044;
  wire [13:0] _GEN_5046 = 14'h13b6 == index ? 14'h27 : _GEN_5045;
  wire [13:0] _GEN_5047 = 14'h13b7 == index ? 14'h27 : _GEN_5046;
  wire [13:0] _GEN_5048 = 14'h13b8 == index ? 14'h27 : _GEN_5047;
  wire [13:0] _GEN_5049 = 14'h13b9 == index ? 14'h27 : _GEN_5048;
  wire [13:0] _GEN_5050 = 14'h13ba == index ? 14'h27 : _GEN_5049;
  wire [13:0] _GEN_5051 = 14'h13bb == index ? 14'h27 : _GEN_5050;
  wire [13:0] _GEN_5052 = 14'h13bc == index ? 14'h27 : _GEN_5051;
  wire [13:0] _GEN_5053 = 14'h13bd == index ? 14'h27 : _GEN_5052;
  wire [13:0] _GEN_5054 = 14'h13be == index ? 14'h27 : _GEN_5053;
  wire [13:0] _GEN_5055 = 14'h13bf == index ? 14'h27 : _GEN_5054;
  wire [13:0] _GEN_5056 = 14'h13c0 == index ? 14'h27 : _GEN_5055;
  wire [13:0] _GEN_5057 = 14'h13c1 == index ? 14'h27 : _GEN_5056;
  wire [13:0] _GEN_5058 = 14'h13c2 == index ? 14'h27 : _GEN_5057;
  wire [13:0] _GEN_5059 = 14'h13c3 == index ? 14'h27 : _GEN_5058;
  wire [13:0] _GEN_5060 = 14'h13c4 == index ? 14'h27 : _GEN_5059;
  wire [13:0] _GEN_5061 = 14'h13c5 == index ? 14'h27 : _GEN_5060;
  wire [13:0] _GEN_5062 = 14'h13c6 == index ? 14'h27 : _GEN_5061;
  wire [13:0] _GEN_5063 = 14'h13c7 == index ? 14'h27 : _GEN_5062;
  wire [13:0] _GEN_5064 = 14'h13c8 == index ? 14'h27 : _GEN_5063;
  wire [13:0] _GEN_5065 = 14'h13c9 == index ? 14'h27 : _GEN_5064;
  wire [13:0] _GEN_5066 = 14'h13ca == index ? 14'h27 : _GEN_5065;
  wire [13:0] _GEN_5067 = 14'h13cb == index ? 14'h27 : _GEN_5066;
  wire [13:0] _GEN_5068 = 14'h13cc == index ? 14'h27 : _GEN_5067;
  wire [13:0] _GEN_5069 = 14'h13cd == index ? 14'h27 : _GEN_5068;
  wire [13:0] _GEN_5070 = 14'h13ce == index ? 14'h27 : _GEN_5069;
  wire [13:0] _GEN_5071 = 14'h13cf == index ? 14'h27 : _GEN_5070;
  wire [13:0] _GEN_5072 = 14'h13d0 == index ? 14'h27 : _GEN_5071;
  wire [13:0] _GEN_5073 = 14'h13d1 == index ? 14'h27 : _GEN_5072;
  wire [13:0] _GEN_5074 = 14'h13d2 == index ? 14'h27 : _GEN_5073;
  wire [13:0] _GEN_5075 = 14'h13d3 == index ? 14'h27 : _GEN_5074;
  wire [13:0] _GEN_5076 = 14'h13d4 == index ? 14'h27 : _GEN_5075;
  wire [13:0] _GEN_5077 = 14'h13d5 == index ? 14'h27 : _GEN_5076;
  wire [13:0] _GEN_5078 = 14'h13d6 == index ? 14'h27 : _GEN_5077;
  wire [13:0] _GEN_5079 = 14'h13d7 == index ? 14'h27 : _GEN_5078;
  wire [13:0] _GEN_5080 = 14'h13d8 == index ? 14'h27 : _GEN_5079;
  wire [13:0] _GEN_5081 = 14'h13d9 == index ? 14'h27 : _GEN_5080;
  wire [13:0] _GEN_5082 = 14'h13da == index ? 14'h27 : _GEN_5081;
  wire [13:0] _GEN_5083 = 14'h13db == index ? 14'h27 : _GEN_5082;
  wire [13:0] _GEN_5084 = 14'h13dc == index ? 14'h27 : _GEN_5083;
  wire [13:0] _GEN_5085 = 14'h13dd == index ? 14'h27 : _GEN_5084;
  wire [13:0] _GEN_5086 = 14'h13de == index ? 14'h27 : _GEN_5085;
  wire [13:0] _GEN_5087 = 14'h13df == index ? 14'h27 : _GEN_5086;
  wire [13:0] _GEN_5088 = 14'h13e0 == index ? 14'h27 : _GEN_5087;
  wire [13:0] _GEN_5089 = 14'h13e1 == index ? 14'h27 : _GEN_5088;
  wire [13:0] _GEN_5090 = 14'h13e2 == index ? 14'h27 : _GEN_5089;
  wire [13:0] _GEN_5091 = 14'h13e3 == index ? 14'h27 : _GEN_5090;
  wire [13:0] _GEN_5092 = 14'h13e4 == index ? 14'h27 : _GEN_5091;
  wire [13:0] _GEN_5093 = 14'h13e5 == index ? 14'h27 : _GEN_5092;
  wire [13:0] _GEN_5094 = 14'h13e6 == index ? 14'h27 : _GEN_5093;
  wire [13:0] _GEN_5095 = 14'h13e7 == index ? 14'h27 : _GEN_5094;
  wire [13:0] _GEN_5096 = 14'h13e8 == index ? 14'h27 : _GEN_5095;
  wire [13:0] _GEN_5097 = 14'h13e9 == index ? 14'h27 : _GEN_5096;
  wire [13:0] _GEN_5098 = 14'h13ea == index ? 14'h27 : _GEN_5097;
  wire [13:0] _GEN_5099 = 14'h13eb == index ? 14'h27 : _GEN_5098;
  wire [13:0] _GEN_5100 = 14'h13ec == index ? 14'h27 : _GEN_5099;
  wire [13:0] _GEN_5101 = 14'h13ed == index ? 14'h27 : _GEN_5100;
  wire [13:0] _GEN_5102 = 14'h13ee == index ? 14'h27 : _GEN_5101;
  wire [13:0] _GEN_5103 = 14'h13ef == index ? 14'h27 : _GEN_5102;
  wire [13:0] _GEN_5104 = 14'h13f0 == index ? 14'h27 : _GEN_5103;
  wire [13:0] _GEN_5105 = 14'h13f1 == index ? 14'h27 : _GEN_5104;
  wire [13:0] _GEN_5106 = 14'h13f2 == index ? 14'h27 : _GEN_5105;
  wire [13:0] _GEN_5107 = 14'h13f3 == index ? 14'h27 : _GEN_5106;
  wire [13:0] _GEN_5108 = 14'h13f4 == index ? 14'h27 : _GEN_5107;
  wire [13:0] _GEN_5109 = 14'h13f5 == index ? 14'h27 : _GEN_5108;
  wire [13:0] _GEN_5110 = 14'h13f6 == index ? 14'h27 : _GEN_5109;
  wire [13:0] _GEN_5111 = 14'h13f7 == index ? 14'h27 : _GEN_5110;
  wire [13:0] _GEN_5112 = 14'h13f8 == index ? 14'h27 : _GEN_5111;
  wire [13:0] _GEN_5113 = 14'h13f9 == index ? 14'h27 : _GEN_5112;
  wire [13:0] _GEN_5114 = 14'h13fa == index ? 14'h27 : _GEN_5113;
  wire [13:0] _GEN_5115 = 14'h13fb == index ? 14'h27 : _GEN_5114;
  wire [13:0] _GEN_5116 = 14'h13fc == index ? 14'h27 : _GEN_5115;
  wire [13:0] _GEN_5117 = 14'h13fd == index ? 14'h27 : _GEN_5116;
  wire [13:0] _GEN_5118 = 14'h13fe == index ? 14'h27 : _GEN_5117;
  wire [13:0] _GEN_5119 = 14'h13ff == index ? 14'h27 : _GEN_5118;
  wire [13:0] _GEN_5120 = 14'h1400 == index ? 14'h0 : _GEN_5119;
  wire [13:0] _GEN_5121 = 14'h1401 == index ? 14'h1400 : _GEN_5120;
  wire [13:0] _GEN_5122 = 14'h1402 == index ? 14'ha00 : _GEN_5121;
  wire [13:0] _GEN_5123 = 14'h1403 == index ? 14'h681 : _GEN_5122;
  wire [13:0] _GEN_5124 = 14'h1404 == index ? 14'h500 : _GEN_5123;
  wire [13:0] _GEN_5125 = 14'h1405 == index ? 14'h400 : _GEN_5124;
  wire [13:0] _GEN_5126 = 14'h1406 == index ? 14'h304 : _GEN_5125;
  wire [13:0] _GEN_5127 = 14'h1407 == index ? 14'h285 : _GEN_5126;
  wire [13:0] _GEN_5128 = 14'h1408 == index ? 14'h280 : _GEN_5127;
  wire [13:0] _GEN_5129 = 14'h1409 == index ? 14'h204 : _GEN_5128;
  wire [13:0] _GEN_5130 = 14'h140a == index ? 14'h200 : _GEN_5129;
  wire [13:0] _GEN_5131 = 14'h140b == index ? 14'h187 : _GEN_5130;
  wire [13:0] _GEN_5132 = 14'h140c == index ? 14'h184 : _GEN_5131;
  wire [13:0] _GEN_5133 = 14'h140d == index ? 14'h181 : _GEN_5132;
  wire [13:0] _GEN_5134 = 14'h140e == index ? 14'h10c : _GEN_5133;
  wire [13:0] _GEN_5135 = 14'h140f == index ? 14'h10a : _GEN_5134;
  wire [13:0] _GEN_5136 = 14'h1410 == index ? 14'h108 : _GEN_5135;
  wire [13:0] _GEN_5137 = 14'h1411 == index ? 14'h106 : _GEN_5136;
  wire [13:0] _GEN_5138 = 14'h1412 == index ? 14'h104 : _GEN_5137;
  wire [13:0] _GEN_5139 = 14'h1413 == index ? 14'h102 : _GEN_5138;
  wire [13:0] _GEN_5140 = 14'h1414 == index ? 14'h100 : _GEN_5139;
  wire [13:0] _GEN_5141 = 14'h1415 == index ? 14'h93 : _GEN_5140;
  wire [13:0] _GEN_5142 = 14'h1416 == index ? 14'h92 : _GEN_5141;
  wire [13:0] _GEN_5143 = 14'h1417 == index ? 14'h91 : _GEN_5142;
  wire [13:0] _GEN_5144 = 14'h1418 == index ? 14'h90 : _GEN_5143;
  wire [13:0] _GEN_5145 = 14'h1419 == index ? 14'h8f : _GEN_5144;
  wire [13:0] _GEN_5146 = 14'h141a == index ? 14'h8e : _GEN_5145;
  wire [13:0] _GEN_5147 = 14'h141b == index ? 14'h8d : _GEN_5146;
  wire [13:0] _GEN_5148 = 14'h141c == index ? 14'h8c : _GEN_5147;
  wire [13:0] _GEN_5149 = 14'h141d == index ? 14'h8b : _GEN_5148;
  wire [13:0] _GEN_5150 = 14'h141e == index ? 14'h8a : _GEN_5149;
  wire [13:0] _GEN_5151 = 14'h141f == index ? 14'h89 : _GEN_5150;
  wire [13:0] _GEN_5152 = 14'h1420 == index ? 14'h88 : _GEN_5151;
  wire [13:0] _GEN_5153 = 14'h1421 == index ? 14'h87 : _GEN_5152;
  wire [13:0] _GEN_5154 = 14'h1422 == index ? 14'h86 : _GEN_5153;
  wire [13:0] _GEN_5155 = 14'h1423 == index ? 14'h85 : _GEN_5154;
  wire [13:0] _GEN_5156 = 14'h1424 == index ? 14'h84 : _GEN_5155;
  wire [13:0] _GEN_5157 = 14'h1425 == index ? 14'h83 : _GEN_5156;
  wire [13:0] _GEN_5158 = 14'h1426 == index ? 14'h82 : _GEN_5157;
  wire [13:0] _GEN_5159 = 14'h1427 == index ? 14'h81 : _GEN_5158;
  wire [13:0] _GEN_5160 = 14'h1428 == index ? 14'h80 : _GEN_5159;
  wire [13:0] _GEN_5161 = 14'h1429 == index ? 14'h28 : _GEN_5160;
  wire [13:0] _GEN_5162 = 14'h142a == index ? 14'h28 : _GEN_5161;
  wire [13:0] _GEN_5163 = 14'h142b == index ? 14'h28 : _GEN_5162;
  wire [13:0] _GEN_5164 = 14'h142c == index ? 14'h28 : _GEN_5163;
  wire [13:0] _GEN_5165 = 14'h142d == index ? 14'h28 : _GEN_5164;
  wire [13:0] _GEN_5166 = 14'h142e == index ? 14'h28 : _GEN_5165;
  wire [13:0] _GEN_5167 = 14'h142f == index ? 14'h28 : _GEN_5166;
  wire [13:0] _GEN_5168 = 14'h1430 == index ? 14'h28 : _GEN_5167;
  wire [13:0] _GEN_5169 = 14'h1431 == index ? 14'h28 : _GEN_5168;
  wire [13:0] _GEN_5170 = 14'h1432 == index ? 14'h28 : _GEN_5169;
  wire [13:0] _GEN_5171 = 14'h1433 == index ? 14'h28 : _GEN_5170;
  wire [13:0] _GEN_5172 = 14'h1434 == index ? 14'h28 : _GEN_5171;
  wire [13:0] _GEN_5173 = 14'h1435 == index ? 14'h28 : _GEN_5172;
  wire [13:0] _GEN_5174 = 14'h1436 == index ? 14'h28 : _GEN_5173;
  wire [13:0] _GEN_5175 = 14'h1437 == index ? 14'h28 : _GEN_5174;
  wire [13:0] _GEN_5176 = 14'h1438 == index ? 14'h28 : _GEN_5175;
  wire [13:0] _GEN_5177 = 14'h1439 == index ? 14'h28 : _GEN_5176;
  wire [13:0] _GEN_5178 = 14'h143a == index ? 14'h28 : _GEN_5177;
  wire [13:0] _GEN_5179 = 14'h143b == index ? 14'h28 : _GEN_5178;
  wire [13:0] _GEN_5180 = 14'h143c == index ? 14'h28 : _GEN_5179;
  wire [13:0] _GEN_5181 = 14'h143d == index ? 14'h28 : _GEN_5180;
  wire [13:0] _GEN_5182 = 14'h143e == index ? 14'h28 : _GEN_5181;
  wire [13:0] _GEN_5183 = 14'h143f == index ? 14'h28 : _GEN_5182;
  wire [13:0] _GEN_5184 = 14'h1440 == index ? 14'h28 : _GEN_5183;
  wire [13:0] _GEN_5185 = 14'h1441 == index ? 14'h28 : _GEN_5184;
  wire [13:0] _GEN_5186 = 14'h1442 == index ? 14'h28 : _GEN_5185;
  wire [13:0] _GEN_5187 = 14'h1443 == index ? 14'h28 : _GEN_5186;
  wire [13:0] _GEN_5188 = 14'h1444 == index ? 14'h28 : _GEN_5187;
  wire [13:0] _GEN_5189 = 14'h1445 == index ? 14'h28 : _GEN_5188;
  wire [13:0] _GEN_5190 = 14'h1446 == index ? 14'h28 : _GEN_5189;
  wire [13:0] _GEN_5191 = 14'h1447 == index ? 14'h28 : _GEN_5190;
  wire [13:0] _GEN_5192 = 14'h1448 == index ? 14'h28 : _GEN_5191;
  wire [13:0] _GEN_5193 = 14'h1449 == index ? 14'h28 : _GEN_5192;
  wire [13:0] _GEN_5194 = 14'h144a == index ? 14'h28 : _GEN_5193;
  wire [13:0] _GEN_5195 = 14'h144b == index ? 14'h28 : _GEN_5194;
  wire [13:0] _GEN_5196 = 14'h144c == index ? 14'h28 : _GEN_5195;
  wire [13:0] _GEN_5197 = 14'h144d == index ? 14'h28 : _GEN_5196;
  wire [13:0] _GEN_5198 = 14'h144e == index ? 14'h28 : _GEN_5197;
  wire [13:0] _GEN_5199 = 14'h144f == index ? 14'h28 : _GEN_5198;
  wire [13:0] _GEN_5200 = 14'h1450 == index ? 14'h28 : _GEN_5199;
  wire [13:0] _GEN_5201 = 14'h1451 == index ? 14'h28 : _GEN_5200;
  wire [13:0] _GEN_5202 = 14'h1452 == index ? 14'h28 : _GEN_5201;
  wire [13:0] _GEN_5203 = 14'h1453 == index ? 14'h28 : _GEN_5202;
  wire [13:0] _GEN_5204 = 14'h1454 == index ? 14'h28 : _GEN_5203;
  wire [13:0] _GEN_5205 = 14'h1455 == index ? 14'h28 : _GEN_5204;
  wire [13:0] _GEN_5206 = 14'h1456 == index ? 14'h28 : _GEN_5205;
  wire [13:0] _GEN_5207 = 14'h1457 == index ? 14'h28 : _GEN_5206;
  wire [13:0] _GEN_5208 = 14'h1458 == index ? 14'h28 : _GEN_5207;
  wire [13:0] _GEN_5209 = 14'h1459 == index ? 14'h28 : _GEN_5208;
  wire [13:0] _GEN_5210 = 14'h145a == index ? 14'h28 : _GEN_5209;
  wire [13:0] _GEN_5211 = 14'h145b == index ? 14'h28 : _GEN_5210;
  wire [13:0] _GEN_5212 = 14'h145c == index ? 14'h28 : _GEN_5211;
  wire [13:0] _GEN_5213 = 14'h145d == index ? 14'h28 : _GEN_5212;
  wire [13:0] _GEN_5214 = 14'h145e == index ? 14'h28 : _GEN_5213;
  wire [13:0] _GEN_5215 = 14'h145f == index ? 14'h28 : _GEN_5214;
  wire [13:0] _GEN_5216 = 14'h1460 == index ? 14'h28 : _GEN_5215;
  wire [13:0] _GEN_5217 = 14'h1461 == index ? 14'h28 : _GEN_5216;
  wire [13:0] _GEN_5218 = 14'h1462 == index ? 14'h28 : _GEN_5217;
  wire [13:0] _GEN_5219 = 14'h1463 == index ? 14'h28 : _GEN_5218;
  wire [13:0] _GEN_5220 = 14'h1464 == index ? 14'h28 : _GEN_5219;
  wire [13:0] _GEN_5221 = 14'h1465 == index ? 14'h28 : _GEN_5220;
  wire [13:0] _GEN_5222 = 14'h1466 == index ? 14'h28 : _GEN_5221;
  wire [13:0] _GEN_5223 = 14'h1467 == index ? 14'h28 : _GEN_5222;
  wire [13:0] _GEN_5224 = 14'h1468 == index ? 14'h28 : _GEN_5223;
  wire [13:0] _GEN_5225 = 14'h1469 == index ? 14'h28 : _GEN_5224;
  wire [13:0] _GEN_5226 = 14'h146a == index ? 14'h28 : _GEN_5225;
  wire [13:0] _GEN_5227 = 14'h146b == index ? 14'h28 : _GEN_5226;
  wire [13:0] _GEN_5228 = 14'h146c == index ? 14'h28 : _GEN_5227;
  wire [13:0] _GEN_5229 = 14'h146d == index ? 14'h28 : _GEN_5228;
  wire [13:0] _GEN_5230 = 14'h146e == index ? 14'h28 : _GEN_5229;
  wire [13:0] _GEN_5231 = 14'h146f == index ? 14'h28 : _GEN_5230;
  wire [13:0] _GEN_5232 = 14'h1470 == index ? 14'h28 : _GEN_5231;
  wire [13:0] _GEN_5233 = 14'h1471 == index ? 14'h28 : _GEN_5232;
  wire [13:0] _GEN_5234 = 14'h1472 == index ? 14'h28 : _GEN_5233;
  wire [13:0] _GEN_5235 = 14'h1473 == index ? 14'h28 : _GEN_5234;
  wire [13:0] _GEN_5236 = 14'h1474 == index ? 14'h28 : _GEN_5235;
  wire [13:0] _GEN_5237 = 14'h1475 == index ? 14'h28 : _GEN_5236;
  wire [13:0] _GEN_5238 = 14'h1476 == index ? 14'h28 : _GEN_5237;
  wire [13:0] _GEN_5239 = 14'h1477 == index ? 14'h28 : _GEN_5238;
  wire [13:0] _GEN_5240 = 14'h1478 == index ? 14'h28 : _GEN_5239;
  wire [13:0] _GEN_5241 = 14'h1479 == index ? 14'h28 : _GEN_5240;
  wire [13:0] _GEN_5242 = 14'h147a == index ? 14'h28 : _GEN_5241;
  wire [13:0] _GEN_5243 = 14'h147b == index ? 14'h28 : _GEN_5242;
  wire [13:0] _GEN_5244 = 14'h147c == index ? 14'h28 : _GEN_5243;
  wire [13:0] _GEN_5245 = 14'h147d == index ? 14'h28 : _GEN_5244;
  wire [13:0] _GEN_5246 = 14'h147e == index ? 14'h28 : _GEN_5245;
  wire [13:0] _GEN_5247 = 14'h147f == index ? 14'h28 : _GEN_5246;
  wire [13:0] _GEN_5248 = 14'h1480 == index ? 14'h0 : _GEN_5247;
  wire [13:0] _GEN_5249 = 14'h1481 == index ? 14'h1480 : _GEN_5248;
  wire [13:0] _GEN_5250 = 14'h1482 == index ? 14'ha01 : _GEN_5249;
  wire [13:0] _GEN_5251 = 14'h1483 == index ? 14'h682 : _GEN_5250;
  wire [13:0] _GEN_5252 = 14'h1484 == index ? 14'h501 : _GEN_5251;
  wire [13:0] _GEN_5253 = 14'h1485 == index ? 14'h401 : _GEN_5252;
  wire [13:0] _GEN_5254 = 14'h1486 == index ? 14'h305 : _GEN_5253;
  wire [13:0] _GEN_5255 = 14'h1487 == index ? 14'h286 : _GEN_5254;
  wire [13:0] _GEN_5256 = 14'h1488 == index ? 14'h281 : _GEN_5255;
  wire [13:0] _GEN_5257 = 14'h1489 == index ? 14'h205 : _GEN_5256;
  wire [13:0] _GEN_5258 = 14'h148a == index ? 14'h201 : _GEN_5257;
  wire [13:0] _GEN_5259 = 14'h148b == index ? 14'h188 : _GEN_5258;
  wire [13:0] _GEN_5260 = 14'h148c == index ? 14'h185 : _GEN_5259;
  wire [13:0] _GEN_5261 = 14'h148d == index ? 14'h182 : _GEN_5260;
  wire [13:0] _GEN_5262 = 14'h148e == index ? 14'h10d : _GEN_5261;
  wire [13:0] _GEN_5263 = 14'h148f == index ? 14'h10b : _GEN_5262;
  wire [13:0] _GEN_5264 = 14'h1490 == index ? 14'h109 : _GEN_5263;
  wire [13:0] _GEN_5265 = 14'h1491 == index ? 14'h107 : _GEN_5264;
  wire [13:0] _GEN_5266 = 14'h1492 == index ? 14'h105 : _GEN_5265;
  wire [13:0] _GEN_5267 = 14'h1493 == index ? 14'h103 : _GEN_5266;
  wire [13:0] _GEN_5268 = 14'h1494 == index ? 14'h101 : _GEN_5267;
  wire [13:0] _GEN_5269 = 14'h1495 == index ? 14'h94 : _GEN_5268;
  wire [13:0] _GEN_5270 = 14'h1496 == index ? 14'h93 : _GEN_5269;
  wire [13:0] _GEN_5271 = 14'h1497 == index ? 14'h92 : _GEN_5270;
  wire [13:0] _GEN_5272 = 14'h1498 == index ? 14'h91 : _GEN_5271;
  wire [13:0] _GEN_5273 = 14'h1499 == index ? 14'h90 : _GEN_5272;
  wire [13:0] _GEN_5274 = 14'h149a == index ? 14'h8f : _GEN_5273;
  wire [13:0] _GEN_5275 = 14'h149b == index ? 14'h8e : _GEN_5274;
  wire [13:0] _GEN_5276 = 14'h149c == index ? 14'h8d : _GEN_5275;
  wire [13:0] _GEN_5277 = 14'h149d == index ? 14'h8c : _GEN_5276;
  wire [13:0] _GEN_5278 = 14'h149e == index ? 14'h8b : _GEN_5277;
  wire [13:0] _GEN_5279 = 14'h149f == index ? 14'h8a : _GEN_5278;
  wire [13:0] _GEN_5280 = 14'h14a0 == index ? 14'h89 : _GEN_5279;
  wire [13:0] _GEN_5281 = 14'h14a1 == index ? 14'h88 : _GEN_5280;
  wire [13:0] _GEN_5282 = 14'h14a2 == index ? 14'h87 : _GEN_5281;
  wire [13:0] _GEN_5283 = 14'h14a3 == index ? 14'h86 : _GEN_5282;
  wire [13:0] _GEN_5284 = 14'h14a4 == index ? 14'h85 : _GEN_5283;
  wire [13:0] _GEN_5285 = 14'h14a5 == index ? 14'h84 : _GEN_5284;
  wire [13:0] _GEN_5286 = 14'h14a6 == index ? 14'h83 : _GEN_5285;
  wire [13:0] _GEN_5287 = 14'h14a7 == index ? 14'h82 : _GEN_5286;
  wire [13:0] _GEN_5288 = 14'h14a8 == index ? 14'h81 : _GEN_5287;
  wire [13:0] _GEN_5289 = 14'h14a9 == index ? 14'h80 : _GEN_5288;
  wire [13:0] _GEN_5290 = 14'h14aa == index ? 14'h29 : _GEN_5289;
  wire [13:0] _GEN_5291 = 14'h14ab == index ? 14'h29 : _GEN_5290;
  wire [13:0] _GEN_5292 = 14'h14ac == index ? 14'h29 : _GEN_5291;
  wire [13:0] _GEN_5293 = 14'h14ad == index ? 14'h29 : _GEN_5292;
  wire [13:0] _GEN_5294 = 14'h14ae == index ? 14'h29 : _GEN_5293;
  wire [13:0] _GEN_5295 = 14'h14af == index ? 14'h29 : _GEN_5294;
  wire [13:0] _GEN_5296 = 14'h14b0 == index ? 14'h29 : _GEN_5295;
  wire [13:0] _GEN_5297 = 14'h14b1 == index ? 14'h29 : _GEN_5296;
  wire [13:0] _GEN_5298 = 14'h14b2 == index ? 14'h29 : _GEN_5297;
  wire [13:0] _GEN_5299 = 14'h14b3 == index ? 14'h29 : _GEN_5298;
  wire [13:0] _GEN_5300 = 14'h14b4 == index ? 14'h29 : _GEN_5299;
  wire [13:0] _GEN_5301 = 14'h14b5 == index ? 14'h29 : _GEN_5300;
  wire [13:0] _GEN_5302 = 14'h14b6 == index ? 14'h29 : _GEN_5301;
  wire [13:0] _GEN_5303 = 14'h14b7 == index ? 14'h29 : _GEN_5302;
  wire [13:0] _GEN_5304 = 14'h14b8 == index ? 14'h29 : _GEN_5303;
  wire [13:0] _GEN_5305 = 14'h14b9 == index ? 14'h29 : _GEN_5304;
  wire [13:0] _GEN_5306 = 14'h14ba == index ? 14'h29 : _GEN_5305;
  wire [13:0] _GEN_5307 = 14'h14bb == index ? 14'h29 : _GEN_5306;
  wire [13:0] _GEN_5308 = 14'h14bc == index ? 14'h29 : _GEN_5307;
  wire [13:0] _GEN_5309 = 14'h14bd == index ? 14'h29 : _GEN_5308;
  wire [13:0] _GEN_5310 = 14'h14be == index ? 14'h29 : _GEN_5309;
  wire [13:0] _GEN_5311 = 14'h14bf == index ? 14'h29 : _GEN_5310;
  wire [13:0] _GEN_5312 = 14'h14c0 == index ? 14'h29 : _GEN_5311;
  wire [13:0] _GEN_5313 = 14'h14c1 == index ? 14'h29 : _GEN_5312;
  wire [13:0] _GEN_5314 = 14'h14c2 == index ? 14'h29 : _GEN_5313;
  wire [13:0] _GEN_5315 = 14'h14c3 == index ? 14'h29 : _GEN_5314;
  wire [13:0] _GEN_5316 = 14'h14c4 == index ? 14'h29 : _GEN_5315;
  wire [13:0] _GEN_5317 = 14'h14c5 == index ? 14'h29 : _GEN_5316;
  wire [13:0] _GEN_5318 = 14'h14c6 == index ? 14'h29 : _GEN_5317;
  wire [13:0] _GEN_5319 = 14'h14c7 == index ? 14'h29 : _GEN_5318;
  wire [13:0] _GEN_5320 = 14'h14c8 == index ? 14'h29 : _GEN_5319;
  wire [13:0] _GEN_5321 = 14'h14c9 == index ? 14'h29 : _GEN_5320;
  wire [13:0] _GEN_5322 = 14'h14ca == index ? 14'h29 : _GEN_5321;
  wire [13:0] _GEN_5323 = 14'h14cb == index ? 14'h29 : _GEN_5322;
  wire [13:0] _GEN_5324 = 14'h14cc == index ? 14'h29 : _GEN_5323;
  wire [13:0] _GEN_5325 = 14'h14cd == index ? 14'h29 : _GEN_5324;
  wire [13:0] _GEN_5326 = 14'h14ce == index ? 14'h29 : _GEN_5325;
  wire [13:0] _GEN_5327 = 14'h14cf == index ? 14'h29 : _GEN_5326;
  wire [13:0] _GEN_5328 = 14'h14d0 == index ? 14'h29 : _GEN_5327;
  wire [13:0] _GEN_5329 = 14'h14d1 == index ? 14'h29 : _GEN_5328;
  wire [13:0] _GEN_5330 = 14'h14d2 == index ? 14'h29 : _GEN_5329;
  wire [13:0] _GEN_5331 = 14'h14d3 == index ? 14'h29 : _GEN_5330;
  wire [13:0] _GEN_5332 = 14'h14d4 == index ? 14'h29 : _GEN_5331;
  wire [13:0] _GEN_5333 = 14'h14d5 == index ? 14'h29 : _GEN_5332;
  wire [13:0] _GEN_5334 = 14'h14d6 == index ? 14'h29 : _GEN_5333;
  wire [13:0] _GEN_5335 = 14'h14d7 == index ? 14'h29 : _GEN_5334;
  wire [13:0] _GEN_5336 = 14'h14d8 == index ? 14'h29 : _GEN_5335;
  wire [13:0] _GEN_5337 = 14'h14d9 == index ? 14'h29 : _GEN_5336;
  wire [13:0] _GEN_5338 = 14'h14da == index ? 14'h29 : _GEN_5337;
  wire [13:0] _GEN_5339 = 14'h14db == index ? 14'h29 : _GEN_5338;
  wire [13:0] _GEN_5340 = 14'h14dc == index ? 14'h29 : _GEN_5339;
  wire [13:0] _GEN_5341 = 14'h14dd == index ? 14'h29 : _GEN_5340;
  wire [13:0] _GEN_5342 = 14'h14de == index ? 14'h29 : _GEN_5341;
  wire [13:0] _GEN_5343 = 14'h14df == index ? 14'h29 : _GEN_5342;
  wire [13:0] _GEN_5344 = 14'h14e0 == index ? 14'h29 : _GEN_5343;
  wire [13:0] _GEN_5345 = 14'h14e1 == index ? 14'h29 : _GEN_5344;
  wire [13:0] _GEN_5346 = 14'h14e2 == index ? 14'h29 : _GEN_5345;
  wire [13:0] _GEN_5347 = 14'h14e3 == index ? 14'h29 : _GEN_5346;
  wire [13:0] _GEN_5348 = 14'h14e4 == index ? 14'h29 : _GEN_5347;
  wire [13:0] _GEN_5349 = 14'h14e5 == index ? 14'h29 : _GEN_5348;
  wire [13:0] _GEN_5350 = 14'h14e6 == index ? 14'h29 : _GEN_5349;
  wire [13:0] _GEN_5351 = 14'h14e7 == index ? 14'h29 : _GEN_5350;
  wire [13:0] _GEN_5352 = 14'h14e8 == index ? 14'h29 : _GEN_5351;
  wire [13:0] _GEN_5353 = 14'h14e9 == index ? 14'h29 : _GEN_5352;
  wire [13:0] _GEN_5354 = 14'h14ea == index ? 14'h29 : _GEN_5353;
  wire [13:0] _GEN_5355 = 14'h14eb == index ? 14'h29 : _GEN_5354;
  wire [13:0] _GEN_5356 = 14'h14ec == index ? 14'h29 : _GEN_5355;
  wire [13:0] _GEN_5357 = 14'h14ed == index ? 14'h29 : _GEN_5356;
  wire [13:0] _GEN_5358 = 14'h14ee == index ? 14'h29 : _GEN_5357;
  wire [13:0] _GEN_5359 = 14'h14ef == index ? 14'h29 : _GEN_5358;
  wire [13:0] _GEN_5360 = 14'h14f0 == index ? 14'h29 : _GEN_5359;
  wire [13:0] _GEN_5361 = 14'h14f1 == index ? 14'h29 : _GEN_5360;
  wire [13:0] _GEN_5362 = 14'h14f2 == index ? 14'h29 : _GEN_5361;
  wire [13:0] _GEN_5363 = 14'h14f3 == index ? 14'h29 : _GEN_5362;
  wire [13:0] _GEN_5364 = 14'h14f4 == index ? 14'h29 : _GEN_5363;
  wire [13:0] _GEN_5365 = 14'h14f5 == index ? 14'h29 : _GEN_5364;
  wire [13:0] _GEN_5366 = 14'h14f6 == index ? 14'h29 : _GEN_5365;
  wire [13:0] _GEN_5367 = 14'h14f7 == index ? 14'h29 : _GEN_5366;
  wire [13:0] _GEN_5368 = 14'h14f8 == index ? 14'h29 : _GEN_5367;
  wire [13:0] _GEN_5369 = 14'h14f9 == index ? 14'h29 : _GEN_5368;
  wire [13:0] _GEN_5370 = 14'h14fa == index ? 14'h29 : _GEN_5369;
  wire [13:0] _GEN_5371 = 14'h14fb == index ? 14'h29 : _GEN_5370;
  wire [13:0] _GEN_5372 = 14'h14fc == index ? 14'h29 : _GEN_5371;
  wire [13:0] _GEN_5373 = 14'h14fd == index ? 14'h29 : _GEN_5372;
  wire [13:0] _GEN_5374 = 14'h14fe == index ? 14'h29 : _GEN_5373;
  wire [13:0] _GEN_5375 = 14'h14ff == index ? 14'h29 : _GEN_5374;
  wire [13:0] _GEN_5376 = 14'h1500 == index ? 14'h0 : _GEN_5375;
  wire [13:0] _GEN_5377 = 14'h1501 == index ? 14'h1500 : _GEN_5376;
  wire [13:0] _GEN_5378 = 14'h1502 == index ? 14'ha80 : _GEN_5377;
  wire [13:0] _GEN_5379 = 14'h1503 == index ? 14'h700 : _GEN_5378;
  wire [13:0] _GEN_5380 = 14'h1504 == index ? 14'h502 : _GEN_5379;
  wire [13:0] _GEN_5381 = 14'h1505 == index ? 14'h402 : _GEN_5380;
  wire [13:0] _GEN_5382 = 14'h1506 == index ? 14'h380 : _GEN_5381;
  wire [13:0] _GEN_5383 = 14'h1507 == index ? 14'h300 : _GEN_5382;
  wire [13:0] _GEN_5384 = 14'h1508 == index ? 14'h282 : _GEN_5383;
  wire [13:0] _GEN_5385 = 14'h1509 == index ? 14'h206 : _GEN_5384;
  wire [13:0] _GEN_5386 = 14'h150a == index ? 14'h202 : _GEN_5385;
  wire [13:0] _GEN_5387 = 14'h150b == index ? 14'h189 : _GEN_5386;
  wire [13:0] _GEN_5388 = 14'h150c == index ? 14'h186 : _GEN_5387;
  wire [13:0] _GEN_5389 = 14'h150d == index ? 14'h183 : _GEN_5388;
  wire [13:0] _GEN_5390 = 14'h150e == index ? 14'h180 : _GEN_5389;
  wire [13:0] _GEN_5391 = 14'h150f == index ? 14'h10c : _GEN_5390;
  wire [13:0] _GEN_5392 = 14'h1510 == index ? 14'h10a : _GEN_5391;
  wire [13:0] _GEN_5393 = 14'h1511 == index ? 14'h108 : _GEN_5392;
  wire [13:0] _GEN_5394 = 14'h1512 == index ? 14'h106 : _GEN_5393;
  wire [13:0] _GEN_5395 = 14'h1513 == index ? 14'h104 : _GEN_5394;
  wire [13:0] _GEN_5396 = 14'h1514 == index ? 14'h102 : _GEN_5395;
  wire [13:0] _GEN_5397 = 14'h1515 == index ? 14'h100 : _GEN_5396;
  wire [13:0] _GEN_5398 = 14'h1516 == index ? 14'h94 : _GEN_5397;
  wire [13:0] _GEN_5399 = 14'h1517 == index ? 14'h93 : _GEN_5398;
  wire [13:0] _GEN_5400 = 14'h1518 == index ? 14'h92 : _GEN_5399;
  wire [13:0] _GEN_5401 = 14'h1519 == index ? 14'h91 : _GEN_5400;
  wire [13:0] _GEN_5402 = 14'h151a == index ? 14'h90 : _GEN_5401;
  wire [13:0] _GEN_5403 = 14'h151b == index ? 14'h8f : _GEN_5402;
  wire [13:0] _GEN_5404 = 14'h151c == index ? 14'h8e : _GEN_5403;
  wire [13:0] _GEN_5405 = 14'h151d == index ? 14'h8d : _GEN_5404;
  wire [13:0] _GEN_5406 = 14'h151e == index ? 14'h8c : _GEN_5405;
  wire [13:0] _GEN_5407 = 14'h151f == index ? 14'h8b : _GEN_5406;
  wire [13:0] _GEN_5408 = 14'h1520 == index ? 14'h8a : _GEN_5407;
  wire [13:0] _GEN_5409 = 14'h1521 == index ? 14'h89 : _GEN_5408;
  wire [13:0] _GEN_5410 = 14'h1522 == index ? 14'h88 : _GEN_5409;
  wire [13:0] _GEN_5411 = 14'h1523 == index ? 14'h87 : _GEN_5410;
  wire [13:0] _GEN_5412 = 14'h1524 == index ? 14'h86 : _GEN_5411;
  wire [13:0] _GEN_5413 = 14'h1525 == index ? 14'h85 : _GEN_5412;
  wire [13:0] _GEN_5414 = 14'h1526 == index ? 14'h84 : _GEN_5413;
  wire [13:0] _GEN_5415 = 14'h1527 == index ? 14'h83 : _GEN_5414;
  wire [13:0] _GEN_5416 = 14'h1528 == index ? 14'h82 : _GEN_5415;
  wire [13:0] _GEN_5417 = 14'h1529 == index ? 14'h81 : _GEN_5416;
  wire [13:0] _GEN_5418 = 14'h152a == index ? 14'h80 : _GEN_5417;
  wire [13:0] _GEN_5419 = 14'h152b == index ? 14'h2a : _GEN_5418;
  wire [13:0] _GEN_5420 = 14'h152c == index ? 14'h2a : _GEN_5419;
  wire [13:0] _GEN_5421 = 14'h152d == index ? 14'h2a : _GEN_5420;
  wire [13:0] _GEN_5422 = 14'h152e == index ? 14'h2a : _GEN_5421;
  wire [13:0] _GEN_5423 = 14'h152f == index ? 14'h2a : _GEN_5422;
  wire [13:0] _GEN_5424 = 14'h1530 == index ? 14'h2a : _GEN_5423;
  wire [13:0] _GEN_5425 = 14'h1531 == index ? 14'h2a : _GEN_5424;
  wire [13:0] _GEN_5426 = 14'h1532 == index ? 14'h2a : _GEN_5425;
  wire [13:0] _GEN_5427 = 14'h1533 == index ? 14'h2a : _GEN_5426;
  wire [13:0] _GEN_5428 = 14'h1534 == index ? 14'h2a : _GEN_5427;
  wire [13:0] _GEN_5429 = 14'h1535 == index ? 14'h2a : _GEN_5428;
  wire [13:0] _GEN_5430 = 14'h1536 == index ? 14'h2a : _GEN_5429;
  wire [13:0] _GEN_5431 = 14'h1537 == index ? 14'h2a : _GEN_5430;
  wire [13:0] _GEN_5432 = 14'h1538 == index ? 14'h2a : _GEN_5431;
  wire [13:0] _GEN_5433 = 14'h1539 == index ? 14'h2a : _GEN_5432;
  wire [13:0] _GEN_5434 = 14'h153a == index ? 14'h2a : _GEN_5433;
  wire [13:0] _GEN_5435 = 14'h153b == index ? 14'h2a : _GEN_5434;
  wire [13:0] _GEN_5436 = 14'h153c == index ? 14'h2a : _GEN_5435;
  wire [13:0] _GEN_5437 = 14'h153d == index ? 14'h2a : _GEN_5436;
  wire [13:0] _GEN_5438 = 14'h153e == index ? 14'h2a : _GEN_5437;
  wire [13:0] _GEN_5439 = 14'h153f == index ? 14'h2a : _GEN_5438;
  wire [13:0] _GEN_5440 = 14'h1540 == index ? 14'h2a : _GEN_5439;
  wire [13:0] _GEN_5441 = 14'h1541 == index ? 14'h2a : _GEN_5440;
  wire [13:0] _GEN_5442 = 14'h1542 == index ? 14'h2a : _GEN_5441;
  wire [13:0] _GEN_5443 = 14'h1543 == index ? 14'h2a : _GEN_5442;
  wire [13:0] _GEN_5444 = 14'h1544 == index ? 14'h2a : _GEN_5443;
  wire [13:0] _GEN_5445 = 14'h1545 == index ? 14'h2a : _GEN_5444;
  wire [13:0] _GEN_5446 = 14'h1546 == index ? 14'h2a : _GEN_5445;
  wire [13:0] _GEN_5447 = 14'h1547 == index ? 14'h2a : _GEN_5446;
  wire [13:0] _GEN_5448 = 14'h1548 == index ? 14'h2a : _GEN_5447;
  wire [13:0] _GEN_5449 = 14'h1549 == index ? 14'h2a : _GEN_5448;
  wire [13:0] _GEN_5450 = 14'h154a == index ? 14'h2a : _GEN_5449;
  wire [13:0] _GEN_5451 = 14'h154b == index ? 14'h2a : _GEN_5450;
  wire [13:0] _GEN_5452 = 14'h154c == index ? 14'h2a : _GEN_5451;
  wire [13:0] _GEN_5453 = 14'h154d == index ? 14'h2a : _GEN_5452;
  wire [13:0] _GEN_5454 = 14'h154e == index ? 14'h2a : _GEN_5453;
  wire [13:0] _GEN_5455 = 14'h154f == index ? 14'h2a : _GEN_5454;
  wire [13:0] _GEN_5456 = 14'h1550 == index ? 14'h2a : _GEN_5455;
  wire [13:0] _GEN_5457 = 14'h1551 == index ? 14'h2a : _GEN_5456;
  wire [13:0] _GEN_5458 = 14'h1552 == index ? 14'h2a : _GEN_5457;
  wire [13:0] _GEN_5459 = 14'h1553 == index ? 14'h2a : _GEN_5458;
  wire [13:0] _GEN_5460 = 14'h1554 == index ? 14'h2a : _GEN_5459;
  wire [13:0] _GEN_5461 = 14'h1555 == index ? 14'h2a : _GEN_5460;
  wire [13:0] _GEN_5462 = 14'h1556 == index ? 14'h2a : _GEN_5461;
  wire [13:0] _GEN_5463 = 14'h1557 == index ? 14'h2a : _GEN_5462;
  wire [13:0] _GEN_5464 = 14'h1558 == index ? 14'h2a : _GEN_5463;
  wire [13:0] _GEN_5465 = 14'h1559 == index ? 14'h2a : _GEN_5464;
  wire [13:0] _GEN_5466 = 14'h155a == index ? 14'h2a : _GEN_5465;
  wire [13:0] _GEN_5467 = 14'h155b == index ? 14'h2a : _GEN_5466;
  wire [13:0] _GEN_5468 = 14'h155c == index ? 14'h2a : _GEN_5467;
  wire [13:0] _GEN_5469 = 14'h155d == index ? 14'h2a : _GEN_5468;
  wire [13:0] _GEN_5470 = 14'h155e == index ? 14'h2a : _GEN_5469;
  wire [13:0] _GEN_5471 = 14'h155f == index ? 14'h2a : _GEN_5470;
  wire [13:0] _GEN_5472 = 14'h1560 == index ? 14'h2a : _GEN_5471;
  wire [13:0] _GEN_5473 = 14'h1561 == index ? 14'h2a : _GEN_5472;
  wire [13:0] _GEN_5474 = 14'h1562 == index ? 14'h2a : _GEN_5473;
  wire [13:0] _GEN_5475 = 14'h1563 == index ? 14'h2a : _GEN_5474;
  wire [13:0] _GEN_5476 = 14'h1564 == index ? 14'h2a : _GEN_5475;
  wire [13:0] _GEN_5477 = 14'h1565 == index ? 14'h2a : _GEN_5476;
  wire [13:0] _GEN_5478 = 14'h1566 == index ? 14'h2a : _GEN_5477;
  wire [13:0] _GEN_5479 = 14'h1567 == index ? 14'h2a : _GEN_5478;
  wire [13:0] _GEN_5480 = 14'h1568 == index ? 14'h2a : _GEN_5479;
  wire [13:0] _GEN_5481 = 14'h1569 == index ? 14'h2a : _GEN_5480;
  wire [13:0] _GEN_5482 = 14'h156a == index ? 14'h2a : _GEN_5481;
  wire [13:0] _GEN_5483 = 14'h156b == index ? 14'h2a : _GEN_5482;
  wire [13:0] _GEN_5484 = 14'h156c == index ? 14'h2a : _GEN_5483;
  wire [13:0] _GEN_5485 = 14'h156d == index ? 14'h2a : _GEN_5484;
  wire [13:0] _GEN_5486 = 14'h156e == index ? 14'h2a : _GEN_5485;
  wire [13:0] _GEN_5487 = 14'h156f == index ? 14'h2a : _GEN_5486;
  wire [13:0] _GEN_5488 = 14'h1570 == index ? 14'h2a : _GEN_5487;
  wire [13:0] _GEN_5489 = 14'h1571 == index ? 14'h2a : _GEN_5488;
  wire [13:0] _GEN_5490 = 14'h1572 == index ? 14'h2a : _GEN_5489;
  wire [13:0] _GEN_5491 = 14'h1573 == index ? 14'h2a : _GEN_5490;
  wire [13:0] _GEN_5492 = 14'h1574 == index ? 14'h2a : _GEN_5491;
  wire [13:0] _GEN_5493 = 14'h1575 == index ? 14'h2a : _GEN_5492;
  wire [13:0] _GEN_5494 = 14'h1576 == index ? 14'h2a : _GEN_5493;
  wire [13:0] _GEN_5495 = 14'h1577 == index ? 14'h2a : _GEN_5494;
  wire [13:0] _GEN_5496 = 14'h1578 == index ? 14'h2a : _GEN_5495;
  wire [13:0] _GEN_5497 = 14'h1579 == index ? 14'h2a : _GEN_5496;
  wire [13:0] _GEN_5498 = 14'h157a == index ? 14'h2a : _GEN_5497;
  wire [13:0] _GEN_5499 = 14'h157b == index ? 14'h2a : _GEN_5498;
  wire [13:0] _GEN_5500 = 14'h157c == index ? 14'h2a : _GEN_5499;
  wire [13:0] _GEN_5501 = 14'h157d == index ? 14'h2a : _GEN_5500;
  wire [13:0] _GEN_5502 = 14'h157e == index ? 14'h2a : _GEN_5501;
  wire [13:0] _GEN_5503 = 14'h157f == index ? 14'h2a : _GEN_5502;
  wire [13:0] _GEN_5504 = 14'h1580 == index ? 14'h0 : _GEN_5503;
  wire [13:0] _GEN_5505 = 14'h1581 == index ? 14'h1580 : _GEN_5504;
  wire [13:0] _GEN_5506 = 14'h1582 == index ? 14'ha81 : _GEN_5505;
  wire [13:0] _GEN_5507 = 14'h1583 == index ? 14'h701 : _GEN_5506;
  wire [13:0] _GEN_5508 = 14'h1584 == index ? 14'h503 : _GEN_5507;
  wire [13:0] _GEN_5509 = 14'h1585 == index ? 14'h403 : _GEN_5508;
  wire [13:0] _GEN_5510 = 14'h1586 == index ? 14'h381 : _GEN_5509;
  wire [13:0] _GEN_5511 = 14'h1587 == index ? 14'h301 : _GEN_5510;
  wire [13:0] _GEN_5512 = 14'h1588 == index ? 14'h283 : _GEN_5511;
  wire [13:0] _GEN_5513 = 14'h1589 == index ? 14'h207 : _GEN_5512;
  wire [13:0] _GEN_5514 = 14'h158a == index ? 14'h203 : _GEN_5513;
  wire [13:0] _GEN_5515 = 14'h158b == index ? 14'h18a : _GEN_5514;
  wire [13:0] _GEN_5516 = 14'h158c == index ? 14'h187 : _GEN_5515;
  wire [13:0] _GEN_5517 = 14'h158d == index ? 14'h184 : _GEN_5516;
  wire [13:0] _GEN_5518 = 14'h158e == index ? 14'h181 : _GEN_5517;
  wire [13:0] _GEN_5519 = 14'h158f == index ? 14'h10d : _GEN_5518;
  wire [13:0] _GEN_5520 = 14'h1590 == index ? 14'h10b : _GEN_5519;
  wire [13:0] _GEN_5521 = 14'h1591 == index ? 14'h109 : _GEN_5520;
  wire [13:0] _GEN_5522 = 14'h1592 == index ? 14'h107 : _GEN_5521;
  wire [13:0] _GEN_5523 = 14'h1593 == index ? 14'h105 : _GEN_5522;
  wire [13:0] _GEN_5524 = 14'h1594 == index ? 14'h103 : _GEN_5523;
  wire [13:0] _GEN_5525 = 14'h1595 == index ? 14'h101 : _GEN_5524;
  wire [13:0] _GEN_5526 = 14'h1596 == index ? 14'h95 : _GEN_5525;
  wire [13:0] _GEN_5527 = 14'h1597 == index ? 14'h94 : _GEN_5526;
  wire [13:0] _GEN_5528 = 14'h1598 == index ? 14'h93 : _GEN_5527;
  wire [13:0] _GEN_5529 = 14'h1599 == index ? 14'h92 : _GEN_5528;
  wire [13:0] _GEN_5530 = 14'h159a == index ? 14'h91 : _GEN_5529;
  wire [13:0] _GEN_5531 = 14'h159b == index ? 14'h90 : _GEN_5530;
  wire [13:0] _GEN_5532 = 14'h159c == index ? 14'h8f : _GEN_5531;
  wire [13:0] _GEN_5533 = 14'h159d == index ? 14'h8e : _GEN_5532;
  wire [13:0] _GEN_5534 = 14'h159e == index ? 14'h8d : _GEN_5533;
  wire [13:0] _GEN_5535 = 14'h159f == index ? 14'h8c : _GEN_5534;
  wire [13:0] _GEN_5536 = 14'h15a0 == index ? 14'h8b : _GEN_5535;
  wire [13:0] _GEN_5537 = 14'h15a1 == index ? 14'h8a : _GEN_5536;
  wire [13:0] _GEN_5538 = 14'h15a2 == index ? 14'h89 : _GEN_5537;
  wire [13:0] _GEN_5539 = 14'h15a3 == index ? 14'h88 : _GEN_5538;
  wire [13:0] _GEN_5540 = 14'h15a4 == index ? 14'h87 : _GEN_5539;
  wire [13:0] _GEN_5541 = 14'h15a5 == index ? 14'h86 : _GEN_5540;
  wire [13:0] _GEN_5542 = 14'h15a6 == index ? 14'h85 : _GEN_5541;
  wire [13:0] _GEN_5543 = 14'h15a7 == index ? 14'h84 : _GEN_5542;
  wire [13:0] _GEN_5544 = 14'h15a8 == index ? 14'h83 : _GEN_5543;
  wire [13:0] _GEN_5545 = 14'h15a9 == index ? 14'h82 : _GEN_5544;
  wire [13:0] _GEN_5546 = 14'h15aa == index ? 14'h81 : _GEN_5545;
  wire [13:0] _GEN_5547 = 14'h15ab == index ? 14'h80 : _GEN_5546;
  wire [13:0] _GEN_5548 = 14'h15ac == index ? 14'h2b : _GEN_5547;
  wire [13:0] _GEN_5549 = 14'h15ad == index ? 14'h2b : _GEN_5548;
  wire [13:0] _GEN_5550 = 14'h15ae == index ? 14'h2b : _GEN_5549;
  wire [13:0] _GEN_5551 = 14'h15af == index ? 14'h2b : _GEN_5550;
  wire [13:0] _GEN_5552 = 14'h15b0 == index ? 14'h2b : _GEN_5551;
  wire [13:0] _GEN_5553 = 14'h15b1 == index ? 14'h2b : _GEN_5552;
  wire [13:0] _GEN_5554 = 14'h15b2 == index ? 14'h2b : _GEN_5553;
  wire [13:0] _GEN_5555 = 14'h15b3 == index ? 14'h2b : _GEN_5554;
  wire [13:0] _GEN_5556 = 14'h15b4 == index ? 14'h2b : _GEN_5555;
  wire [13:0] _GEN_5557 = 14'h15b5 == index ? 14'h2b : _GEN_5556;
  wire [13:0] _GEN_5558 = 14'h15b6 == index ? 14'h2b : _GEN_5557;
  wire [13:0] _GEN_5559 = 14'h15b7 == index ? 14'h2b : _GEN_5558;
  wire [13:0] _GEN_5560 = 14'h15b8 == index ? 14'h2b : _GEN_5559;
  wire [13:0] _GEN_5561 = 14'h15b9 == index ? 14'h2b : _GEN_5560;
  wire [13:0] _GEN_5562 = 14'h15ba == index ? 14'h2b : _GEN_5561;
  wire [13:0] _GEN_5563 = 14'h15bb == index ? 14'h2b : _GEN_5562;
  wire [13:0] _GEN_5564 = 14'h15bc == index ? 14'h2b : _GEN_5563;
  wire [13:0] _GEN_5565 = 14'h15bd == index ? 14'h2b : _GEN_5564;
  wire [13:0] _GEN_5566 = 14'h15be == index ? 14'h2b : _GEN_5565;
  wire [13:0] _GEN_5567 = 14'h15bf == index ? 14'h2b : _GEN_5566;
  wire [13:0] _GEN_5568 = 14'h15c0 == index ? 14'h2b : _GEN_5567;
  wire [13:0] _GEN_5569 = 14'h15c1 == index ? 14'h2b : _GEN_5568;
  wire [13:0] _GEN_5570 = 14'h15c2 == index ? 14'h2b : _GEN_5569;
  wire [13:0] _GEN_5571 = 14'h15c3 == index ? 14'h2b : _GEN_5570;
  wire [13:0] _GEN_5572 = 14'h15c4 == index ? 14'h2b : _GEN_5571;
  wire [13:0] _GEN_5573 = 14'h15c5 == index ? 14'h2b : _GEN_5572;
  wire [13:0] _GEN_5574 = 14'h15c6 == index ? 14'h2b : _GEN_5573;
  wire [13:0] _GEN_5575 = 14'h15c7 == index ? 14'h2b : _GEN_5574;
  wire [13:0] _GEN_5576 = 14'h15c8 == index ? 14'h2b : _GEN_5575;
  wire [13:0] _GEN_5577 = 14'h15c9 == index ? 14'h2b : _GEN_5576;
  wire [13:0] _GEN_5578 = 14'h15ca == index ? 14'h2b : _GEN_5577;
  wire [13:0] _GEN_5579 = 14'h15cb == index ? 14'h2b : _GEN_5578;
  wire [13:0] _GEN_5580 = 14'h15cc == index ? 14'h2b : _GEN_5579;
  wire [13:0] _GEN_5581 = 14'h15cd == index ? 14'h2b : _GEN_5580;
  wire [13:0] _GEN_5582 = 14'h15ce == index ? 14'h2b : _GEN_5581;
  wire [13:0] _GEN_5583 = 14'h15cf == index ? 14'h2b : _GEN_5582;
  wire [13:0] _GEN_5584 = 14'h15d0 == index ? 14'h2b : _GEN_5583;
  wire [13:0] _GEN_5585 = 14'h15d1 == index ? 14'h2b : _GEN_5584;
  wire [13:0] _GEN_5586 = 14'h15d2 == index ? 14'h2b : _GEN_5585;
  wire [13:0] _GEN_5587 = 14'h15d3 == index ? 14'h2b : _GEN_5586;
  wire [13:0] _GEN_5588 = 14'h15d4 == index ? 14'h2b : _GEN_5587;
  wire [13:0] _GEN_5589 = 14'h15d5 == index ? 14'h2b : _GEN_5588;
  wire [13:0] _GEN_5590 = 14'h15d6 == index ? 14'h2b : _GEN_5589;
  wire [13:0] _GEN_5591 = 14'h15d7 == index ? 14'h2b : _GEN_5590;
  wire [13:0] _GEN_5592 = 14'h15d8 == index ? 14'h2b : _GEN_5591;
  wire [13:0] _GEN_5593 = 14'h15d9 == index ? 14'h2b : _GEN_5592;
  wire [13:0] _GEN_5594 = 14'h15da == index ? 14'h2b : _GEN_5593;
  wire [13:0] _GEN_5595 = 14'h15db == index ? 14'h2b : _GEN_5594;
  wire [13:0] _GEN_5596 = 14'h15dc == index ? 14'h2b : _GEN_5595;
  wire [13:0] _GEN_5597 = 14'h15dd == index ? 14'h2b : _GEN_5596;
  wire [13:0] _GEN_5598 = 14'h15de == index ? 14'h2b : _GEN_5597;
  wire [13:0] _GEN_5599 = 14'h15df == index ? 14'h2b : _GEN_5598;
  wire [13:0] _GEN_5600 = 14'h15e0 == index ? 14'h2b : _GEN_5599;
  wire [13:0] _GEN_5601 = 14'h15e1 == index ? 14'h2b : _GEN_5600;
  wire [13:0] _GEN_5602 = 14'h15e2 == index ? 14'h2b : _GEN_5601;
  wire [13:0] _GEN_5603 = 14'h15e3 == index ? 14'h2b : _GEN_5602;
  wire [13:0] _GEN_5604 = 14'h15e4 == index ? 14'h2b : _GEN_5603;
  wire [13:0] _GEN_5605 = 14'h15e5 == index ? 14'h2b : _GEN_5604;
  wire [13:0] _GEN_5606 = 14'h15e6 == index ? 14'h2b : _GEN_5605;
  wire [13:0] _GEN_5607 = 14'h15e7 == index ? 14'h2b : _GEN_5606;
  wire [13:0] _GEN_5608 = 14'h15e8 == index ? 14'h2b : _GEN_5607;
  wire [13:0] _GEN_5609 = 14'h15e9 == index ? 14'h2b : _GEN_5608;
  wire [13:0] _GEN_5610 = 14'h15ea == index ? 14'h2b : _GEN_5609;
  wire [13:0] _GEN_5611 = 14'h15eb == index ? 14'h2b : _GEN_5610;
  wire [13:0] _GEN_5612 = 14'h15ec == index ? 14'h2b : _GEN_5611;
  wire [13:0] _GEN_5613 = 14'h15ed == index ? 14'h2b : _GEN_5612;
  wire [13:0] _GEN_5614 = 14'h15ee == index ? 14'h2b : _GEN_5613;
  wire [13:0] _GEN_5615 = 14'h15ef == index ? 14'h2b : _GEN_5614;
  wire [13:0] _GEN_5616 = 14'h15f0 == index ? 14'h2b : _GEN_5615;
  wire [13:0] _GEN_5617 = 14'h15f1 == index ? 14'h2b : _GEN_5616;
  wire [13:0] _GEN_5618 = 14'h15f2 == index ? 14'h2b : _GEN_5617;
  wire [13:0] _GEN_5619 = 14'h15f3 == index ? 14'h2b : _GEN_5618;
  wire [13:0] _GEN_5620 = 14'h15f4 == index ? 14'h2b : _GEN_5619;
  wire [13:0] _GEN_5621 = 14'h15f5 == index ? 14'h2b : _GEN_5620;
  wire [13:0] _GEN_5622 = 14'h15f6 == index ? 14'h2b : _GEN_5621;
  wire [13:0] _GEN_5623 = 14'h15f7 == index ? 14'h2b : _GEN_5622;
  wire [13:0] _GEN_5624 = 14'h15f8 == index ? 14'h2b : _GEN_5623;
  wire [13:0] _GEN_5625 = 14'h15f9 == index ? 14'h2b : _GEN_5624;
  wire [13:0] _GEN_5626 = 14'h15fa == index ? 14'h2b : _GEN_5625;
  wire [13:0] _GEN_5627 = 14'h15fb == index ? 14'h2b : _GEN_5626;
  wire [13:0] _GEN_5628 = 14'h15fc == index ? 14'h2b : _GEN_5627;
  wire [13:0] _GEN_5629 = 14'h15fd == index ? 14'h2b : _GEN_5628;
  wire [13:0] _GEN_5630 = 14'h15fe == index ? 14'h2b : _GEN_5629;
  wire [13:0] _GEN_5631 = 14'h15ff == index ? 14'h2b : _GEN_5630;
  wire [13:0] _GEN_5632 = 14'h1600 == index ? 14'h0 : _GEN_5631;
  wire [13:0] _GEN_5633 = 14'h1601 == index ? 14'h1600 : _GEN_5632;
  wire [13:0] _GEN_5634 = 14'h1602 == index ? 14'hb00 : _GEN_5633;
  wire [13:0] _GEN_5635 = 14'h1603 == index ? 14'h702 : _GEN_5634;
  wire [13:0] _GEN_5636 = 14'h1604 == index ? 14'h580 : _GEN_5635;
  wire [13:0] _GEN_5637 = 14'h1605 == index ? 14'h404 : _GEN_5636;
  wire [13:0] _GEN_5638 = 14'h1606 == index ? 14'h382 : _GEN_5637;
  wire [13:0] _GEN_5639 = 14'h1607 == index ? 14'h302 : _GEN_5638;
  wire [13:0] _GEN_5640 = 14'h1608 == index ? 14'h284 : _GEN_5639;
  wire [13:0] _GEN_5641 = 14'h1609 == index ? 14'h208 : _GEN_5640;
  wire [13:0] _GEN_5642 = 14'h160a == index ? 14'h204 : _GEN_5641;
  wire [13:0] _GEN_5643 = 14'h160b == index ? 14'h200 : _GEN_5642;
  wire [13:0] _GEN_5644 = 14'h160c == index ? 14'h188 : _GEN_5643;
  wire [13:0] _GEN_5645 = 14'h160d == index ? 14'h185 : _GEN_5644;
  wire [13:0] _GEN_5646 = 14'h160e == index ? 14'h182 : _GEN_5645;
  wire [13:0] _GEN_5647 = 14'h160f == index ? 14'h10e : _GEN_5646;
  wire [13:0] _GEN_5648 = 14'h1610 == index ? 14'h10c : _GEN_5647;
  wire [13:0] _GEN_5649 = 14'h1611 == index ? 14'h10a : _GEN_5648;
  wire [13:0] _GEN_5650 = 14'h1612 == index ? 14'h108 : _GEN_5649;
  wire [13:0] _GEN_5651 = 14'h1613 == index ? 14'h106 : _GEN_5650;
  wire [13:0] _GEN_5652 = 14'h1614 == index ? 14'h104 : _GEN_5651;
  wire [13:0] _GEN_5653 = 14'h1615 == index ? 14'h102 : _GEN_5652;
  wire [13:0] _GEN_5654 = 14'h1616 == index ? 14'h100 : _GEN_5653;
  wire [13:0] _GEN_5655 = 14'h1617 == index ? 14'h95 : _GEN_5654;
  wire [13:0] _GEN_5656 = 14'h1618 == index ? 14'h94 : _GEN_5655;
  wire [13:0] _GEN_5657 = 14'h1619 == index ? 14'h93 : _GEN_5656;
  wire [13:0] _GEN_5658 = 14'h161a == index ? 14'h92 : _GEN_5657;
  wire [13:0] _GEN_5659 = 14'h161b == index ? 14'h91 : _GEN_5658;
  wire [13:0] _GEN_5660 = 14'h161c == index ? 14'h90 : _GEN_5659;
  wire [13:0] _GEN_5661 = 14'h161d == index ? 14'h8f : _GEN_5660;
  wire [13:0] _GEN_5662 = 14'h161e == index ? 14'h8e : _GEN_5661;
  wire [13:0] _GEN_5663 = 14'h161f == index ? 14'h8d : _GEN_5662;
  wire [13:0] _GEN_5664 = 14'h1620 == index ? 14'h8c : _GEN_5663;
  wire [13:0] _GEN_5665 = 14'h1621 == index ? 14'h8b : _GEN_5664;
  wire [13:0] _GEN_5666 = 14'h1622 == index ? 14'h8a : _GEN_5665;
  wire [13:0] _GEN_5667 = 14'h1623 == index ? 14'h89 : _GEN_5666;
  wire [13:0] _GEN_5668 = 14'h1624 == index ? 14'h88 : _GEN_5667;
  wire [13:0] _GEN_5669 = 14'h1625 == index ? 14'h87 : _GEN_5668;
  wire [13:0] _GEN_5670 = 14'h1626 == index ? 14'h86 : _GEN_5669;
  wire [13:0] _GEN_5671 = 14'h1627 == index ? 14'h85 : _GEN_5670;
  wire [13:0] _GEN_5672 = 14'h1628 == index ? 14'h84 : _GEN_5671;
  wire [13:0] _GEN_5673 = 14'h1629 == index ? 14'h83 : _GEN_5672;
  wire [13:0] _GEN_5674 = 14'h162a == index ? 14'h82 : _GEN_5673;
  wire [13:0] _GEN_5675 = 14'h162b == index ? 14'h81 : _GEN_5674;
  wire [13:0] _GEN_5676 = 14'h162c == index ? 14'h80 : _GEN_5675;
  wire [13:0] _GEN_5677 = 14'h162d == index ? 14'h2c : _GEN_5676;
  wire [13:0] _GEN_5678 = 14'h162e == index ? 14'h2c : _GEN_5677;
  wire [13:0] _GEN_5679 = 14'h162f == index ? 14'h2c : _GEN_5678;
  wire [13:0] _GEN_5680 = 14'h1630 == index ? 14'h2c : _GEN_5679;
  wire [13:0] _GEN_5681 = 14'h1631 == index ? 14'h2c : _GEN_5680;
  wire [13:0] _GEN_5682 = 14'h1632 == index ? 14'h2c : _GEN_5681;
  wire [13:0] _GEN_5683 = 14'h1633 == index ? 14'h2c : _GEN_5682;
  wire [13:0] _GEN_5684 = 14'h1634 == index ? 14'h2c : _GEN_5683;
  wire [13:0] _GEN_5685 = 14'h1635 == index ? 14'h2c : _GEN_5684;
  wire [13:0] _GEN_5686 = 14'h1636 == index ? 14'h2c : _GEN_5685;
  wire [13:0] _GEN_5687 = 14'h1637 == index ? 14'h2c : _GEN_5686;
  wire [13:0] _GEN_5688 = 14'h1638 == index ? 14'h2c : _GEN_5687;
  wire [13:0] _GEN_5689 = 14'h1639 == index ? 14'h2c : _GEN_5688;
  wire [13:0] _GEN_5690 = 14'h163a == index ? 14'h2c : _GEN_5689;
  wire [13:0] _GEN_5691 = 14'h163b == index ? 14'h2c : _GEN_5690;
  wire [13:0] _GEN_5692 = 14'h163c == index ? 14'h2c : _GEN_5691;
  wire [13:0] _GEN_5693 = 14'h163d == index ? 14'h2c : _GEN_5692;
  wire [13:0] _GEN_5694 = 14'h163e == index ? 14'h2c : _GEN_5693;
  wire [13:0] _GEN_5695 = 14'h163f == index ? 14'h2c : _GEN_5694;
  wire [13:0] _GEN_5696 = 14'h1640 == index ? 14'h2c : _GEN_5695;
  wire [13:0] _GEN_5697 = 14'h1641 == index ? 14'h2c : _GEN_5696;
  wire [13:0] _GEN_5698 = 14'h1642 == index ? 14'h2c : _GEN_5697;
  wire [13:0] _GEN_5699 = 14'h1643 == index ? 14'h2c : _GEN_5698;
  wire [13:0] _GEN_5700 = 14'h1644 == index ? 14'h2c : _GEN_5699;
  wire [13:0] _GEN_5701 = 14'h1645 == index ? 14'h2c : _GEN_5700;
  wire [13:0] _GEN_5702 = 14'h1646 == index ? 14'h2c : _GEN_5701;
  wire [13:0] _GEN_5703 = 14'h1647 == index ? 14'h2c : _GEN_5702;
  wire [13:0] _GEN_5704 = 14'h1648 == index ? 14'h2c : _GEN_5703;
  wire [13:0] _GEN_5705 = 14'h1649 == index ? 14'h2c : _GEN_5704;
  wire [13:0] _GEN_5706 = 14'h164a == index ? 14'h2c : _GEN_5705;
  wire [13:0] _GEN_5707 = 14'h164b == index ? 14'h2c : _GEN_5706;
  wire [13:0] _GEN_5708 = 14'h164c == index ? 14'h2c : _GEN_5707;
  wire [13:0] _GEN_5709 = 14'h164d == index ? 14'h2c : _GEN_5708;
  wire [13:0] _GEN_5710 = 14'h164e == index ? 14'h2c : _GEN_5709;
  wire [13:0] _GEN_5711 = 14'h164f == index ? 14'h2c : _GEN_5710;
  wire [13:0] _GEN_5712 = 14'h1650 == index ? 14'h2c : _GEN_5711;
  wire [13:0] _GEN_5713 = 14'h1651 == index ? 14'h2c : _GEN_5712;
  wire [13:0] _GEN_5714 = 14'h1652 == index ? 14'h2c : _GEN_5713;
  wire [13:0] _GEN_5715 = 14'h1653 == index ? 14'h2c : _GEN_5714;
  wire [13:0] _GEN_5716 = 14'h1654 == index ? 14'h2c : _GEN_5715;
  wire [13:0] _GEN_5717 = 14'h1655 == index ? 14'h2c : _GEN_5716;
  wire [13:0] _GEN_5718 = 14'h1656 == index ? 14'h2c : _GEN_5717;
  wire [13:0] _GEN_5719 = 14'h1657 == index ? 14'h2c : _GEN_5718;
  wire [13:0] _GEN_5720 = 14'h1658 == index ? 14'h2c : _GEN_5719;
  wire [13:0] _GEN_5721 = 14'h1659 == index ? 14'h2c : _GEN_5720;
  wire [13:0] _GEN_5722 = 14'h165a == index ? 14'h2c : _GEN_5721;
  wire [13:0] _GEN_5723 = 14'h165b == index ? 14'h2c : _GEN_5722;
  wire [13:0] _GEN_5724 = 14'h165c == index ? 14'h2c : _GEN_5723;
  wire [13:0] _GEN_5725 = 14'h165d == index ? 14'h2c : _GEN_5724;
  wire [13:0] _GEN_5726 = 14'h165e == index ? 14'h2c : _GEN_5725;
  wire [13:0] _GEN_5727 = 14'h165f == index ? 14'h2c : _GEN_5726;
  wire [13:0] _GEN_5728 = 14'h1660 == index ? 14'h2c : _GEN_5727;
  wire [13:0] _GEN_5729 = 14'h1661 == index ? 14'h2c : _GEN_5728;
  wire [13:0] _GEN_5730 = 14'h1662 == index ? 14'h2c : _GEN_5729;
  wire [13:0] _GEN_5731 = 14'h1663 == index ? 14'h2c : _GEN_5730;
  wire [13:0] _GEN_5732 = 14'h1664 == index ? 14'h2c : _GEN_5731;
  wire [13:0] _GEN_5733 = 14'h1665 == index ? 14'h2c : _GEN_5732;
  wire [13:0] _GEN_5734 = 14'h1666 == index ? 14'h2c : _GEN_5733;
  wire [13:0] _GEN_5735 = 14'h1667 == index ? 14'h2c : _GEN_5734;
  wire [13:0] _GEN_5736 = 14'h1668 == index ? 14'h2c : _GEN_5735;
  wire [13:0] _GEN_5737 = 14'h1669 == index ? 14'h2c : _GEN_5736;
  wire [13:0] _GEN_5738 = 14'h166a == index ? 14'h2c : _GEN_5737;
  wire [13:0] _GEN_5739 = 14'h166b == index ? 14'h2c : _GEN_5738;
  wire [13:0] _GEN_5740 = 14'h166c == index ? 14'h2c : _GEN_5739;
  wire [13:0] _GEN_5741 = 14'h166d == index ? 14'h2c : _GEN_5740;
  wire [13:0] _GEN_5742 = 14'h166e == index ? 14'h2c : _GEN_5741;
  wire [13:0] _GEN_5743 = 14'h166f == index ? 14'h2c : _GEN_5742;
  wire [13:0] _GEN_5744 = 14'h1670 == index ? 14'h2c : _GEN_5743;
  wire [13:0] _GEN_5745 = 14'h1671 == index ? 14'h2c : _GEN_5744;
  wire [13:0] _GEN_5746 = 14'h1672 == index ? 14'h2c : _GEN_5745;
  wire [13:0] _GEN_5747 = 14'h1673 == index ? 14'h2c : _GEN_5746;
  wire [13:0] _GEN_5748 = 14'h1674 == index ? 14'h2c : _GEN_5747;
  wire [13:0] _GEN_5749 = 14'h1675 == index ? 14'h2c : _GEN_5748;
  wire [13:0] _GEN_5750 = 14'h1676 == index ? 14'h2c : _GEN_5749;
  wire [13:0] _GEN_5751 = 14'h1677 == index ? 14'h2c : _GEN_5750;
  wire [13:0] _GEN_5752 = 14'h1678 == index ? 14'h2c : _GEN_5751;
  wire [13:0] _GEN_5753 = 14'h1679 == index ? 14'h2c : _GEN_5752;
  wire [13:0] _GEN_5754 = 14'h167a == index ? 14'h2c : _GEN_5753;
  wire [13:0] _GEN_5755 = 14'h167b == index ? 14'h2c : _GEN_5754;
  wire [13:0] _GEN_5756 = 14'h167c == index ? 14'h2c : _GEN_5755;
  wire [13:0] _GEN_5757 = 14'h167d == index ? 14'h2c : _GEN_5756;
  wire [13:0] _GEN_5758 = 14'h167e == index ? 14'h2c : _GEN_5757;
  wire [13:0] _GEN_5759 = 14'h167f == index ? 14'h2c : _GEN_5758;
  wire [13:0] _GEN_5760 = 14'h1680 == index ? 14'h0 : _GEN_5759;
  wire [13:0] _GEN_5761 = 14'h1681 == index ? 14'h1680 : _GEN_5760;
  wire [13:0] _GEN_5762 = 14'h1682 == index ? 14'hb01 : _GEN_5761;
  wire [13:0] _GEN_5763 = 14'h1683 == index ? 14'h780 : _GEN_5762;
  wire [13:0] _GEN_5764 = 14'h1684 == index ? 14'h581 : _GEN_5763;
  wire [13:0] _GEN_5765 = 14'h1685 == index ? 14'h480 : _GEN_5764;
  wire [13:0] _GEN_5766 = 14'h1686 == index ? 14'h383 : _GEN_5765;
  wire [13:0] _GEN_5767 = 14'h1687 == index ? 14'h303 : _GEN_5766;
  wire [13:0] _GEN_5768 = 14'h1688 == index ? 14'h285 : _GEN_5767;
  wire [13:0] _GEN_5769 = 14'h1689 == index ? 14'h280 : _GEN_5768;
  wire [13:0] _GEN_5770 = 14'h168a == index ? 14'h205 : _GEN_5769;
  wire [13:0] _GEN_5771 = 14'h168b == index ? 14'h201 : _GEN_5770;
  wire [13:0] _GEN_5772 = 14'h168c == index ? 14'h189 : _GEN_5771;
  wire [13:0] _GEN_5773 = 14'h168d == index ? 14'h186 : _GEN_5772;
  wire [13:0] _GEN_5774 = 14'h168e == index ? 14'h183 : _GEN_5773;
  wire [13:0] _GEN_5775 = 14'h168f == index ? 14'h180 : _GEN_5774;
  wire [13:0] _GEN_5776 = 14'h1690 == index ? 14'h10d : _GEN_5775;
  wire [13:0] _GEN_5777 = 14'h1691 == index ? 14'h10b : _GEN_5776;
  wire [13:0] _GEN_5778 = 14'h1692 == index ? 14'h109 : _GEN_5777;
  wire [13:0] _GEN_5779 = 14'h1693 == index ? 14'h107 : _GEN_5778;
  wire [13:0] _GEN_5780 = 14'h1694 == index ? 14'h105 : _GEN_5779;
  wire [13:0] _GEN_5781 = 14'h1695 == index ? 14'h103 : _GEN_5780;
  wire [13:0] _GEN_5782 = 14'h1696 == index ? 14'h101 : _GEN_5781;
  wire [13:0] _GEN_5783 = 14'h1697 == index ? 14'h96 : _GEN_5782;
  wire [13:0] _GEN_5784 = 14'h1698 == index ? 14'h95 : _GEN_5783;
  wire [13:0] _GEN_5785 = 14'h1699 == index ? 14'h94 : _GEN_5784;
  wire [13:0] _GEN_5786 = 14'h169a == index ? 14'h93 : _GEN_5785;
  wire [13:0] _GEN_5787 = 14'h169b == index ? 14'h92 : _GEN_5786;
  wire [13:0] _GEN_5788 = 14'h169c == index ? 14'h91 : _GEN_5787;
  wire [13:0] _GEN_5789 = 14'h169d == index ? 14'h90 : _GEN_5788;
  wire [13:0] _GEN_5790 = 14'h169e == index ? 14'h8f : _GEN_5789;
  wire [13:0] _GEN_5791 = 14'h169f == index ? 14'h8e : _GEN_5790;
  wire [13:0] _GEN_5792 = 14'h16a0 == index ? 14'h8d : _GEN_5791;
  wire [13:0] _GEN_5793 = 14'h16a1 == index ? 14'h8c : _GEN_5792;
  wire [13:0] _GEN_5794 = 14'h16a2 == index ? 14'h8b : _GEN_5793;
  wire [13:0] _GEN_5795 = 14'h16a3 == index ? 14'h8a : _GEN_5794;
  wire [13:0] _GEN_5796 = 14'h16a4 == index ? 14'h89 : _GEN_5795;
  wire [13:0] _GEN_5797 = 14'h16a5 == index ? 14'h88 : _GEN_5796;
  wire [13:0] _GEN_5798 = 14'h16a6 == index ? 14'h87 : _GEN_5797;
  wire [13:0] _GEN_5799 = 14'h16a7 == index ? 14'h86 : _GEN_5798;
  wire [13:0] _GEN_5800 = 14'h16a8 == index ? 14'h85 : _GEN_5799;
  wire [13:0] _GEN_5801 = 14'h16a9 == index ? 14'h84 : _GEN_5800;
  wire [13:0] _GEN_5802 = 14'h16aa == index ? 14'h83 : _GEN_5801;
  wire [13:0] _GEN_5803 = 14'h16ab == index ? 14'h82 : _GEN_5802;
  wire [13:0] _GEN_5804 = 14'h16ac == index ? 14'h81 : _GEN_5803;
  wire [13:0] _GEN_5805 = 14'h16ad == index ? 14'h80 : _GEN_5804;
  wire [13:0] _GEN_5806 = 14'h16ae == index ? 14'h2d : _GEN_5805;
  wire [13:0] _GEN_5807 = 14'h16af == index ? 14'h2d : _GEN_5806;
  wire [13:0] _GEN_5808 = 14'h16b0 == index ? 14'h2d : _GEN_5807;
  wire [13:0] _GEN_5809 = 14'h16b1 == index ? 14'h2d : _GEN_5808;
  wire [13:0] _GEN_5810 = 14'h16b2 == index ? 14'h2d : _GEN_5809;
  wire [13:0] _GEN_5811 = 14'h16b3 == index ? 14'h2d : _GEN_5810;
  wire [13:0] _GEN_5812 = 14'h16b4 == index ? 14'h2d : _GEN_5811;
  wire [13:0] _GEN_5813 = 14'h16b5 == index ? 14'h2d : _GEN_5812;
  wire [13:0] _GEN_5814 = 14'h16b6 == index ? 14'h2d : _GEN_5813;
  wire [13:0] _GEN_5815 = 14'h16b7 == index ? 14'h2d : _GEN_5814;
  wire [13:0] _GEN_5816 = 14'h16b8 == index ? 14'h2d : _GEN_5815;
  wire [13:0] _GEN_5817 = 14'h16b9 == index ? 14'h2d : _GEN_5816;
  wire [13:0] _GEN_5818 = 14'h16ba == index ? 14'h2d : _GEN_5817;
  wire [13:0] _GEN_5819 = 14'h16bb == index ? 14'h2d : _GEN_5818;
  wire [13:0] _GEN_5820 = 14'h16bc == index ? 14'h2d : _GEN_5819;
  wire [13:0] _GEN_5821 = 14'h16bd == index ? 14'h2d : _GEN_5820;
  wire [13:0] _GEN_5822 = 14'h16be == index ? 14'h2d : _GEN_5821;
  wire [13:0] _GEN_5823 = 14'h16bf == index ? 14'h2d : _GEN_5822;
  wire [13:0] _GEN_5824 = 14'h16c0 == index ? 14'h2d : _GEN_5823;
  wire [13:0] _GEN_5825 = 14'h16c1 == index ? 14'h2d : _GEN_5824;
  wire [13:0] _GEN_5826 = 14'h16c2 == index ? 14'h2d : _GEN_5825;
  wire [13:0] _GEN_5827 = 14'h16c3 == index ? 14'h2d : _GEN_5826;
  wire [13:0] _GEN_5828 = 14'h16c4 == index ? 14'h2d : _GEN_5827;
  wire [13:0] _GEN_5829 = 14'h16c5 == index ? 14'h2d : _GEN_5828;
  wire [13:0] _GEN_5830 = 14'h16c6 == index ? 14'h2d : _GEN_5829;
  wire [13:0] _GEN_5831 = 14'h16c7 == index ? 14'h2d : _GEN_5830;
  wire [13:0] _GEN_5832 = 14'h16c8 == index ? 14'h2d : _GEN_5831;
  wire [13:0] _GEN_5833 = 14'h16c9 == index ? 14'h2d : _GEN_5832;
  wire [13:0] _GEN_5834 = 14'h16ca == index ? 14'h2d : _GEN_5833;
  wire [13:0] _GEN_5835 = 14'h16cb == index ? 14'h2d : _GEN_5834;
  wire [13:0] _GEN_5836 = 14'h16cc == index ? 14'h2d : _GEN_5835;
  wire [13:0] _GEN_5837 = 14'h16cd == index ? 14'h2d : _GEN_5836;
  wire [13:0] _GEN_5838 = 14'h16ce == index ? 14'h2d : _GEN_5837;
  wire [13:0] _GEN_5839 = 14'h16cf == index ? 14'h2d : _GEN_5838;
  wire [13:0] _GEN_5840 = 14'h16d0 == index ? 14'h2d : _GEN_5839;
  wire [13:0] _GEN_5841 = 14'h16d1 == index ? 14'h2d : _GEN_5840;
  wire [13:0] _GEN_5842 = 14'h16d2 == index ? 14'h2d : _GEN_5841;
  wire [13:0] _GEN_5843 = 14'h16d3 == index ? 14'h2d : _GEN_5842;
  wire [13:0] _GEN_5844 = 14'h16d4 == index ? 14'h2d : _GEN_5843;
  wire [13:0] _GEN_5845 = 14'h16d5 == index ? 14'h2d : _GEN_5844;
  wire [13:0] _GEN_5846 = 14'h16d6 == index ? 14'h2d : _GEN_5845;
  wire [13:0] _GEN_5847 = 14'h16d7 == index ? 14'h2d : _GEN_5846;
  wire [13:0] _GEN_5848 = 14'h16d8 == index ? 14'h2d : _GEN_5847;
  wire [13:0] _GEN_5849 = 14'h16d9 == index ? 14'h2d : _GEN_5848;
  wire [13:0] _GEN_5850 = 14'h16da == index ? 14'h2d : _GEN_5849;
  wire [13:0] _GEN_5851 = 14'h16db == index ? 14'h2d : _GEN_5850;
  wire [13:0] _GEN_5852 = 14'h16dc == index ? 14'h2d : _GEN_5851;
  wire [13:0] _GEN_5853 = 14'h16dd == index ? 14'h2d : _GEN_5852;
  wire [13:0] _GEN_5854 = 14'h16de == index ? 14'h2d : _GEN_5853;
  wire [13:0] _GEN_5855 = 14'h16df == index ? 14'h2d : _GEN_5854;
  wire [13:0] _GEN_5856 = 14'h16e0 == index ? 14'h2d : _GEN_5855;
  wire [13:0] _GEN_5857 = 14'h16e1 == index ? 14'h2d : _GEN_5856;
  wire [13:0] _GEN_5858 = 14'h16e2 == index ? 14'h2d : _GEN_5857;
  wire [13:0] _GEN_5859 = 14'h16e3 == index ? 14'h2d : _GEN_5858;
  wire [13:0] _GEN_5860 = 14'h16e4 == index ? 14'h2d : _GEN_5859;
  wire [13:0] _GEN_5861 = 14'h16e5 == index ? 14'h2d : _GEN_5860;
  wire [13:0] _GEN_5862 = 14'h16e6 == index ? 14'h2d : _GEN_5861;
  wire [13:0] _GEN_5863 = 14'h16e7 == index ? 14'h2d : _GEN_5862;
  wire [13:0] _GEN_5864 = 14'h16e8 == index ? 14'h2d : _GEN_5863;
  wire [13:0] _GEN_5865 = 14'h16e9 == index ? 14'h2d : _GEN_5864;
  wire [13:0] _GEN_5866 = 14'h16ea == index ? 14'h2d : _GEN_5865;
  wire [13:0] _GEN_5867 = 14'h16eb == index ? 14'h2d : _GEN_5866;
  wire [13:0] _GEN_5868 = 14'h16ec == index ? 14'h2d : _GEN_5867;
  wire [13:0] _GEN_5869 = 14'h16ed == index ? 14'h2d : _GEN_5868;
  wire [13:0] _GEN_5870 = 14'h16ee == index ? 14'h2d : _GEN_5869;
  wire [13:0] _GEN_5871 = 14'h16ef == index ? 14'h2d : _GEN_5870;
  wire [13:0] _GEN_5872 = 14'h16f0 == index ? 14'h2d : _GEN_5871;
  wire [13:0] _GEN_5873 = 14'h16f1 == index ? 14'h2d : _GEN_5872;
  wire [13:0] _GEN_5874 = 14'h16f2 == index ? 14'h2d : _GEN_5873;
  wire [13:0] _GEN_5875 = 14'h16f3 == index ? 14'h2d : _GEN_5874;
  wire [13:0] _GEN_5876 = 14'h16f4 == index ? 14'h2d : _GEN_5875;
  wire [13:0] _GEN_5877 = 14'h16f5 == index ? 14'h2d : _GEN_5876;
  wire [13:0] _GEN_5878 = 14'h16f6 == index ? 14'h2d : _GEN_5877;
  wire [13:0] _GEN_5879 = 14'h16f7 == index ? 14'h2d : _GEN_5878;
  wire [13:0] _GEN_5880 = 14'h16f8 == index ? 14'h2d : _GEN_5879;
  wire [13:0] _GEN_5881 = 14'h16f9 == index ? 14'h2d : _GEN_5880;
  wire [13:0] _GEN_5882 = 14'h16fa == index ? 14'h2d : _GEN_5881;
  wire [13:0] _GEN_5883 = 14'h16fb == index ? 14'h2d : _GEN_5882;
  wire [13:0] _GEN_5884 = 14'h16fc == index ? 14'h2d : _GEN_5883;
  wire [13:0] _GEN_5885 = 14'h16fd == index ? 14'h2d : _GEN_5884;
  wire [13:0] _GEN_5886 = 14'h16fe == index ? 14'h2d : _GEN_5885;
  wire [13:0] _GEN_5887 = 14'h16ff == index ? 14'h2d : _GEN_5886;
  wire [13:0] _GEN_5888 = 14'h1700 == index ? 14'h0 : _GEN_5887;
  wire [13:0] _GEN_5889 = 14'h1701 == index ? 14'h1700 : _GEN_5888;
  wire [13:0] _GEN_5890 = 14'h1702 == index ? 14'hb80 : _GEN_5889;
  wire [13:0] _GEN_5891 = 14'h1703 == index ? 14'h781 : _GEN_5890;
  wire [13:0] _GEN_5892 = 14'h1704 == index ? 14'h582 : _GEN_5891;
  wire [13:0] _GEN_5893 = 14'h1705 == index ? 14'h481 : _GEN_5892;
  wire [13:0] _GEN_5894 = 14'h1706 == index ? 14'h384 : _GEN_5893;
  wire [13:0] _GEN_5895 = 14'h1707 == index ? 14'h304 : _GEN_5894;
  wire [13:0] _GEN_5896 = 14'h1708 == index ? 14'h286 : _GEN_5895;
  wire [13:0] _GEN_5897 = 14'h1709 == index ? 14'h281 : _GEN_5896;
  wire [13:0] _GEN_5898 = 14'h170a == index ? 14'h206 : _GEN_5897;
  wire [13:0] _GEN_5899 = 14'h170b == index ? 14'h202 : _GEN_5898;
  wire [13:0] _GEN_5900 = 14'h170c == index ? 14'h18a : _GEN_5899;
  wire [13:0] _GEN_5901 = 14'h170d == index ? 14'h187 : _GEN_5900;
  wire [13:0] _GEN_5902 = 14'h170e == index ? 14'h184 : _GEN_5901;
  wire [13:0] _GEN_5903 = 14'h170f == index ? 14'h181 : _GEN_5902;
  wire [13:0] _GEN_5904 = 14'h1710 == index ? 14'h10e : _GEN_5903;
  wire [13:0] _GEN_5905 = 14'h1711 == index ? 14'h10c : _GEN_5904;
  wire [13:0] _GEN_5906 = 14'h1712 == index ? 14'h10a : _GEN_5905;
  wire [13:0] _GEN_5907 = 14'h1713 == index ? 14'h108 : _GEN_5906;
  wire [13:0] _GEN_5908 = 14'h1714 == index ? 14'h106 : _GEN_5907;
  wire [13:0] _GEN_5909 = 14'h1715 == index ? 14'h104 : _GEN_5908;
  wire [13:0] _GEN_5910 = 14'h1716 == index ? 14'h102 : _GEN_5909;
  wire [13:0] _GEN_5911 = 14'h1717 == index ? 14'h100 : _GEN_5910;
  wire [13:0] _GEN_5912 = 14'h1718 == index ? 14'h96 : _GEN_5911;
  wire [13:0] _GEN_5913 = 14'h1719 == index ? 14'h95 : _GEN_5912;
  wire [13:0] _GEN_5914 = 14'h171a == index ? 14'h94 : _GEN_5913;
  wire [13:0] _GEN_5915 = 14'h171b == index ? 14'h93 : _GEN_5914;
  wire [13:0] _GEN_5916 = 14'h171c == index ? 14'h92 : _GEN_5915;
  wire [13:0] _GEN_5917 = 14'h171d == index ? 14'h91 : _GEN_5916;
  wire [13:0] _GEN_5918 = 14'h171e == index ? 14'h90 : _GEN_5917;
  wire [13:0] _GEN_5919 = 14'h171f == index ? 14'h8f : _GEN_5918;
  wire [13:0] _GEN_5920 = 14'h1720 == index ? 14'h8e : _GEN_5919;
  wire [13:0] _GEN_5921 = 14'h1721 == index ? 14'h8d : _GEN_5920;
  wire [13:0] _GEN_5922 = 14'h1722 == index ? 14'h8c : _GEN_5921;
  wire [13:0] _GEN_5923 = 14'h1723 == index ? 14'h8b : _GEN_5922;
  wire [13:0] _GEN_5924 = 14'h1724 == index ? 14'h8a : _GEN_5923;
  wire [13:0] _GEN_5925 = 14'h1725 == index ? 14'h89 : _GEN_5924;
  wire [13:0] _GEN_5926 = 14'h1726 == index ? 14'h88 : _GEN_5925;
  wire [13:0] _GEN_5927 = 14'h1727 == index ? 14'h87 : _GEN_5926;
  wire [13:0] _GEN_5928 = 14'h1728 == index ? 14'h86 : _GEN_5927;
  wire [13:0] _GEN_5929 = 14'h1729 == index ? 14'h85 : _GEN_5928;
  wire [13:0] _GEN_5930 = 14'h172a == index ? 14'h84 : _GEN_5929;
  wire [13:0] _GEN_5931 = 14'h172b == index ? 14'h83 : _GEN_5930;
  wire [13:0] _GEN_5932 = 14'h172c == index ? 14'h82 : _GEN_5931;
  wire [13:0] _GEN_5933 = 14'h172d == index ? 14'h81 : _GEN_5932;
  wire [13:0] _GEN_5934 = 14'h172e == index ? 14'h80 : _GEN_5933;
  wire [13:0] _GEN_5935 = 14'h172f == index ? 14'h2e : _GEN_5934;
  wire [13:0] _GEN_5936 = 14'h1730 == index ? 14'h2e : _GEN_5935;
  wire [13:0] _GEN_5937 = 14'h1731 == index ? 14'h2e : _GEN_5936;
  wire [13:0] _GEN_5938 = 14'h1732 == index ? 14'h2e : _GEN_5937;
  wire [13:0] _GEN_5939 = 14'h1733 == index ? 14'h2e : _GEN_5938;
  wire [13:0] _GEN_5940 = 14'h1734 == index ? 14'h2e : _GEN_5939;
  wire [13:0] _GEN_5941 = 14'h1735 == index ? 14'h2e : _GEN_5940;
  wire [13:0] _GEN_5942 = 14'h1736 == index ? 14'h2e : _GEN_5941;
  wire [13:0] _GEN_5943 = 14'h1737 == index ? 14'h2e : _GEN_5942;
  wire [13:0] _GEN_5944 = 14'h1738 == index ? 14'h2e : _GEN_5943;
  wire [13:0] _GEN_5945 = 14'h1739 == index ? 14'h2e : _GEN_5944;
  wire [13:0] _GEN_5946 = 14'h173a == index ? 14'h2e : _GEN_5945;
  wire [13:0] _GEN_5947 = 14'h173b == index ? 14'h2e : _GEN_5946;
  wire [13:0] _GEN_5948 = 14'h173c == index ? 14'h2e : _GEN_5947;
  wire [13:0] _GEN_5949 = 14'h173d == index ? 14'h2e : _GEN_5948;
  wire [13:0] _GEN_5950 = 14'h173e == index ? 14'h2e : _GEN_5949;
  wire [13:0] _GEN_5951 = 14'h173f == index ? 14'h2e : _GEN_5950;
  wire [13:0] _GEN_5952 = 14'h1740 == index ? 14'h2e : _GEN_5951;
  wire [13:0] _GEN_5953 = 14'h1741 == index ? 14'h2e : _GEN_5952;
  wire [13:0] _GEN_5954 = 14'h1742 == index ? 14'h2e : _GEN_5953;
  wire [13:0] _GEN_5955 = 14'h1743 == index ? 14'h2e : _GEN_5954;
  wire [13:0] _GEN_5956 = 14'h1744 == index ? 14'h2e : _GEN_5955;
  wire [13:0] _GEN_5957 = 14'h1745 == index ? 14'h2e : _GEN_5956;
  wire [13:0] _GEN_5958 = 14'h1746 == index ? 14'h2e : _GEN_5957;
  wire [13:0] _GEN_5959 = 14'h1747 == index ? 14'h2e : _GEN_5958;
  wire [13:0] _GEN_5960 = 14'h1748 == index ? 14'h2e : _GEN_5959;
  wire [13:0] _GEN_5961 = 14'h1749 == index ? 14'h2e : _GEN_5960;
  wire [13:0] _GEN_5962 = 14'h174a == index ? 14'h2e : _GEN_5961;
  wire [13:0] _GEN_5963 = 14'h174b == index ? 14'h2e : _GEN_5962;
  wire [13:0] _GEN_5964 = 14'h174c == index ? 14'h2e : _GEN_5963;
  wire [13:0] _GEN_5965 = 14'h174d == index ? 14'h2e : _GEN_5964;
  wire [13:0] _GEN_5966 = 14'h174e == index ? 14'h2e : _GEN_5965;
  wire [13:0] _GEN_5967 = 14'h174f == index ? 14'h2e : _GEN_5966;
  wire [13:0] _GEN_5968 = 14'h1750 == index ? 14'h2e : _GEN_5967;
  wire [13:0] _GEN_5969 = 14'h1751 == index ? 14'h2e : _GEN_5968;
  wire [13:0] _GEN_5970 = 14'h1752 == index ? 14'h2e : _GEN_5969;
  wire [13:0] _GEN_5971 = 14'h1753 == index ? 14'h2e : _GEN_5970;
  wire [13:0] _GEN_5972 = 14'h1754 == index ? 14'h2e : _GEN_5971;
  wire [13:0] _GEN_5973 = 14'h1755 == index ? 14'h2e : _GEN_5972;
  wire [13:0] _GEN_5974 = 14'h1756 == index ? 14'h2e : _GEN_5973;
  wire [13:0] _GEN_5975 = 14'h1757 == index ? 14'h2e : _GEN_5974;
  wire [13:0] _GEN_5976 = 14'h1758 == index ? 14'h2e : _GEN_5975;
  wire [13:0] _GEN_5977 = 14'h1759 == index ? 14'h2e : _GEN_5976;
  wire [13:0] _GEN_5978 = 14'h175a == index ? 14'h2e : _GEN_5977;
  wire [13:0] _GEN_5979 = 14'h175b == index ? 14'h2e : _GEN_5978;
  wire [13:0] _GEN_5980 = 14'h175c == index ? 14'h2e : _GEN_5979;
  wire [13:0] _GEN_5981 = 14'h175d == index ? 14'h2e : _GEN_5980;
  wire [13:0] _GEN_5982 = 14'h175e == index ? 14'h2e : _GEN_5981;
  wire [13:0] _GEN_5983 = 14'h175f == index ? 14'h2e : _GEN_5982;
  wire [13:0] _GEN_5984 = 14'h1760 == index ? 14'h2e : _GEN_5983;
  wire [13:0] _GEN_5985 = 14'h1761 == index ? 14'h2e : _GEN_5984;
  wire [13:0] _GEN_5986 = 14'h1762 == index ? 14'h2e : _GEN_5985;
  wire [13:0] _GEN_5987 = 14'h1763 == index ? 14'h2e : _GEN_5986;
  wire [13:0] _GEN_5988 = 14'h1764 == index ? 14'h2e : _GEN_5987;
  wire [13:0] _GEN_5989 = 14'h1765 == index ? 14'h2e : _GEN_5988;
  wire [13:0] _GEN_5990 = 14'h1766 == index ? 14'h2e : _GEN_5989;
  wire [13:0] _GEN_5991 = 14'h1767 == index ? 14'h2e : _GEN_5990;
  wire [13:0] _GEN_5992 = 14'h1768 == index ? 14'h2e : _GEN_5991;
  wire [13:0] _GEN_5993 = 14'h1769 == index ? 14'h2e : _GEN_5992;
  wire [13:0] _GEN_5994 = 14'h176a == index ? 14'h2e : _GEN_5993;
  wire [13:0] _GEN_5995 = 14'h176b == index ? 14'h2e : _GEN_5994;
  wire [13:0] _GEN_5996 = 14'h176c == index ? 14'h2e : _GEN_5995;
  wire [13:0] _GEN_5997 = 14'h176d == index ? 14'h2e : _GEN_5996;
  wire [13:0] _GEN_5998 = 14'h176e == index ? 14'h2e : _GEN_5997;
  wire [13:0] _GEN_5999 = 14'h176f == index ? 14'h2e : _GEN_5998;
  wire [13:0] _GEN_6000 = 14'h1770 == index ? 14'h2e : _GEN_5999;
  wire [13:0] _GEN_6001 = 14'h1771 == index ? 14'h2e : _GEN_6000;
  wire [13:0] _GEN_6002 = 14'h1772 == index ? 14'h2e : _GEN_6001;
  wire [13:0] _GEN_6003 = 14'h1773 == index ? 14'h2e : _GEN_6002;
  wire [13:0] _GEN_6004 = 14'h1774 == index ? 14'h2e : _GEN_6003;
  wire [13:0] _GEN_6005 = 14'h1775 == index ? 14'h2e : _GEN_6004;
  wire [13:0] _GEN_6006 = 14'h1776 == index ? 14'h2e : _GEN_6005;
  wire [13:0] _GEN_6007 = 14'h1777 == index ? 14'h2e : _GEN_6006;
  wire [13:0] _GEN_6008 = 14'h1778 == index ? 14'h2e : _GEN_6007;
  wire [13:0] _GEN_6009 = 14'h1779 == index ? 14'h2e : _GEN_6008;
  wire [13:0] _GEN_6010 = 14'h177a == index ? 14'h2e : _GEN_6009;
  wire [13:0] _GEN_6011 = 14'h177b == index ? 14'h2e : _GEN_6010;
  wire [13:0] _GEN_6012 = 14'h177c == index ? 14'h2e : _GEN_6011;
  wire [13:0] _GEN_6013 = 14'h177d == index ? 14'h2e : _GEN_6012;
  wire [13:0] _GEN_6014 = 14'h177e == index ? 14'h2e : _GEN_6013;
  wire [13:0] _GEN_6015 = 14'h177f == index ? 14'h2e : _GEN_6014;
  wire [13:0] _GEN_6016 = 14'h1780 == index ? 14'h0 : _GEN_6015;
  wire [13:0] _GEN_6017 = 14'h1781 == index ? 14'h1780 : _GEN_6016;
  wire [13:0] _GEN_6018 = 14'h1782 == index ? 14'hb81 : _GEN_6017;
  wire [13:0] _GEN_6019 = 14'h1783 == index ? 14'h782 : _GEN_6018;
  wire [13:0] _GEN_6020 = 14'h1784 == index ? 14'h583 : _GEN_6019;
  wire [13:0] _GEN_6021 = 14'h1785 == index ? 14'h482 : _GEN_6020;
  wire [13:0] _GEN_6022 = 14'h1786 == index ? 14'h385 : _GEN_6021;
  wire [13:0] _GEN_6023 = 14'h1787 == index ? 14'h305 : _GEN_6022;
  wire [13:0] _GEN_6024 = 14'h1788 == index ? 14'h287 : _GEN_6023;
  wire [13:0] _GEN_6025 = 14'h1789 == index ? 14'h282 : _GEN_6024;
  wire [13:0] _GEN_6026 = 14'h178a == index ? 14'h207 : _GEN_6025;
  wire [13:0] _GEN_6027 = 14'h178b == index ? 14'h203 : _GEN_6026;
  wire [13:0] _GEN_6028 = 14'h178c == index ? 14'h18b : _GEN_6027;
  wire [13:0] _GEN_6029 = 14'h178d == index ? 14'h188 : _GEN_6028;
  wire [13:0] _GEN_6030 = 14'h178e == index ? 14'h185 : _GEN_6029;
  wire [13:0] _GEN_6031 = 14'h178f == index ? 14'h182 : _GEN_6030;
  wire [13:0] _GEN_6032 = 14'h1790 == index ? 14'h10f : _GEN_6031;
  wire [13:0] _GEN_6033 = 14'h1791 == index ? 14'h10d : _GEN_6032;
  wire [13:0] _GEN_6034 = 14'h1792 == index ? 14'h10b : _GEN_6033;
  wire [13:0] _GEN_6035 = 14'h1793 == index ? 14'h109 : _GEN_6034;
  wire [13:0] _GEN_6036 = 14'h1794 == index ? 14'h107 : _GEN_6035;
  wire [13:0] _GEN_6037 = 14'h1795 == index ? 14'h105 : _GEN_6036;
  wire [13:0] _GEN_6038 = 14'h1796 == index ? 14'h103 : _GEN_6037;
  wire [13:0] _GEN_6039 = 14'h1797 == index ? 14'h101 : _GEN_6038;
  wire [13:0] _GEN_6040 = 14'h1798 == index ? 14'h97 : _GEN_6039;
  wire [13:0] _GEN_6041 = 14'h1799 == index ? 14'h96 : _GEN_6040;
  wire [13:0] _GEN_6042 = 14'h179a == index ? 14'h95 : _GEN_6041;
  wire [13:0] _GEN_6043 = 14'h179b == index ? 14'h94 : _GEN_6042;
  wire [13:0] _GEN_6044 = 14'h179c == index ? 14'h93 : _GEN_6043;
  wire [13:0] _GEN_6045 = 14'h179d == index ? 14'h92 : _GEN_6044;
  wire [13:0] _GEN_6046 = 14'h179e == index ? 14'h91 : _GEN_6045;
  wire [13:0] _GEN_6047 = 14'h179f == index ? 14'h90 : _GEN_6046;
  wire [13:0] _GEN_6048 = 14'h17a0 == index ? 14'h8f : _GEN_6047;
  wire [13:0] _GEN_6049 = 14'h17a1 == index ? 14'h8e : _GEN_6048;
  wire [13:0] _GEN_6050 = 14'h17a2 == index ? 14'h8d : _GEN_6049;
  wire [13:0] _GEN_6051 = 14'h17a3 == index ? 14'h8c : _GEN_6050;
  wire [13:0] _GEN_6052 = 14'h17a4 == index ? 14'h8b : _GEN_6051;
  wire [13:0] _GEN_6053 = 14'h17a5 == index ? 14'h8a : _GEN_6052;
  wire [13:0] _GEN_6054 = 14'h17a6 == index ? 14'h89 : _GEN_6053;
  wire [13:0] _GEN_6055 = 14'h17a7 == index ? 14'h88 : _GEN_6054;
  wire [13:0] _GEN_6056 = 14'h17a8 == index ? 14'h87 : _GEN_6055;
  wire [13:0] _GEN_6057 = 14'h17a9 == index ? 14'h86 : _GEN_6056;
  wire [13:0] _GEN_6058 = 14'h17aa == index ? 14'h85 : _GEN_6057;
  wire [13:0] _GEN_6059 = 14'h17ab == index ? 14'h84 : _GEN_6058;
  wire [13:0] _GEN_6060 = 14'h17ac == index ? 14'h83 : _GEN_6059;
  wire [13:0] _GEN_6061 = 14'h17ad == index ? 14'h82 : _GEN_6060;
  wire [13:0] _GEN_6062 = 14'h17ae == index ? 14'h81 : _GEN_6061;
  wire [13:0] _GEN_6063 = 14'h17af == index ? 14'h80 : _GEN_6062;
  wire [13:0] _GEN_6064 = 14'h17b0 == index ? 14'h2f : _GEN_6063;
  wire [13:0] _GEN_6065 = 14'h17b1 == index ? 14'h2f : _GEN_6064;
  wire [13:0] _GEN_6066 = 14'h17b2 == index ? 14'h2f : _GEN_6065;
  wire [13:0] _GEN_6067 = 14'h17b3 == index ? 14'h2f : _GEN_6066;
  wire [13:0] _GEN_6068 = 14'h17b4 == index ? 14'h2f : _GEN_6067;
  wire [13:0] _GEN_6069 = 14'h17b5 == index ? 14'h2f : _GEN_6068;
  wire [13:0] _GEN_6070 = 14'h17b6 == index ? 14'h2f : _GEN_6069;
  wire [13:0] _GEN_6071 = 14'h17b7 == index ? 14'h2f : _GEN_6070;
  wire [13:0] _GEN_6072 = 14'h17b8 == index ? 14'h2f : _GEN_6071;
  wire [13:0] _GEN_6073 = 14'h17b9 == index ? 14'h2f : _GEN_6072;
  wire [13:0] _GEN_6074 = 14'h17ba == index ? 14'h2f : _GEN_6073;
  wire [13:0] _GEN_6075 = 14'h17bb == index ? 14'h2f : _GEN_6074;
  wire [13:0] _GEN_6076 = 14'h17bc == index ? 14'h2f : _GEN_6075;
  wire [13:0] _GEN_6077 = 14'h17bd == index ? 14'h2f : _GEN_6076;
  wire [13:0] _GEN_6078 = 14'h17be == index ? 14'h2f : _GEN_6077;
  wire [13:0] _GEN_6079 = 14'h17bf == index ? 14'h2f : _GEN_6078;
  wire [13:0] _GEN_6080 = 14'h17c0 == index ? 14'h2f : _GEN_6079;
  wire [13:0] _GEN_6081 = 14'h17c1 == index ? 14'h2f : _GEN_6080;
  wire [13:0] _GEN_6082 = 14'h17c2 == index ? 14'h2f : _GEN_6081;
  wire [13:0] _GEN_6083 = 14'h17c3 == index ? 14'h2f : _GEN_6082;
  wire [13:0] _GEN_6084 = 14'h17c4 == index ? 14'h2f : _GEN_6083;
  wire [13:0] _GEN_6085 = 14'h17c5 == index ? 14'h2f : _GEN_6084;
  wire [13:0] _GEN_6086 = 14'h17c6 == index ? 14'h2f : _GEN_6085;
  wire [13:0] _GEN_6087 = 14'h17c7 == index ? 14'h2f : _GEN_6086;
  wire [13:0] _GEN_6088 = 14'h17c8 == index ? 14'h2f : _GEN_6087;
  wire [13:0] _GEN_6089 = 14'h17c9 == index ? 14'h2f : _GEN_6088;
  wire [13:0] _GEN_6090 = 14'h17ca == index ? 14'h2f : _GEN_6089;
  wire [13:0] _GEN_6091 = 14'h17cb == index ? 14'h2f : _GEN_6090;
  wire [13:0] _GEN_6092 = 14'h17cc == index ? 14'h2f : _GEN_6091;
  wire [13:0] _GEN_6093 = 14'h17cd == index ? 14'h2f : _GEN_6092;
  wire [13:0] _GEN_6094 = 14'h17ce == index ? 14'h2f : _GEN_6093;
  wire [13:0] _GEN_6095 = 14'h17cf == index ? 14'h2f : _GEN_6094;
  wire [13:0] _GEN_6096 = 14'h17d0 == index ? 14'h2f : _GEN_6095;
  wire [13:0] _GEN_6097 = 14'h17d1 == index ? 14'h2f : _GEN_6096;
  wire [13:0] _GEN_6098 = 14'h17d2 == index ? 14'h2f : _GEN_6097;
  wire [13:0] _GEN_6099 = 14'h17d3 == index ? 14'h2f : _GEN_6098;
  wire [13:0] _GEN_6100 = 14'h17d4 == index ? 14'h2f : _GEN_6099;
  wire [13:0] _GEN_6101 = 14'h17d5 == index ? 14'h2f : _GEN_6100;
  wire [13:0] _GEN_6102 = 14'h17d6 == index ? 14'h2f : _GEN_6101;
  wire [13:0] _GEN_6103 = 14'h17d7 == index ? 14'h2f : _GEN_6102;
  wire [13:0] _GEN_6104 = 14'h17d8 == index ? 14'h2f : _GEN_6103;
  wire [13:0] _GEN_6105 = 14'h17d9 == index ? 14'h2f : _GEN_6104;
  wire [13:0] _GEN_6106 = 14'h17da == index ? 14'h2f : _GEN_6105;
  wire [13:0] _GEN_6107 = 14'h17db == index ? 14'h2f : _GEN_6106;
  wire [13:0] _GEN_6108 = 14'h17dc == index ? 14'h2f : _GEN_6107;
  wire [13:0] _GEN_6109 = 14'h17dd == index ? 14'h2f : _GEN_6108;
  wire [13:0] _GEN_6110 = 14'h17de == index ? 14'h2f : _GEN_6109;
  wire [13:0] _GEN_6111 = 14'h17df == index ? 14'h2f : _GEN_6110;
  wire [13:0] _GEN_6112 = 14'h17e0 == index ? 14'h2f : _GEN_6111;
  wire [13:0] _GEN_6113 = 14'h17e1 == index ? 14'h2f : _GEN_6112;
  wire [13:0] _GEN_6114 = 14'h17e2 == index ? 14'h2f : _GEN_6113;
  wire [13:0] _GEN_6115 = 14'h17e3 == index ? 14'h2f : _GEN_6114;
  wire [13:0] _GEN_6116 = 14'h17e4 == index ? 14'h2f : _GEN_6115;
  wire [13:0] _GEN_6117 = 14'h17e5 == index ? 14'h2f : _GEN_6116;
  wire [13:0] _GEN_6118 = 14'h17e6 == index ? 14'h2f : _GEN_6117;
  wire [13:0] _GEN_6119 = 14'h17e7 == index ? 14'h2f : _GEN_6118;
  wire [13:0] _GEN_6120 = 14'h17e8 == index ? 14'h2f : _GEN_6119;
  wire [13:0] _GEN_6121 = 14'h17e9 == index ? 14'h2f : _GEN_6120;
  wire [13:0] _GEN_6122 = 14'h17ea == index ? 14'h2f : _GEN_6121;
  wire [13:0] _GEN_6123 = 14'h17eb == index ? 14'h2f : _GEN_6122;
  wire [13:0] _GEN_6124 = 14'h17ec == index ? 14'h2f : _GEN_6123;
  wire [13:0] _GEN_6125 = 14'h17ed == index ? 14'h2f : _GEN_6124;
  wire [13:0] _GEN_6126 = 14'h17ee == index ? 14'h2f : _GEN_6125;
  wire [13:0] _GEN_6127 = 14'h17ef == index ? 14'h2f : _GEN_6126;
  wire [13:0] _GEN_6128 = 14'h17f0 == index ? 14'h2f : _GEN_6127;
  wire [13:0] _GEN_6129 = 14'h17f1 == index ? 14'h2f : _GEN_6128;
  wire [13:0] _GEN_6130 = 14'h17f2 == index ? 14'h2f : _GEN_6129;
  wire [13:0] _GEN_6131 = 14'h17f3 == index ? 14'h2f : _GEN_6130;
  wire [13:0] _GEN_6132 = 14'h17f4 == index ? 14'h2f : _GEN_6131;
  wire [13:0] _GEN_6133 = 14'h17f5 == index ? 14'h2f : _GEN_6132;
  wire [13:0] _GEN_6134 = 14'h17f6 == index ? 14'h2f : _GEN_6133;
  wire [13:0] _GEN_6135 = 14'h17f7 == index ? 14'h2f : _GEN_6134;
  wire [13:0] _GEN_6136 = 14'h17f8 == index ? 14'h2f : _GEN_6135;
  wire [13:0] _GEN_6137 = 14'h17f9 == index ? 14'h2f : _GEN_6136;
  wire [13:0] _GEN_6138 = 14'h17fa == index ? 14'h2f : _GEN_6137;
  wire [13:0] _GEN_6139 = 14'h17fb == index ? 14'h2f : _GEN_6138;
  wire [13:0] _GEN_6140 = 14'h17fc == index ? 14'h2f : _GEN_6139;
  wire [13:0] _GEN_6141 = 14'h17fd == index ? 14'h2f : _GEN_6140;
  wire [13:0] _GEN_6142 = 14'h17fe == index ? 14'h2f : _GEN_6141;
  wire [13:0] _GEN_6143 = 14'h17ff == index ? 14'h2f : _GEN_6142;
  wire [13:0] _GEN_6144 = 14'h1800 == index ? 14'h0 : _GEN_6143;
  wire [13:0] _GEN_6145 = 14'h1801 == index ? 14'h1800 : _GEN_6144;
  wire [13:0] _GEN_6146 = 14'h1802 == index ? 14'hc00 : _GEN_6145;
  wire [13:0] _GEN_6147 = 14'h1803 == index ? 14'h800 : _GEN_6146;
  wire [13:0] _GEN_6148 = 14'h1804 == index ? 14'h600 : _GEN_6147;
  wire [13:0] _GEN_6149 = 14'h1805 == index ? 14'h483 : _GEN_6148;
  wire [13:0] _GEN_6150 = 14'h1806 == index ? 14'h400 : _GEN_6149;
  wire [13:0] _GEN_6151 = 14'h1807 == index ? 14'h306 : _GEN_6150;
  wire [13:0] _GEN_6152 = 14'h1808 == index ? 14'h300 : _GEN_6151;
  wire [13:0] _GEN_6153 = 14'h1809 == index ? 14'h283 : _GEN_6152;
  wire [13:0] _GEN_6154 = 14'h180a == index ? 14'h208 : _GEN_6153;
  wire [13:0] _GEN_6155 = 14'h180b == index ? 14'h204 : _GEN_6154;
  wire [13:0] _GEN_6156 = 14'h180c == index ? 14'h200 : _GEN_6155;
  wire [13:0] _GEN_6157 = 14'h180d == index ? 14'h189 : _GEN_6156;
  wire [13:0] _GEN_6158 = 14'h180e == index ? 14'h186 : _GEN_6157;
  wire [13:0] _GEN_6159 = 14'h180f == index ? 14'h183 : _GEN_6158;
  wire [13:0] _GEN_6160 = 14'h1810 == index ? 14'h180 : _GEN_6159;
  wire [13:0] _GEN_6161 = 14'h1811 == index ? 14'h10e : _GEN_6160;
  wire [13:0] _GEN_6162 = 14'h1812 == index ? 14'h10c : _GEN_6161;
  wire [13:0] _GEN_6163 = 14'h1813 == index ? 14'h10a : _GEN_6162;
  wire [13:0] _GEN_6164 = 14'h1814 == index ? 14'h108 : _GEN_6163;
  wire [13:0] _GEN_6165 = 14'h1815 == index ? 14'h106 : _GEN_6164;
  wire [13:0] _GEN_6166 = 14'h1816 == index ? 14'h104 : _GEN_6165;
  wire [13:0] _GEN_6167 = 14'h1817 == index ? 14'h102 : _GEN_6166;
  wire [13:0] _GEN_6168 = 14'h1818 == index ? 14'h100 : _GEN_6167;
  wire [13:0] _GEN_6169 = 14'h1819 == index ? 14'h97 : _GEN_6168;
  wire [13:0] _GEN_6170 = 14'h181a == index ? 14'h96 : _GEN_6169;
  wire [13:0] _GEN_6171 = 14'h181b == index ? 14'h95 : _GEN_6170;
  wire [13:0] _GEN_6172 = 14'h181c == index ? 14'h94 : _GEN_6171;
  wire [13:0] _GEN_6173 = 14'h181d == index ? 14'h93 : _GEN_6172;
  wire [13:0] _GEN_6174 = 14'h181e == index ? 14'h92 : _GEN_6173;
  wire [13:0] _GEN_6175 = 14'h181f == index ? 14'h91 : _GEN_6174;
  wire [13:0] _GEN_6176 = 14'h1820 == index ? 14'h90 : _GEN_6175;
  wire [13:0] _GEN_6177 = 14'h1821 == index ? 14'h8f : _GEN_6176;
  wire [13:0] _GEN_6178 = 14'h1822 == index ? 14'h8e : _GEN_6177;
  wire [13:0] _GEN_6179 = 14'h1823 == index ? 14'h8d : _GEN_6178;
  wire [13:0] _GEN_6180 = 14'h1824 == index ? 14'h8c : _GEN_6179;
  wire [13:0] _GEN_6181 = 14'h1825 == index ? 14'h8b : _GEN_6180;
  wire [13:0] _GEN_6182 = 14'h1826 == index ? 14'h8a : _GEN_6181;
  wire [13:0] _GEN_6183 = 14'h1827 == index ? 14'h89 : _GEN_6182;
  wire [13:0] _GEN_6184 = 14'h1828 == index ? 14'h88 : _GEN_6183;
  wire [13:0] _GEN_6185 = 14'h1829 == index ? 14'h87 : _GEN_6184;
  wire [13:0] _GEN_6186 = 14'h182a == index ? 14'h86 : _GEN_6185;
  wire [13:0] _GEN_6187 = 14'h182b == index ? 14'h85 : _GEN_6186;
  wire [13:0] _GEN_6188 = 14'h182c == index ? 14'h84 : _GEN_6187;
  wire [13:0] _GEN_6189 = 14'h182d == index ? 14'h83 : _GEN_6188;
  wire [13:0] _GEN_6190 = 14'h182e == index ? 14'h82 : _GEN_6189;
  wire [13:0] _GEN_6191 = 14'h182f == index ? 14'h81 : _GEN_6190;
  wire [13:0] _GEN_6192 = 14'h1830 == index ? 14'h80 : _GEN_6191;
  wire [13:0] _GEN_6193 = 14'h1831 == index ? 14'h30 : _GEN_6192;
  wire [13:0] _GEN_6194 = 14'h1832 == index ? 14'h30 : _GEN_6193;
  wire [13:0] _GEN_6195 = 14'h1833 == index ? 14'h30 : _GEN_6194;
  wire [13:0] _GEN_6196 = 14'h1834 == index ? 14'h30 : _GEN_6195;
  wire [13:0] _GEN_6197 = 14'h1835 == index ? 14'h30 : _GEN_6196;
  wire [13:0] _GEN_6198 = 14'h1836 == index ? 14'h30 : _GEN_6197;
  wire [13:0] _GEN_6199 = 14'h1837 == index ? 14'h30 : _GEN_6198;
  wire [13:0] _GEN_6200 = 14'h1838 == index ? 14'h30 : _GEN_6199;
  wire [13:0] _GEN_6201 = 14'h1839 == index ? 14'h30 : _GEN_6200;
  wire [13:0] _GEN_6202 = 14'h183a == index ? 14'h30 : _GEN_6201;
  wire [13:0] _GEN_6203 = 14'h183b == index ? 14'h30 : _GEN_6202;
  wire [13:0] _GEN_6204 = 14'h183c == index ? 14'h30 : _GEN_6203;
  wire [13:0] _GEN_6205 = 14'h183d == index ? 14'h30 : _GEN_6204;
  wire [13:0] _GEN_6206 = 14'h183e == index ? 14'h30 : _GEN_6205;
  wire [13:0] _GEN_6207 = 14'h183f == index ? 14'h30 : _GEN_6206;
  wire [13:0] _GEN_6208 = 14'h1840 == index ? 14'h30 : _GEN_6207;
  wire [13:0] _GEN_6209 = 14'h1841 == index ? 14'h30 : _GEN_6208;
  wire [13:0] _GEN_6210 = 14'h1842 == index ? 14'h30 : _GEN_6209;
  wire [13:0] _GEN_6211 = 14'h1843 == index ? 14'h30 : _GEN_6210;
  wire [13:0] _GEN_6212 = 14'h1844 == index ? 14'h30 : _GEN_6211;
  wire [13:0] _GEN_6213 = 14'h1845 == index ? 14'h30 : _GEN_6212;
  wire [13:0] _GEN_6214 = 14'h1846 == index ? 14'h30 : _GEN_6213;
  wire [13:0] _GEN_6215 = 14'h1847 == index ? 14'h30 : _GEN_6214;
  wire [13:0] _GEN_6216 = 14'h1848 == index ? 14'h30 : _GEN_6215;
  wire [13:0] _GEN_6217 = 14'h1849 == index ? 14'h30 : _GEN_6216;
  wire [13:0] _GEN_6218 = 14'h184a == index ? 14'h30 : _GEN_6217;
  wire [13:0] _GEN_6219 = 14'h184b == index ? 14'h30 : _GEN_6218;
  wire [13:0] _GEN_6220 = 14'h184c == index ? 14'h30 : _GEN_6219;
  wire [13:0] _GEN_6221 = 14'h184d == index ? 14'h30 : _GEN_6220;
  wire [13:0] _GEN_6222 = 14'h184e == index ? 14'h30 : _GEN_6221;
  wire [13:0] _GEN_6223 = 14'h184f == index ? 14'h30 : _GEN_6222;
  wire [13:0] _GEN_6224 = 14'h1850 == index ? 14'h30 : _GEN_6223;
  wire [13:0] _GEN_6225 = 14'h1851 == index ? 14'h30 : _GEN_6224;
  wire [13:0] _GEN_6226 = 14'h1852 == index ? 14'h30 : _GEN_6225;
  wire [13:0] _GEN_6227 = 14'h1853 == index ? 14'h30 : _GEN_6226;
  wire [13:0] _GEN_6228 = 14'h1854 == index ? 14'h30 : _GEN_6227;
  wire [13:0] _GEN_6229 = 14'h1855 == index ? 14'h30 : _GEN_6228;
  wire [13:0] _GEN_6230 = 14'h1856 == index ? 14'h30 : _GEN_6229;
  wire [13:0] _GEN_6231 = 14'h1857 == index ? 14'h30 : _GEN_6230;
  wire [13:0] _GEN_6232 = 14'h1858 == index ? 14'h30 : _GEN_6231;
  wire [13:0] _GEN_6233 = 14'h1859 == index ? 14'h30 : _GEN_6232;
  wire [13:0] _GEN_6234 = 14'h185a == index ? 14'h30 : _GEN_6233;
  wire [13:0] _GEN_6235 = 14'h185b == index ? 14'h30 : _GEN_6234;
  wire [13:0] _GEN_6236 = 14'h185c == index ? 14'h30 : _GEN_6235;
  wire [13:0] _GEN_6237 = 14'h185d == index ? 14'h30 : _GEN_6236;
  wire [13:0] _GEN_6238 = 14'h185e == index ? 14'h30 : _GEN_6237;
  wire [13:0] _GEN_6239 = 14'h185f == index ? 14'h30 : _GEN_6238;
  wire [13:0] _GEN_6240 = 14'h1860 == index ? 14'h30 : _GEN_6239;
  wire [13:0] _GEN_6241 = 14'h1861 == index ? 14'h30 : _GEN_6240;
  wire [13:0] _GEN_6242 = 14'h1862 == index ? 14'h30 : _GEN_6241;
  wire [13:0] _GEN_6243 = 14'h1863 == index ? 14'h30 : _GEN_6242;
  wire [13:0] _GEN_6244 = 14'h1864 == index ? 14'h30 : _GEN_6243;
  wire [13:0] _GEN_6245 = 14'h1865 == index ? 14'h30 : _GEN_6244;
  wire [13:0] _GEN_6246 = 14'h1866 == index ? 14'h30 : _GEN_6245;
  wire [13:0] _GEN_6247 = 14'h1867 == index ? 14'h30 : _GEN_6246;
  wire [13:0] _GEN_6248 = 14'h1868 == index ? 14'h30 : _GEN_6247;
  wire [13:0] _GEN_6249 = 14'h1869 == index ? 14'h30 : _GEN_6248;
  wire [13:0] _GEN_6250 = 14'h186a == index ? 14'h30 : _GEN_6249;
  wire [13:0] _GEN_6251 = 14'h186b == index ? 14'h30 : _GEN_6250;
  wire [13:0] _GEN_6252 = 14'h186c == index ? 14'h30 : _GEN_6251;
  wire [13:0] _GEN_6253 = 14'h186d == index ? 14'h30 : _GEN_6252;
  wire [13:0] _GEN_6254 = 14'h186e == index ? 14'h30 : _GEN_6253;
  wire [13:0] _GEN_6255 = 14'h186f == index ? 14'h30 : _GEN_6254;
  wire [13:0] _GEN_6256 = 14'h1870 == index ? 14'h30 : _GEN_6255;
  wire [13:0] _GEN_6257 = 14'h1871 == index ? 14'h30 : _GEN_6256;
  wire [13:0] _GEN_6258 = 14'h1872 == index ? 14'h30 : _GEN_6257;
  wire [13:0] _GEN_6259 = 14'h1873 == index ? 14'h30 : _GEN_6258;
  wire [13:0] _GEN_6260 = 14'h1874 == index ? 14'h30 : _GEN_6259;
  wire [13:0] _GEN_6261 = 14'h1875 == index ? 14'h30 : _GEN_6260;
  wire [13:0] _GEN_6262 = 14'h1876 == index ? 14'h30 : _GEN_6261;
  wire [13:0] _GEN_6263 = 14'h1877 == index ? 14'h30 : _GEN_6262;
  wire [13:0] _GEN_6264 = 14'h1878 == index ? 14'h30 : _GEN_6263;
  wire [13:0] _GEN_6265 = 14'h1879 == index ? 14'h30 : _GEN_6264;
  wire [13:0] _GEN_6266 = 14'h187a == index ? 14'h30 : _GEN_6265;
  wire [13:0] _GEN_6267 = 14'h187b == index ? 14'h30 : _GEN_6266;
  wire [13:0] _GEN_6268 = 14'h187c == index ? 14'h30 : _GEN_6267;
  wire [13:0] _GEN_6269 = 14'h187d == index ? 14'h30 : _GEN_6268;
  wire [13:0] _GEN_6270 = 14'h187e == index ? 14'h30 : _GEN_6269;
  wire [13:0] _GEN_6271 = 14'h187f == index ? 14'h30 : _GEN_6270;
  wire [13:0] _GEN_6272 = 14'h1880 == index ? 14'h0 : _GEN_6271;
  wire [13:0] _GEN_6273 = 14'h1881 == index ? 14'h1880 : _GEN_6272;
  wire [13:0] _GEN_6274 = 14'h1882 == index ? 14'hc01 : _GEN_6273;
  wire [13:0] _GEN_6275 = 14'h1883 == index ? 14'h801 : _GEN_6274;
  wire [13:0] _GEN_6276 = 14'h1884 == index ? 14'h601 : _GEN_6275;
  wire [13:0] _GEN_6277 = 14'h1885 == index ? 14'h484 : _GEN_6276;
  wire [13:0] _GEN_6278 = 14'h1886 == index ? 14'h401 : _GEN_6277;
  wire [13:0] _GEN_6279 = 14'h1887 == index ? 14'h380 : _GEN_6278;
  wire [13:0] _GEN_6280 = 14'h1888 == index ? 14'h301 : _GEN_6279;
  wire [13:0] _GEN_6281 = 14'h1889 == index ? 14'h284 : _GEN_6280;
  wire [13:0] _GEN_6282 = 14'h188a == index ? 14'h209 : _GEN_6281;
  wire [13:0] _GEN_6283 = 14'h188b == index ? 14'h205 : _GEN_6282;
  wire [13:0] _GEN_6284 = 14'h188c == index ? 14'h201 : _GEN_6283;
  wire [13:0] _GEN_6285 = 14'h188d == index ? 14'h18a : _GEN_6284;
  wire [13:0] _GEN_6286 = 14'h188e == index ? 14'h187 : _GEN_6285;
  wire [13:0] _GEN_6287 = 14'h188f == index ? 14'h184 : _GEN_6286;
  wire [13:0] _GEN_6288 = 14'h1890 == index ? 14'h181 : _GEN_6287;
  wire [13:0] _GEN_6289 = 14'h1891 == index ? 14'h10f : _GEN_6288;
  wire [13:0] _GEN_6290 = 14'h1892 == index ? 14'h10d : _GEN_6289;
  wire [13:0] _GEN_6291 = 14'h1893 == index ? 14'h10b : _GEN_6290;
  wire [13:0] _GEN_6292 = 14'h1894 == index ? 14'h109 : _GEN_6291;
  wire [13:0] _GEN_6293 = 14'h1895 == index ? 14'h107 : _GEN_6292;
  wire [13:0] _GEN_6294 = 14'h1896 == index ? 14'h105 : _GEN_6293;
  wire [13:0] _GEN_6295 = 14'h1897 == index ? 14'h103 : _GEN_6294;
  wire [13:0] _GEN_6296 = 14'h1898 == index ? 14'h101 : _GEN_6295;
  wire [13:0] _GEN_6297 = 14'h1899 == index ? 14'h98 : _GEN_6296;
  wire [13:0] _GEN_6298 = 14'h189a == index ? 14'h97 : _GEN_6297;
  wire [13:0] _GEN_6299 = 14'h189b == index ? 14'h96 : _GEN_6298;
  wire [13:0] _GEN_6300 = 14'h189c == index ? 14'h95 : _GEN_6299;
  wire [13:0] _GEN_6301 = 14'h189d == index ? 14'h94 : _GEN_6300;
  wire [13:0] _GEN_6302 = 14'h189e == index ? 14'h93 : _GEN_6301;
  wire [13:0] _GEN_6303 = 14'h189f == index ? 14'h92 : _GEN_6302;
  wire [13:0] _GEN_6304 = 14'h18a0 == index ? 14'h91 : _GEN_6303;
  wire [13:0] _GEN_6305 = 14'h18a1 == index ? 14'h90 : _GEN_6304;
  wire [13:0] _GEN_6306 = 14'h18a2 == index ? 14'h8f : _GEN_6305;
  wire [13:0] _GEN_6307 = 14'h18a3 == index ? 14'h8e : _GEN_6306;
  wire [13:0] _GEN_6308 = 14'h18a4 == index ? 14'h8d : _GEN_6307;
  wire [13:0] _GEN_6309 = 14'h18a5 == index ? 14'h8c : _GEN_6308;
  wire [13:0] _GEN_6310 = 14'h18a6 == index ? 14'h8b : _GEN_6309;
  wire [13:0] _GEN_6311 = 14'h18a7 == index ? 14'h8a : _GEN_6310;
  wire [13:0] _GEN_6312 = 14'h18a8 == index ? 14'h89 : _GEN_6311;
  wire [13:0] _GEN_6313 = 14'h18a9 == index ? 14'h88 : _GEN_6312;
  wire [13:0] _GEN_6314 = 14'h18aa == index ? 14'h87 : _GEN_6313;
  wire [13:0] _GEN_6315 = 14'h18ab == index ? 14'h86 : _GEN_6314;
  wire [13:0] _GEN_6316 = 14'h18ac == index ? 14'h85 : _GEN_6315;
  wire [13:0] _GEN_6317 = 14'h18ad == index ? 14'h84 : _GEN_6316;
  wire [13:0] _GEN_6318 = 14'h18ae == index ? 14'h83 : _GEN_6317;
  wire [13:0] _GEN_6319 = 14'h18af == index ? 14'h82 : _GEN_6318;
  wire [13:0] _GEN_6320 = 14'h18b0 == index ? 14'h81 : _GEN_6319;
  wire [13:0] _GEN_6321 = 14'h18b1 == index ? 14'h80 : _GEN_6320;
  wire [13:0] _GEN_6322 = 14'h18b2 == index ? 14'h31 : _GEN_6321;
  wire [13:0] _GEN_6323 = 14'h18b3 == index ? 14'h31 : _GEN_6322;
  wire [13:0] _GEN_6324 = 14'h18b4 == index ? 14'h31 : _GEN_6323;
  wire [13:0] _GEN_6325 = 14'h18b5 == index ? 14'h31 : _GEN_6324;
  wire [13:0] _GEN_6326 = 14'h18b6 == index ? 14'h31 : _GEN_6325;
  wire [13:0] _GEN_6327 = 14'h18b7 == index ? 14'h31 : _GEN_6326;
  wire [13:0] _GEN_6328 = 14'h18b8 == index ? 14'h31 : _GEN_6327;
  wire [13:0] _GEN_6329 = 14'h18b9 == index ? 14'h31 : _GEN_6328;
  wire [13:0] _GEN_6330 = 14'h18ba == index ? 14'h31 : _GEN_6329;
  wire [13:0] _GEN_6331 = 14'h18bb == index ? 14'h31 : _GEN_6330;
  wire [13:0] _GEN_6332 = 14'h18bc == index ? 14'h31 : _GEN_6331;
  wire [13:0] _GEN_6333 = 14'h18bd == index ? 14'h31 : _GEN_6332;
  wire [13:0] _GEN_6334 = 14'h18be == index ? 14'h31 : _GEN_6333;
  wire [13:0] _GEN_6335 = 14'h18bf == index ? 14'h31 : _GEN_6334;
  wire [13:0] _GEN_6336 = 14'h18c0 == index ? 14'h31 : _GEN_6335;
  wire [13:0] _GEN_6337 = 14'h18c1 == index ? 14'h31 : _GEN_6336;
  wire [13:0] _GEN_6338 = 14'h18c2 == index ? 14'h31 : _GEN_6337;
  wire [13:0] _GEN_6339 = 14'h18c3 == index ? 14'h31 : _GEN_6338;
  wire [13:0] _GEN_6340 = 14'h18c4 == index ? 14'h31 : _GEN_6339;
  wire [13:0] _GEN_6341 = 14'h18c5 == index ? 14'h31 : _GEN_6340;
  wire [13:0] _GEN_6342 = 14'h18c6 == index ? 14'h31 : _GEN_6341;
  wire [13:0] _GEN_6343 = 14'h18c7 == index ? 14'h31 : _GEN_6342;
  wire [13:0] _GEN_6344 = 14'h18c8 == index ? 14'h31 : _GEN_6343;
  wire [13:0] _GEN_6345 = 14'h18c9 == index ? 14'h31 : _GEN_6344;
  wire [13:0] _GEN_6346 = 14'h18ca == index ? 14'h31 : _GEN_6345;
  wire [13:0] _GEN_6347 = 14'h18cb == index ? 14'h31 : _GEN_6346;
  wire [13:0] _GEN_6348 = 14'h18cc == index ? 14'h31 : _GEN_6347;
  wire [13:0] _GEN_6349 = 14'h18cd == index ? 14'h31 : _GEN_6348;
  wire [13:0] _GEN_6350 = 14'h18ce == index ? 14'h31 : _GEN_6349;
  wire [13:0] _GEN_6351 = 14'h18cf == index ? 14'h31 : _GEN_6350;
  wire [13:0] _GEN_6352 = 14'h18d0 == index ? 14'h31 : _GEN_6351;
  wire [13:0] _GEN_6353 = 14'h18d1 == index ? 14'h31 : _GEN_6352;
  wire [13:0] _GEN_6354 = 14'h18d2 == index ? 14'h31 : _GEN_6353;
  wire [13:0] _GEN_6355 = 14'h18d3 == index ? 14'h31 : _GEN_6354;
  wire [13:0] _GEN_6356 = 14'h18d4 == index ? 14'h31 : _GEN_6355;
  wire [13:0] _GEN_6357 = 14'h18d5 == index ? 14'h31 : _GEN_6356;
  wire [13:0] _GEN_6358 = 14'h18d6 == index ? 14'h31 : _GEN_6357;
  wire [13:0] _GEN_6359 = 14'h18d7 == index ? 14'h31 : _GEN_6358;
  wire [13:0] _GEN_6360 = 14'h18d8 == index ? 14'h31 : _GEN_6359;
  wire [13:0] _GEN_6361 = 14'h18d9 == index ? 14'h31 : _GEN_6360;
  wire [13:0] _GEN_6362 = 14'h18da == index ? 14'h31 : _GEN_6361;
  wire [13:0] _GEN_6363 = 14'h18db == index ? 14'h31 : _GEN_6362;
  wire [13:0] _GEN_6364 = 14'h18dc == index ? 14'h31 : _GEN_6363;
  wire [13:0] _GEN_6365 = 14'h18dd == index ? 14'h31 : _GEN_6364;
  wire [13:0] _GEN_6366 = 14'h18de == index ? 14'h31 : _GEN_6365;
  wire [13:0] _GEN_6367 = 14'h18df == index ? 14'h31 : _GEN_6366;
  wire [13:0] _GEN_6368 = 14'h18e0 == index ? 14'h31 : _GEN_6367;
  wire [13:0] _GEN_6369 = 14'h18e1 == index ? 14'h31 : _GEN_6368;
  wire [13:0] _GEN_6370 = 14'h18e2 == index ? 14'h31 : _GEN_6369;
  wire [13:0] _GEN_6371 = 14'h18e3 == index ? 14'h31 : _GEN_6370;
  wire [13:0] _GEN_6372 = 14'h18e4 == index ? 14'h31 : _GEN_6371;
  wire [13:0] _GEN_6373 = 14'h18e5 == index ? 14'h31 : _GEN_6372;
  wire [13:0] _GEN_6374 = 14'h18e6 == index ? 14'h31 : _GEN_6373;
  wire [13:0] _GEN_6375 = 14'h18e7 == index ? 14'h31 : _GEN_6374;
  wire [13:0] _GEN_6376 = 14'h18e8 == index ? 14'h31 : _GEN_6375;
  wire [13:0] _GEN_6377 = 14'h18e9 == index ? 14'h31 : _GEN_6376;
  wire [13:0] _GEN_6378 = 14'h18ea == index ? 14'h31 : _GEN_6377;
  wire [13:0] _GEN_6379 = 14'h18eb == index ? 14'h31 : _GEN_6378;
  wire [13:0] _GEN_6380 = 14'h18ec == index ? 14'h31 : _GEN_6379;
  wire [13:0] _GEN_6381 = 14'h18ed == index ? 14'h31 : _GEN_6380;
  wire [13:0] _GEN_6382 = 14'h18ee == index ? 14'h31 : _GEN_6381;
  wire [13:0] _GEN_6383 = 14'h18ef == index ? 14'h31 : _GEN_6382;
  wire [13:0] _GEN_6384 = 14'h18f0 == index ? 14'h31 : _GEN_6383;
  wire [13:0] _GEN_6385 = 14'h18f1 == index ? 14'h31 : _GEN_6384;
  wire [13:0] _GEN_6386 = 14'h18f2 == index ? 14'h31 : _GEN_6385;
  wire [13:0] _GEN_6387 = 14'h18f3 == index ? 14'h31 : _GEN_6386;
  wire [13:0] _GEN_6388 = 14'h18f4 == index ? 14'h31 : _GEN_6387;
  wire [13:0] _GEN_6389 = 14'h18f5 == index ? 14'h31 : _GEN_6388;
  wire [13:0] _GEN_6390 = 14'h18f6 == index ? 14'h31 : _GEN_6389;
  wire [13:0] _GEN_6391 = 14'h18f7 == index ? 14'h31 : _GEN_6390;
  wire [13:0] _GEN_6392 = 14'h18f8 == index ? 14'h31 : _GEN_6391;
  wire [13:0] _GEN_6393 = 14'h18f9 == index ? 14'h31 : _GEN_6392;
  wire [13:0] _GEN_6394 = 14'h18fa == index ? 14'h31 : _GEN_6393;
  wire [13:0] _GEN_6395 = 14'h18fb == index ? 14'h31 : _GEN_6394;
  wire [13:0] _GEN_6396 = 14'h18fc == index ? 14'h31 : _GEN_6395;
  wire [13:0] _GEN_6397 = 14'h18fd == index ? 14'h31 : _GEN_6396;
  wire [13:0] _GEN_6398 = 14'h18fe == index ? 14'h31 : _GEN_6397;
  wire [13:0] _GEN_6399 = 14'h18ff == index ? 14'h31 : _GEN_6398;
  wire [13:0] _GEN_6400 = 14'h1900 == index ? 14'h0 : _GEN_6399;
  wire [13:0] _GEN_6401 = 14'h1901 == index ? 14'h1900 : _GEN_6400;
  wire [13:0] _GEN_6402 = 14'h1902 == index ? 14'hc80 : _GEN_6401;
  wire [13:0] _GEN_6403 = 14'h1903 == index ? 14'h802 : _GEN_6402;
  wire [13:0] _GEN_6404 = 14'h1904 == index ? 14'h602 : _GEN_6403;
  wire [13:0] _GEN_6405 = 14'h1905 == index ? 14'h500 : _GEN_6404;
  wire [13:0] _GEN_6406 = 14'h1906 == index ? 14'h402 : _GEN_6405;
  wire [13:0] _GEN_6407 = 14'h1907 == index ? 14'h381 : _GEN_6406;
  wire [13:0] _GEN_6408 = 14'h1908 == index ? 14'h302 : _GEN_6407;
  wire [13:0] _GEN_6409 = 14'h1909 == index ? 14'h285 : _GEN_6408;
  wire [13:0] _GEN_6410 = 14'h190a == index ? 14'h280 : _GEN_6409;
  wire [13:0] _GEN_6411 = 14'h190b == index ? 14'h206 : _GEN_6410;
  wire [13:0] _GEN_6412 = 14'h190c == index ? 14'h202 : _GEN_6411;
  wire [13:0] _GEN_6413 = 14'h190d == index ? 14'h18b : _GEN_6412;
  wire [13:0] _GEN_6414 = 14'h190e == index ? 14'h188 : _GEN_6413;
  wire [13:0] _GEN_6415 = 14'h190f == index ? 14'h185 : _GEN_6414;
  wire [13:0] _GEN_6416 = 14'h1910 == index ? 14'h182 : _GEN_6415;
  wire [13:0] _GEN_6417 = 14'h1911 == index ? 14'h110 : _GEN_6416;
  wire [13:0] _GEN_6418 = 14'h1912 == index ? 14'h10e : _GEN_6417;
  wire [13:0] _GEN_6419 = 14'h1913 == index ? 14'h10c : _GEN_6418;
  wire [13:0] _GEN_6420 = 14'h1914 == index ? 14'h10a : _GEN_6419;
  wire [13:0] _GEN_6421 = 14'h1915 == index ? 14'h108 : _GEN_6420;
  wire [13:0] _GEN_6422 = 14'h1916 == index ? 14'h106 : _GEN_6421;
  wire [13:0] _GEN_6423 = 14'h1917 == index ? 14'h104 : _GEN_6422;
  wire [13:0] _GEN_6424 = 14'h1918 == index ? 14'h102 : _GEN_6423;
  wire [13:0] _GEN_6425 = 14'h1919 == index ? 14'h100 : _GEN_6424;
  wire [13:0] _GEN_6426 = 14'h191a == index ? 14'h98 : _GEN_6425;
  wire [13:0] _GEN_6427 = 14'h191b == index ? 14'h97 : _GEN_6426;
  wire [13:0] _GEN_6428 = 14'h191c == index ? 14'h96 : _GEN_6427;
  wire [13:0] _GEN_6429 = 14'h191d == index ? 14'h95 : _GEN_6428;
  wire [13:0] _GEN_6430 = 14'h191e == index ? 14'h94 : _GEN_6429;
  wire [13:0] _GEN_6431 = 14'h191f == index ? 14'h93 : _GEN_6430;
  wire [13:0] _GEN_6432 = 14'h1920 == index ? 14'h92 : _GEN_6431;
  wire [13:0] _GEN_6433 = 14'h1921 == index ? 14'h91 : _GEN_6432;
  wire [13:0] _GEN_6434 = 14'h1922 == index ? 14'h90 : _GEN_6433;
  wire [13:0] _GEN_6435 = 14'h1923 == index ? 14'h8f : _GEN_6434;
  wire [13:0] _GEN_6436 = 14'h1924 == index ? 14'h8e : _GEN_6435;
  wire [13:0] _GEN_6437 = 14'h1925 == index ? 14'h8d : _GEN_6436;
  wire [13:0] _GEN_6438 = 14'h1926 == index ? 14'h8c : _GEN_6437;
  wire [13:0] _GEN_6439 = 14'h1927 == index ? 14'h8b : _GEN_6438;
  wire [13:0] _GEN_6440 = 14'h1928 == index ? 14'h8a : _GEN_6439;
  wire [13:0] _GEN_6441 = 14'h1929 == index ? 14'h89 : _GEN_6440;
  wire [13:0] _GEN_6442 = 14'h192a == index ? 14'h88 : _GEN_6441;
  wire [13:0] _GEN_6443 = 14'h192b == index ? 14'h87 : _GEN_6442;
  wire [13:0] _GEN_6444 = 14'h192c == index ? 14'h86 : _GEN_6443;
  wire [13:0] _GEN_6445 = 14'h192d == index ? 14'h85 : _GEN_6444;
  wire [13:0] _GEN_6446 = 14'h192e == index ? 14'h84 : _GEN_6445;
  wire [13:0] _GEN_6447 = 14'h192f == index ? 14'h83 : _GEN_6446;
  wire [13:0] _GEN_6448 = 14'h1930 == index ? 14'h82 : _GEN_6447;
  wire [13:0] _GEN_6449 = 14'h1931 == index ? 14'h81 : _GEN_6448;
  wire [13:0] _GEN_6450 = 14'h1932 == index ? 14'h80 : _GEN_6449;
  wire [13:0] _GEN_6451 = 14'h1933 == index ? 14'h32 : _GEN_6450;
  wire [13:0] _GEN_6452 = 14'h1934 == index ? 14'h32 : _GEN_6451;
  wire [13:0] _GEN_6453 = 14'h1935 == index ? 14'h32 : _GEN_6452;
  wire [13:0] _GEN_6454 = 14'h1936 == index ? 14'h32 : _GEN_6453;
  wire [13:0] _GEN_6455 = 14'h1937 == index ? 14'h32 : _GEN_6454;
  wire [13:0] _GEN_6456 = 14'h1938 == index ? 14'h32 : _GEN_6455;
  wire [13:0] _GEN_6457 = 14'h1939 == index ? 14'h32 : _GEN_6456;
  wire [13:0] _GEN_6458 = 14'h193a == index ? 14'h32 : _GEN_6457;
  wire [13:0] _GEN_6459 = 14'h193b == index ? 14'h32 : _GEN_6458;
  wire [13:0] _GEN_6460 = 14'h193c == index ? 14'h32 : _GEN_6459;
  wire [13:0] _GEN_6461 = 14'h193d == index ? 14'h32 : _GEN_6460;
  wire [13:0] _GEN_6462 = 14'h193e == index ? 14'h32 : _GEN_6461;
  wire [13:0] _GEN_6463 = 14'h193f == index ? 14'h32 : _GEN_6462;
  wire [13:0] _GEN_6464 = 14'h1940 == index ? 14'h32 : _GEN_6463;
  wire [13:0] _GEN_6465 = 14'h1941 == index ? 14'h32 : _GEN_6464;
  wire [13:0] _GEN_6466 = 14'h1942 == index ? 14'h32 : _GEN_6465;
  wire [13:0] _GEN_6467 = 14'h1943 == index ? 14'h32 : _GEN_6466;
  wire [13:0] _GEN_6468 = 14'h1944 == index ? 14'h32 : _GEN_6467;
  wire [13:0] _GEN_6469 = 14'h1945 == index ? 14'h32 : _GEN_6468;
  wire [13:0] _GEN_6470 = 14'h1946 == index ? 14'h32 : _GEN_6469;
  wire [13:0] _GEN_6471 = 14'h1947 == index ? 14'h32 : _GEN_6470;
  wire [13:0] _GEN_6472 = 14'h1948 == index ? 14'h32 : _GEN_6471;
  wire [13:0] _GEN_6473 = 14'h1949 == index ? 14'h32 : _GEN_6472;
  wire [13:0] _GEN_6474 = 14'h194a == index ? 14'h32 : _GEN_6473;
  wire [13:0] _GEN_6475 = 14'h194b == index ? 14'h32 : _GEN_6474;
  wire [13:0] _GEN_6476 = 14'h194c == index ? 14'h32 : _GEN_6475;
  wire [13:0] _GEN_6477 = 14'h194d == index ? 14'h32 : _GEN_6476;
  wire [13:0] _GEN_6478 = 14'h194e == index ? 14'h32 : _GEN_6477;
  wire [13:0] _GEN_6479 = 14'h194f == index ? 14'h32 : _GEN_6478;
  wire [13:0] _GEN_6480 = 14'h1950 == index ? 14'h32 : _GEN_6479;
  wire [13:0] _GEN_6481 = 14'h1951 == index ? 14'h32 : _GEN_6480;
  wire [13:0] _GEN_6482 = 14'h1952 == index ? 14'h32 : _GEN_6481;
  wire [13:0] _GEN_6483 = 14'h1953 == index ? 14'h32 : _GEN_6482;
  wire [13:0] _GEN_6484 = 14'h1954 == index ? 14'h32 : _GEN_6483;
  wire [13:0] _GEN_6485 = 14'h1955 == index ? 14'h32 : _GEN_6484;
  wire [13:0] _GEN_6486 = 14'h1956 == index ? 14'h32 : _GEN_6485;
  wire [13:0] _GEN_6487 = 14'h1957 == index ? 14'h32 : _GEN_6486;
  wire [13:0] _GEN_6488 = 14'h1958 == index ? 14'h32 : _GEN_6487;
  wire [13:0] _GEN_6489 = 14'h1959 == index ? 14'h32 : _GEN_6488;
  wire [13:0] _GEN_6490 = 14'h195a == index ? 14'h32 : _GEN_6489;
  wire [13:0] _GEN_6491 = 14'h195b == index ? 14'h32 : _GEN_6490;
  wire [13:0] _GEN_6492 = 14'h195c == index ? 14'h32 : _GEN_6491;
  wire [13:0] _GEN_6493 = 14'h195d == index ? 14'h32 : _GEN_6492;
  wire [13:0] _GEN_6494 = 14'h195e == index ? 14'h32 : _GEN_6493;
  wire [13:0] _GEN_6495 = 14'h195f == index ? 14'h32 : _GEN_6494;
  wire [13:0] _GEN_6496 = 14'h1960 == index ? 14'h32 : _GEN_6495;
  wire [13:0] _GEN_6497 = 14'h1961 == index ? 14'h32 : _GEN_6496;
  wire [13:0] _GEN_6498 = 14'h1962 == index ? 14'h32 : _GEN_6497;
  wire [13:0] _GEN_6499 = 14'h1963 == index ? 14'h32 : _GEN_6498;
  wire [13:0] _GEN_6500 = 14'h1964 == index ? 14'h32 : _GEN_6499;
  wire [13:0] _GEN_6501 = 14'h1965 == index ? 14'h32 : _GEN_6500;
  wire [13:0] _GEN_6502 = 14'h1966 == index ? 14'h32 : _GEN_6501;
  wire [13:0] _GEN_6503 = 14'h1967 == index ? 14'h32 : _GEN_6502;
  wire [13:0] _GEN_6504 = 14'h1968 == index ? 14'h32 : _GEN_6503;
  wire [13:0] _GEN_6505 = 14'h1969 == index ? 14'h32 : _GEN_6504;
  wire [13:0] _GEN_6506 = 14'h196a == index ? 14'h32 : _GEN_6505;
  wire [13:0] _GEN_6507 = 14'h196b == index ? 14'h32 : _GEN_6506;
  wire [13:0] _GEN_6508 = 14'h196c == index ? 14'h32 : _GEN_6507;
  wire [13:0] _GEN_6509 = 14'h196d == index ? 14'h32 : _GEN_6508;
  wire [13:0] _GEN_6510 = 14'h196e == index ? 14'h32 : _GEN_6509;
  wire [13:0] _GEN_6511 = 14'h196f == index ? 14'h32 : _GEN_6510;
  wire [13:0] _GEN_6512 = 14'h1970 == index ? 14'h32 : _GEN_6511;
  wire [13:0] _GEN_6513 = 14'h1971 == index ? 14'h32 : _GEN_6512;
  wire [13:0] _GEN_6514 = 14'h1972 == index ? 14'h32 : _GEN_6513;
  wire [13:0] _GEN_6515 = 14'h1973 == index ? 14'h32 : _GEN_6514;
  wire [13:0] _GEN_6516 = 14'h1974 == index ? 14'h32 : _GEN_6515;
  wire [13:0] _GEN_6517 = 14'h1975 == index ? 14'h32 : _GEN_6516;
  wire [13:0] _GEN_6518 = 14'h1976 == index ? 14'h32 : _GEN_6517;
  wire [13:0] _GEN_6519 = 14'h1977 == index ? 14'h32 : _GEN_6518;
  wire [13:0] _GEN_6520 = 14'h1978 == index ? 14'h32 : _GEN_6519;
  wire [13:0] _GEN_6521 = 14'h1979 == index ? 14'h32 : _GEN_6520;
  wire [13:0] _GEN_6522 = 14'h197a == index ? 14'h32 : _GEN_6521;
  wire [13:0] _GEN_6523 = 14'h197b == index ? 14'h32 : _GEN_6522;
  wire [13:0] _GEN_6524 = 14'h197c == index ? 14'h32 : _GEN_6523;
  wire [13:0] _GEN_6525 = 14'h197d == index ? 14'h32 : _GEN_6524;
  wire [13:0] _GEN_6526 = 14'h197e == index ? 14'h32 : _GEN_6525;
  wire [13:0] _GEN_6527 = 14'h197f == index ? 14'h32 : _GEN_6526;
  wire [13:0] _GEN_6528 = 14'h1980 == index ? 14'h0 : _GEN_6527;
  wire [13:0] _GEN_6529 = 14'h1981 == index ? 14'h1980 : _GEN_6528;
  wire [13:0] _GEN_6530 = 14'h1982 == index ? 14'hc81 : _GEN_6529;
  wire [13:0] _GEN_6531 = 14'h1983 == index ? 14'h880 : _GEN_6530;
  wire [13:0] _GEN_6532 = 14'h1984 == index ? 14'h603 : _GEN_6531;
  wire [13:0] _GEN_6533 = 14'h1985 == index ? 14'h501 : _GEN_6532;
  wire [13:0] _GEN_6534 = 14'h1986 == index ? 14'h403 : _GEN_6533;
  wire [13:0] _GEN_6535 = 14'h1987 == index ? 14'h382 : _GEN_6534;
  wire [13:0] _GEN_6536 = 14'h1988 == index ? 14'h303 : _GEN_6535;
  wire [13:0] _GEN_6537 = 14'h1989 == index ? 14'h286 : _GEN_6536;
  wire [13:0] _GEN_6538 = 14'h198a == index ? 14'h281 : _GEN_6537;
  wire [13:0] _GEN_6539 = 14'h198b == index ? 14'h207 : _GEN_6538;
  wire [13:0] _GEN_6540 = 14'h198c == index ? 14'h203 : _GEN_6539;
  wire [13:0] _GEN_6541 = 14'h198d == index ? 14'h18c : _GEN_6540;
  wire [13:0] _GEN_6542 = 14'h198e == index ? 14'h189 : _GEN_6541;
  wire [13:0] _GEN_6543 = 14'h198f == index ? 14'h186 : _GEN_6542;
  wire [13:0] _GEN_6544 = 14'h1990 == index ? 14'h183 : _GEN_6543;
  wire [13:0] _GEN_6545 = 14'h1991 == index ? 14'h180 : _GEN_6544;
  wire [13:0] _GEN_6546 = 14'h1992 == index ? 14'h10f : _GEN_6545;
  wire [13:0] _GEN_6547 = 14'h1993 == index ? 14'h10d : _GEN_6546;
  wire [13:0] _GEN_6548 = 14'h1994 == index ? 14'h10b : _GEN_6547;
  wire [13:0] _GEN_6549 = 14'h1995 == index ? 14'h109 : _GEN_6548;
  wire [13:0] _GEN_6550 = 14'h1996 == index ? 14'h107 : _GEN_6549;
  wire [13:0] _GEN_6551 = 14'h1997 == index ? 14'h105 : _GEN_6550;
  wire [13:0] _GEN_6552 = 14'h1998 == index ? 14'h103 : _GEN_6551;
  wire [13:0] _GEN_6553 = 14'h1999 == index ? 14'h101 : _GEN_6552;
  wire [13:0] _GEN_6554 = 14'h199a == index ? 14'h99 : _GEN_6553;
  wire [13:0] _GEN_6555 = 14'h199b == index ? 14'h98 : _GEN_6554;
  wire [13:0] _GEN_6556 = 14'h199c == index ? 14'h97 : _GEN_6555;
  wire [13:0] _GEN_6557 = 14'h199d == index ? 14'h96 : _GEN_6556;
  wire [13:0] _GEN_6558 = 14'h199e == index ? 14'h95 : _GEN_6557;
  wire [13:0] _GEN_6559 = 14'h199f == index ? 14'h94 : _GEN_6558;
  wire [13:0] _GEN_6560 = 14'h19a0 == index ? 14'h93 : _GEN_6559;
  wire [13:0] _GEN_6561 = 14'h19a1 == index ? 14'h92 : _GEN_6560;
  wire [13:0] _GEN_6562 = 14'h19a2 == index ? 14'h91 : _GEN_6561;
  wire [13:0] _GEN_6563 = 14'h19a3 == index ? 14'h90 : _GEN_6562;
  wire [13:0] _GEN_6564 = 14'h19a4 == index ? 14'h8f : _GEN_6563;
  wire [13:0] _GEN_6565 = 14'h19a5 == index ? 14'h8e : _GEN_6564;
  wire [13:0] _GEN_6566 = 14'h19a6 == index ? 14'h8d : _GEN_6565;
  wire [13:0] _GEN_6567 = 14'h19a7 == index ? 14'h8c : _GEN_6566;
  wire [13:0] _GEN_6568 = 14'h19a8 == index ? 14'h8b : _GEN_6567;
  wire [13:0] _GEN_6569 = 14'h19a9 == index ? 14'h8a : _GEN_6568;
  wire [13:0] _GEN_6570 = 14'h19aa == index ? 14'h89 : _GEN_6569;
  wire [13:0] _GEN_6571 = 14'h19ab == index ? 14'h88 : _GEN_6570;
  wire [13:0] _GEN_6572 = 14'h19ac == index ? 14'h87 : _GEN_6571;
  wire [13:0] _GEN_6573 = 14'h19ad == index ? 14'h86 : _GEN_6572;
  wire [13:0] _GEN_6574 = 14'h19ae == index ? 14'h85 : _GEN_6573;
  wire [13:0] _GEN_6575 = 14'h19af == index ? 14'h84 : _GEN_6574;
  wire [13:0] _GEN_6576 = 14'h19b0 == index ? 14'h83 : _GEN_6575;
  wire [13:0] _GEN_6577 = 14'h19b1 == index ? 14'h82 : _GEN_6576;
  wire [13:0] _GEN_6578 = 14'h19b2 == index ? 14'h81 : _GEN_6577;
  wire [13:0] _GEN_6579 = 14'h19b3 == index ? 14'h80 : _GEN_6578;
  wire [13:0] _GEN_6580 = 14'h19b4 == index ? 14'h33 : _GEN_6579;
  wire [13:0] _GEN_6581 = 14'h19b5 == index ? 14'h33 : _GEN_6580;
  wire [13:0] _GEN_6582 = 14'h19b6 == index ? 14'h33 : _GEN_6581;
  wire [13:0] _GEN_6583 = 14'h19b7 == index ? 14'h33 : _GEN_6582;
  wire [13:0] _GEN_6584 = 14'h19b8 == index ? 14'h33 : _GEN_6583;
  wire [13:0] _GEN_6585 = 14'h19b9 == index ? 14'h33 : _GEN_6584;
  wire [13:0] _GEN_6586 = 14'h19ba == index ? 14'h33 : _GEN_6585;
  wire [13:0] _GEN_6587 = 14'h19bb == index ? 14'h33 : _GEN_6586;
  wire [13:0] _GEN_6588 = 14'h19bc == index ? 14'h33 : _GEN_6587;
  wire [13:0] _GEN_6589 = 14'h19bd == index ? 14'h33 : _GEN_6588;
  wire [13:0] _GEN_6590 = 14'h19be == index ? 14'h33 : _GEN_6589;
  wire [13:0] _GEN_6591 = 14'h19bf == index ? 14'h33 : _GEN_6590;
  wire [13:0] _GEN_6592 = 14'h19c0 == index ? 14'h33 : _GEN_6591;
  wire [13:0] _GEN_6593 = 14'h19c1 == index ? 14'h33 : _GEN_6592;
  wire [13:0] _GEN_6594 = 14'h19c2 == index ? 14'h33 : _GEN_6593;
  wire [13:0] _GEN_6595 = 14'h19c3 == index ? 14'h33 : _GEN_6594;
  wire [13:0] _GEN_6596 = 14'h19c4 == index ? 14'h33 : _GEN_6595;
  wire [13:0] _GEN_6597 = 14'h19c5 == index ? 14'h33 : _GEN_6596;
  wire [13:0] _GEN_6598 = 14'h19c6 == index ? 14'h33 : _GEN_6597;
  wire [13:0] _GEN_6599 = 14'h19c7 == index ? 14'h33 : _GEN_6598;
  wire [13:0] _GEN_6600 = 14'h19c8 == index ? 14'h33 : _GEN_6599;
  wire [13:0] _GEN_6601 = 14'h19c9 == index ? 14'h33 : _GEN_6600;
  wire [13:0] _GEN_6602 = 14'h19ca == index ? 14'h33 : _GEN_6601;
  wire [13:0] _GEN_6603 = 14'h19cb == index ? 14'h33 : _GEN_6602;
  wire [13:0] _GEN_6604 = 14'h19cc == index ? 14'h33 : _GEN_6603;
  wire [13:0] _GEN_6605 = 14'h19cd == index ? 14'h33 : _GEN_6604;
  wire [13:0] _GEN_6606 = 14'h19ce == index ? 14'h33 : _GEN_6605;
  wire [13:0] _GEN_6607 = 14'h19cf == index ? 14'h33 : _GEN_6606;
  wire [13:0] _GEN_6608 = 14'h19d0 == index ? 14'h33 : _GEN_6607;
  wire [13:0] _GEN_6609 = 14'h19d1 == index ? 14'h33 : _GEN_6608;
  wire [13:0] _GEN_6610 = 14'h19d2 == index ? 14'h33 : _GEN_6609;
  wire [13:0] _GEN_6611 = 14'h19d3 == index ? 14'h33 : _GEN_6610;
  wire [13:0] _GEN_6612 = 14'h19d4 == index ? 14'h33 : _GEN_6611;
  wire [13:0] _GEN_6613 = 14'h19d5 == index ? 14'h33 : _GEN_6612;
  wire [13:0] _GEN_6614 = 14'h19d6 == index ? 14'h33 : _GEN_6613;
  wire [13:0] _GEN_6615 = 14'h19d7 == index ? 14'h33 : _GEN_6614;
  wire [13:0] _GEN_6616 = 14'h19d8 == index ? 14'h33 : _GEN_6615;
  wire [13:0] _GEN_6617 = 14'h19d9 == index ? 14'h33 : _GEN_6616;
  wire [13:0] _GEN_6618 = 14'h19da == index ? 14'h33 : _GEN_6617;
  wire [13:0] _GEN_6619 = 14'h19db == index ? 14'h33 : _GEN_6618;
  wire [13:0] _GEN_6620 = 14'h19dc == index ? 14'h33 : _GEN_6619;
  wire [13:0] _GEN_6621 = 14'h19dd == index ? 14'h33 : _GEN_6620;
  wire [13:0] _GEN_6622 = 14'h19de == index ? 14'h33 : _GEN_6621;
  wire [13:0] _GEN_6623 = 14'h19df == index ? 14'h33 : _GEN_6622;
  wire [13:0] _GEN_6624 = 14'h19e0 == index ? 14'h33 : _GEN_6623;
  wire [13:0] _GEN_6625 = 14'h19e1 == index ? 14'h33 : _GEN_6624;
  wire [13:0] _GEN_6626 = 14'h19e2 == index ? 14'h33 : _GEN_6625;
  wire [13:0] _GEN_6627 = 14'h19e3 == index ? 14'h33 : _GEN_6626;
  wire [13:0] _GEN_6628 = 14'h19e4 == index ? 14'h33 : _GEN_6627;
  wire [13:0] _GEN_6629 = 14'h19e5 == index ? 14'h33 : _GEN_6628;
  wire [13:0] _GEN_6630 = 14'h19e6 == index ? 14'h33 : _GEN_6629;
  wire [13:0] _GEN_6631 = 14'h19e7 == index ? 14'h33 : _GEN_6630;
  wire [13:0] _GEN_6632 = 14'h19e8 == index ? 14'h33 : _GEN_6631;
  wire [13:0] _GEN_6633 = 14'h19e9 == index ? 14'h33 : _GEN_6632;
  wire [13:0] _GEN_6634 = 14'h19ea == index ? 14'h33 : _GEN_6633;
  wire [13:0] _GEN_6635 = 14'h19eb == index ? 14'h33 : _GEN_6634;
  wire [13:0] _GEN_6636 = 14'h19ec == index ? 14'h33 : _GEN_6635;
  wire [13:0] _GEN_6637 = 14'h19ed == index ? 14'h33 : _GEN_6636;
  wire [13:0] _GEN_6638 = 14'h19ee == index ? 14'h33 : _GEN_6637;
  wire [13:0] _GEN_6639 = 14'h19ef == index ? 14'h33 : _GEN_6638;
  wire [13:0] _GEN_6640 = 14'h19f0 == index ? 14'h33 : _GEN_6639;
  wire [13:0] _GEN_6641 = 14'h19f1 == index ? 14'h33 : _GEN_6640;
  wire [13:0] _GEN_6642 = 14'h19f2 == index ? 14'h33 : _GEN_6641;
  wire [13:0] _GEN_6643 = 14'h19f3 == index ? 14'h33 : _GEN_6642;
  wire [13:0] _GEN_6644 = 14'h19f4 == index ? 14'h33 : _GEN_6643;
  wire [13:0] _GEN_6645 = 14'h19f5 == index ? 14'h33 : _GEN_6644;
  wire [13:0] _GEN_6646 = 14'h19f6 == index ? 14'h33 : _GEN_6645;
  wire [13:0] _GEN_6647 = 14'h19f7 == index ? 14'h33 : _GEN_6646;
  wire [13:0] _GEN_6648 = 14'h19f8 == index ? 14'h33 : _GEN_6647;
  wire [13:0] _GEN_6649 = 14'h19f9 == index ? 14'h33 : _GEN_6648;
  wire [13:0] _GEN_6650 = 14'h19fa == index ? 14'h33 : _GEN_6649;
  wire [13:0] _GEN_6651 = 14'h19fb == index ? 14'h33 : _GEN_6650;
  wire [13:0] _GEN_6652 = 14'h19fc == index ? 14'h33 : _GEN_6651;
  wire [13:0] _GEN_6653 = 14'h19fd == index ? 14'h33 : _GEN_6652;
  wire [13:0] _GEN_6654 = 14'h19fe == index ? 14'h33 : _GEN_6653;
  wire [13:0] _GEN_6655 = 14'h19ff == index ? 14'h33 : _GEN_6654;
  wire [13:0] _GEN_6656 = 14'h1a00 == index ? 14'h0 : _GEN_6655;
  wire [13:0] _GEN_6657 = 14'h1a01 == index ? 14'h1a00 : _GEN_6656;
  wire [13:0] _GEN_6658 = 14'h1a02 == index ? 14'hd00 : _GEN_6657;
  wire [13:0] _GEN_6659 = 14'h1a03 == index ? 14'h881 : _GEN_6658;
  wire [13:0] _GEN_6660 = 14'h1a04 == index ? 14'h680 : _GEN_6659;
  wire [13:0] _GEN_6661 = 14'h1a05 == index ? 14'h502 : _GEN_6660;
  wire [13:0] _GEN_6662 = 14'h1a06 == index ? 14'h404 : _GEN_6661;
  wire [13:0] _GEN_6663 = 14'h1a07 == index ? 14'h383 : _GEN_6662;
  wire [13:0] _GEN_6664 = 14'h1a08 == index ? 14'h304 : _GEN_6663;
  wire [13:0] _GEN_6665 = 14'h1a09 == index ? 14'h287 : _GEN_6664;
  wire [13:0] _GEN_6666 = 14'h1a0a == index ? 14'h282 : _GEN_6665;
  wire [13:0] _GEN_6667 = 14'h1a0b == index ? 14'h208 : _GEN_6666;
  wire [13:0] _GEN_6668 = 14'h1a0c == index ? 14'h204 : _GEN_6667;
  wire [13:0] _GEN_6669 = 14'h1a0d == index ? 14'h200 : _GEN_6668;
  wire [13:0] _GEN_6670 = 14'h1a0e == index ? 14'h18a : _GEN_6669;
  wire [13:0] _GEN_6671 = 14'h1a0f == index ? 14'h187 : _GEN_6670;
  wire [13:0] _GEN_6672 = 14'h1a10 == index ? 14'h184 : _GEN_6671;
  wire [13:0] _GEN_6673 = 14'h1a11 == index ? 14'h181 : _GEN_6672;
  wire [13:0] _GEN_6674 = 14'h1a12 == index ? 14'h110 : _GEN_6673;
  wire [13:0] _GEN_6675 = 14'h1a13 == index ? 14'h10e : _GEN_6674;
  wire [13:0] _GEN_6676 = 14'h1a14 == index ? 14'h10c : _GEN_6675;
  wire [13:0] _GEN_6677 = 14'h1a15 == index ? 14'h10a : _GEN_6676;
  wire [13:0] _GEN_6678 = 14'h1a16 == index ? 14'h108 : _GEN_6677;
  wire [13:0] _GEN_6679 = 14'h1a17 == index ? 14'h106 : _GEN_6678;
  wire [13:0] _GEN_6680 = 14'h1a18 == index ? 14'h104 : _GEN_6679;
  wire [13:0] _GEN_6681 = 14'h1a19 == index ? 14'h102 : _GEN_6680;
  wire [13:0] _GEN_6682 = 14'h1a1a == index ? 14'h100 : _GEN_6681;
  wire [13:0] _GEN_6683 = 14'h1a1b == index ? 14'h99 : _GEN_6682;
  wire [13:0] _GEN_6684 = 14'h1a1c == index ? 14'h98 : _GEN_6683;
  wire [13:0] _GEN_6685 = 14'h1a1d == index ? 14'h97 : _GEN_6684;
  wire [13:0] _GEN_6686 = 14'h1a1e == index ? 14'h96 : _GEN_6685;
  wire [13:0] _GEN_6687 = 14'h1a1f == index ? 14'h95 : _GEN_6686;
  wire [13:0] _GEN_6688 = 14'h1a20 == index ? 14'h94 : _GEN_6687;
  wire [13:0] _GEN_6689 = 14'h1a21 == index ? 14'h93 : _GEN_6688;
  wire [13:0] _GEN_6690 = 14'h1a22 == index ? 14'h92 : _GEN_6689;
  wire [13:0] _GEN_6691 = 14'h1a23 == index ? 14'h91 : _GEN_6690;
  wire [13:0] _GEN_6692 = 14'h1a24 == index ? 14'h90 : _GEN_6691;
  wire [13:0] _GEN_6693 = 14'h1a25 == index ? 14'h8f : _GEN_6692;
  wire [13:0] _GEN_6694 = 14'h1a26 == index ? 14'h8e : _GEN_6693;
  wire [13:0] _GEN_6695 = 14'h1a27 == index ? 14'h8d : _GEN_6694;
  wire [13:0] _GEN_6696 = 14'h1a28 == index ? 14'h8c : _GEN_6695;
  wire [13:0] _GEN_6697 = 14'h1a29 == index ? 14'h8b : _GEN_6696;
  wire [13:0] _GEN_6698 = 14'h1a2a == index ? 14'h8a : _GEN_6697;
  wire [13:0] _GEN_6699 = 14'h1a2b == index ? 14'h89 : _GEN_6698;
  wire [13:0] _GEN_6700 = 14'h1a2c == index ? 14'h88 : _GEN_6699;
  wire [13:0] _GEN_6701 = 14'h1a2d == index ? 14'h87 : _GEN_6700;
  wire [13:0] _GEN_6702 = 14'h1a2e == index ? 14'h86 : _GEN_6701;
  wire [13:0] _GEN_6703 = 14'h1a2f == index ? 14'h85 : _GEN_6702;
  wire [13:0] _GEN_6704 = 14'h1a30 == index ? 14'h84 : _GEN_6703;
  wire [13:0] _GEN_6705 = 14'h1a31 == index ? 14'h83 : _GEN_6704;
  wire [13:0] _GEN_6706 = 14'h1a32 == index ? 14'h82 : _GEN_6705;
  wire [13:0] _GEN_6707 = 14'h1a33 == index ? 14'h81 : _GEN_6706;
  wire [13:0] _GEN_6708 = 14'h1a34 == index ? 14'h80 : _GEN_6707;
  wire [13:0] _GEN_6709 = 14'h1a35 == index ? 14'h34 : _GEN_6708;
  wire [13:0] _GEN_6710 = 14'h1a36 == index ? 14'h34 : _GEN_6709;
  wire [13:0] _GEN_6711 = 14'h1a37 == index ? 14'h34 : _GEN_6710;
  wire [13:0] _GEN_6712 = 14'h1a38 == index ? 14'h34 : _GEN_6711;
  wire [13:0] _GEN_6713 = 14'h1a39 == index ? 14'h34 : _GEN_6712;
  wire [13:0] _GEN_6714 = 14'h1a3a == index ? 14'h34 : _GEN_6713;
  wire [13:0] _GEN_6715 = 14'h1a3b == index ? 14'h34 : _GEN_6714;
  wire [13:0] _GEN_6716 = 14'h1a3c == index ? 14'h34 : _GEN_6715;
  wire [13:0] _GEN_6717 = 14'h1a3d == index ? 14'h34 : _GEN_6716;
  wire [13:0] _GEN_6718 = 14'h1a3e == index ? 14'h34 : _GEN_6717;
  wire [13:0] _GEN_6719 = 14'h1a3f == index ? 14'h34 : _GEN_6718;
  wire [13:0] _GEN_6720 = 14'h1a40 == index ? 14'h34 : _GEN_6719;
  wire [13:0] _GEN_6721 = 14'h1a41 == index ? 14'h34 : _GEN_6720;
  wire [13:0] _GEN_6722 = 14'h1a42 == index ? 14'h34 : _GEN_6721;
  wire [13:0] _GEN_6723 = 14'h1a43 == index ? 14'h34 : _GEN_6722;
  wire [13:0] _GEN_6724 = 14'h1a44 == index ? 14'h34 : _GEN_6723;
  wire [13:0] _GEN_6725 = 14'h1a45 == index ? 14'h34 : _GEN_6724;
  wire [13:0] _GEN_6726 = 14'h1a46 == index ? 14'h34 : _GEN_6725;
  wire [13:0] _GEN_6727 = 14'h1a47 == index ? 14'h34 : _GEN_6726;
  wire [13:0] _GEN_6728 = 14'h1a48 == index ? 14'h34 : _GEN_6727;
  wire [13:0] _GEN_6729 = 14'h1a49 == index ? 14'h34 : _GEN_6728;
  wire [13:0] _GEN_6730 = 14'h1a4a == index ? 14'h34 : _GEN_6729;
  wire [13:0] _GEN_6731 = 14'h1a4b == index ? 14'h34 : _GEN_6730;
  wire [13:0] _GEN_6732 = 14'h1a4c == index ? 14'h34 : _GEN_6731;
  wire [13:0] _GEN_6733 = 14'h1a4d == index ? 14'h34 : _GEN_6732;
  wire [13:0] _GEN_6734 = 14'h1a4e == index ? 14'h34 : _GEN_6733;
  wire [13:0] _GEN_6735 = 14'h1a4f == index ? 14'h34 : _GEN_6734;
  wire [13:0] _GEN_6736 = 14'h1a50 == index ? 14'h34 : _GEN_6735;
  wire [13:0] _GEN_6737 = 14'h1a51 == index ? 14'h34 : _GEN_6736;
  wire [13:0] _GEN_6738 = 14'h1a52 == index ? 14'h34 : _GEN_6737;
  wire [13:0] _GEN_6739 = 14'h1a53 == index ? 14'h34 : _GEN_6738;
  wire [13:0] _GEN_6740 = 14'h1a54 == index ? 14'h34 : _GEN_6739;
  wire [13:0] _GEN_6741 = 14'h1a55 == index ? 14'h34 : _GEN_6740;
  wire [13:0] _GEN_6742 = 14'h1a56 == index ? 14'h34 : _GEN_6741;
  wire [13:0] _GEN_6743 = 14'h1a57 == index ? 14'h34 : _GEN_6742;
  wire [13:0] _GEN_6744 = 14'h1a58 == index ? 14'h34 : _GEN_6743;
  wire [13:0] _GEN_6745 = 14'h1a59 == index ? 14'h34 : _GEN_6744;
  wire [13:0] _GEN_6746 = 14'h1a5a == index ? 14'h34 : _GEN_6745;
  wire [13:0] _GEN_6747 = 14'h1a5b == index ? 14'h34 : _GEN_6746;
  wire [13:0] _GEN_6748 = 14'h1a5c == index ? 14'h34 : _GEN_6747;
  wire [13:0] _GEN_6749 = 14'h1a5d == index ? 14'h34 : _GEN_6748;
  wire [13:0] _GEN_6750 = 14'h1a5e == index ? 14'h34 : _GEN_6749;
  wire [13:0] _GEN_6751 = 14'h1a5f == index ? 14'h34 : _GEN_6750;
  wire [13:0] _GEN_6752 = 14'h1a60 == index ? 14'h34 : _GEN_6751;
  wire [13:0] _GEN_6753 = 14'h1a61 == index ? 14'h34 : _GEN_6752;
  wire [13:0] _GEN_6754 = 14'h1a62 == index ? 14'h34 : _GEN_6753;
  wire [13:0] _GEN_6755 = 14'h1a63 == index ? 14'h34 : _GEN_6754;
  wire [13:0] _GEN_6756 = 14'h1a64 == index ? 14'h34 : _GEN_6755;
  wire [13:0] _GEN_6757 = 14'h1a65 == index ? 14'h34 : _GEN_6756;
  wire [13:0] _GEN_6758 = 14'h1a66 == index ? 14'h34 : _GEN_6757;
  wire [13:0] _GEN_6759 = 14'h1a67 == index ? 14'h34 : _GEN_6758;
  wire [13:0] _GEN_6760 = 14'h1a68 == index ? 14'h34 : _GEN_6759;
  wire [13:0] _GEN_6761 = 14'h1a69 == index ? 14'h34 : _GEN_6760;
  wire [13:0] _GEN_6762 = 14'h1a6a == index ? 14'h34 : _GEN_6761;
  wire [13:0] _GEN_6763 = 14'h1a6b == index ? 14'h34 : _GEN_6762;
  wire [13:0] _GEN_6764 = 14'h1a6c == index ? 14'h34 : _GEN_6763;
  wire [13:0] _GEN_6765 = 14'h1a6d == index ? 14'h34 : _GEN_6764;
  wire [13:0] _GEN_6766 = 14'h1a6e == index ? 14'h34 : _GEN_6765;
  wire [13:0] _GEN_6767 = 14'h1a6f == index ? 14'h34 : _GEN_6766;
  wire [13:0] _GEN_6768 = 14'h1a70 == index ? 14'h34 : _GEN_6767;
  wire [13:0] _GEN_6769 = 14'h1a71 == index ? 14'h34 : _GEN_6768;
  wire [13:0] _GEN_6770 = 14'h1a72 == index ? 14'h34 : _GEN_6769;
  wire [13:0] _GEN_6771 = 14'h1a73 == index ? 14'h34 : _GEN_6770;
  wire [13:0] _GEN_6772 = 14'h1a74 == index ? 14'h34 : _GEN_6771;
  wire [13:0] _GEN_6773 = 14'h1a75 == index ? 14'h34 : _GEN_6772;
  wire [13:0] _GEN_6774 = 14'h1a76 == index ? 14'h34 : _GEN_6773;
  wire [13:0] _GEN_6775 = 14'h1a77 == index ? 14'h34 : _GEN_6774;
  wire [13:0] _GEN_6776 = 14'h1a78 == index ? 14'h34 : _GEN_6775;
  wire [13:0] _GEN_6777 = 14'h1a79 == index ? 14'h34 : _GEN_6776;
  wire [13:0] _GEN_6778 = 14'h1a7a == index ? 14'h34 : _GEN_6777;
  wire [13:0] _GEN_6779 = 14'h1a7b == index ? 14'h34 : _GEN_6778;
  wire [13:0] _GEN_6780 = 14'h1a7c == index ? 14'h34 : _GEN_6779;
  wire [13:0] _GEN_6781 = 14'h1a7d == index ? 14'h34 : _GEN_6780;
  wire [13:0] _GEN_6782 = 14'h1a7e == index ? 14'h34 : _GEN_6781;
  wire [13:0] _GEN_6783 = 14'h1a7f == index ? 14'h34 : _GEN_6782;
  wire [13:0] _GEN_6784 = 14'h1a80 == index ? 14'h0 : _GEN_6783;
  wire [13:0] _GEN_6785 = 14'h1a81 == index ? 14'h1a80 : _GEN_6784;
  wire [13:0] _GEN_6786 = 14'h1a82 == index ? 14'hd01 : _GEN_6785;
  wire [13:0] _GEN_6787 = 14'h1a83 == index ? 14'h882 : _GEN_6786;
  wire [13:0] _GEN_6788 = 14'h1a84 == index ? 14'h681 : _GEN_6787;
  wire [13:0] _GEN_6789 = 14'h1a85 == index ? 14'h503 : _GEN_6788;
  wire [13:0] _GEN_6790 = 14'h1a86 == index ? 14'h405 : _GEN_6789;
  wire [13:0] _GEN_6791 = 14'h1a87 == index ? 14'h384 : _GEN_6790;
  wire [13:0] _GEN_6792 = 14'h1a88 == index ? 14'h305 : _GEN_6791;
  wire [13:0] _GEN_6793 = 14'h1a89 == index ? 14'h288 : _GEN_6792;
  wire [13:0] _GEN_6794 = 14'h1a8a == index ? 14'h283 : _GEN_6793;
  wire [13:0] _GEN_6795 = 14'h1a8b == index ? 14'h209 : _GEN_6794;
  wire [13:0] _GEN_6796 = 14'h1a8c == index ? 14'h205 : _GEN_6795;
  wire [13:0] _GEN_6797 = 14'h1a8d == index ? 14'h201 : _GEN_6796;
  wire [13:0] _GEN_6798 = 14'h1a8e == index ? 14'h18b : _GEN_6797;
  wire [13:0] _GEN_6799 = 14'h1a8f == index ? 14'h188 : _GEN_6798;
  wire [13:0] _GEN_6800 = 14'h1a90 == index ? 14'h185 : _GEN_6799;
  wire [13:0] _GEN_6801 = 14'h1a91 == index ? 14'h182 : _GEN_6800;
  wire [13:0] _GEN_6802 = 14'h1a92 == index ? 14'h111 : _GEN_6801;
  wire [13:0] _GEN_6803 = 14'h1a93 == index ? 14'h10f : _GEN_6802;
  wire [13:0] _GEN_6804 = 14'h1a94 == index ? 14'h10d : _GEN_6803;
  wire [13:0] _GEN_6805 = 14'h1a95 == index ? 14'h10b : _GEN_6804;
  wire [13:0] _GEN_6806 = 14'h1a96 == index ? 14'h109 : _GEN_6805;
  wire [13:0] _GEN_6807 = 14'h1a97 == index ? 14'h107 : _GEN_6806;
  wire [13:0] _GEN_6808 = 14'h1a98 == index ? 14'h105 : _GEN_6807;
  wire [13:0] _GEN_6809 = 14'h1a99 == index ? 14'h103 : _GEN_6808;
  wire [13:0] _GEN_6810 = 14'h1a9a == index ? 14'h101 : _GEN_6809;
  wire [13:0] _GEN_6811 = 14'h1a9b == index ? 14'h9a : _GEN_6810;
  wire [13:0] _GEN_6812 = 14'h1a9c == index ? 14'h99 : _GEN_6811;
  wire [13:0] _GEN_6813 = 14'h1a9d == index ? 14'h98 : _GEN_6812;
  wire [13:0] _GEN_6814 = 14'h1a9e == index ? 14'h97 : _GEN_6813;
  wire [13:0] _GEN_6815 = 14'h1a9f == index ? 14'h96 : _GEN_6814;
  wire [13:0] _GEN_6816 = 14'h1aa0 == index ? 14'h95 : _GEN_6815;
  wire [13:0] _GEN_6817 = 14'h1aa1 == index ? 14'h94 : _GEN_6816;
  wire [13:0] _GEN_6818 = 14'h1aa2 == index ? 14'h93 : _GEN_6817;
  wire [13:0] _GEN_6819 = 14'h1aa3 == index ? 14'h92 : _GEN_6818;
  wire [13:0] _GEN_6820 = 14'h1aa4 == index ? 14'h91 : _GEN_6819;
  wire [13:0] _GEN_6821 = 14'h1aa5 == index ? 14'h90 : _GEN_6820;
  wire [13:0] _GEN_6822 = 14'h1aa6 == index ? 14'h8f : _GEN_6821;
  wire [13:0] _GEN_6823 = 14'h1aa7 == index ? 14'h8e : _GEN_6822;
  wire [13:0] _GEN_6824 = 14'h1aa8 == index ? 14'h8d : _GEN_6823;
  wire [13:0] _GEN_6825 = 14'h1aa9 == index ? 14'h8c : _GEN_6824;
  wire [13:0] _GEN_6826 = 14'h1aaa == index ? 14'h8b : _GEN_6825;
  wire [13:0] _GEN_6827 = 14'h1aab == index ? 14'h8a : _GEN_6826;
  wire [13:0] _GEN_6828 = 14'h1aac == index ? 14'h89 : _GEN_6827;
  wire [13:0] _GEN_6829 = 14'h1aad == index ? 14'h88 : _GEN_6828;
  wire [13:0] _GEN_6830 = 14'h1aae == index ? 14'h87 : _GEN_6829;
  wire [13:0] _GEN_6831 = 14'h1aaf == index ? 14'h86 : _GEN_6830;
  wire [13:0] _GEN_6832 = 14'h1ab0 == index ? 14'h85 : _GEN_6831;
  wire [13:0] _GEN_6833 = 14'h1ab1 == index ? 14'h84 : _GEN_6832;
  wire [13:0] _GEN_6834 = 14'h1ab2 == index ? 14'h83 : _GEN_6833;
  wire [13:0] _GEN_6835 = 14'h1ab3 == index ? 14'h82 : _GEN_6834;
  wire [13:0] _GEN_6836 = 14'h1ab4 == index ? 14'h81 : _GEN_6835;
  wire [13:0] _GEN_6837 = 14'h1ab5 == index ? 14'h80 : _GEN_6836;
  wire [13:0] _GEN_6838 = 14'h1ab6 == index ? 14'h35 : _GEN_6837;
  wire [13:0] _GEN_6839 = 14'h1ab7 == index ? 14'h35 : _GEN_6838;
  wire [13:0] _GEN_6840 = 14'h1ab8 == index ? 14'h35 : _GEN_6839;
  wire [13:0] _GEN_6841 = 14'h1ab9 == index ? 14'h35 : _GEN_6840;
  wire [13:0] _GEN_6842 = 14'h1aba == index ? 14'h35 : _GEN_6841;
  wire [13:0] _GEN_6843 = 14'h1abb == index ? 14'h35 : _GEN_6842;
  wire [13:0] _GEN_6844 = 14'h1abc == index ? 14'h35 : _GEN_6843;
  wire [13:0] _GEN_6845 = 14'h1abd == index ? 14'h35 : _GEN_6844;
  wire [13:0] _GEN_6846 = 14'h1abe == index ? 14'h35 : _GEN_6845;
  wire [13:0] _GEN_6847 = 14'h1abf == index ? 14'h35 : _GEN_6846;
  wire [13:0] _GEN_6848 = 14'h1ac0 == index ? 14'h35 : _GEN_6847;
  wire [13:0] _GEN_6849 = 14'h1ac1 == index ? 14'h35 : _GEN_6848;
  wire [13:0] _GEN_6850 = 14'h1ac2 == index ? 14'h35 : _GEN_6849;
  wire [13:0] _GEN_6851 = 14'h1ac3 == index ? 14'h35 : _GEN_6850;
  wire [13:0] _GEN_6852 = 14'h1ac4 == index ? 14'h35 : _GEN_6851;
  wire [13:0] _GEN_6853 = 14'h1ac5 == index ? 14'h35 : _GEN_6852;
  wire [13:0] _GEN_6854 = 14'h1ac6 == index ? 14'h35 : _GEN_6853;
  wire [13:0] _GEN_6855 = 14'h1ac7 == index ? 14'h35 : _GEN_6854;
  wire [13:0] _GEN_6856 = 14'h1ac8 == index ? 14'h35 : _GEN_6855;
  wire [13:0] _GEN_6857 = 14'h1ac9 == index ? 14'h35 : _GEN_6856;
  wire [13:0] _GEN_6858 = 14'h1aca == index ? 14'h35 : _GEN_6857;
  wire [13:0] _GEN_6859 = 14'h1acb == index ? 14'h35 : _GEN_6858;
  wire [13:0] _GEN_6860 = 14'h1acc == index ? 14'h35 : _GEN_6859;
  wire [13:0] _GEN_6861 = 14'h1acd == index ? 14'h35 : _GEN_6860;
  wire [13:0] _GEN_6862 = 14'h1ace == index ? 14'h35 : _GEN_6861;
  wire [13:0] _GEN_6863 = 14'h1acf == index ? 14'h35 : _GEN_6862;
  wire [13:0] _GEN_6864 = 14'h1ad0 == index ? 14'h35 : _GEN_6863;
  wire [13:0] _GEN_6865 = 14'h1ad1 == index ? 14'h35 : _GEN_6864;
  wire [13:0] _GEN_6866 = 14'h1ad2 == index ? 14'h35 : _GEN_6865;
  wire [13:0] _GEN_6867 = 14'h1ad3 == index ? 14'h35 : _GEN_6866;
  wire [13:0] _GEN_6868 = 14'h1ad4 == index ? 14'h35 : _GEN_6867;
  wire [13:0] _GEN_6869 = 14'h1ad5 == index ? 14'h35 : _GEN_6868;
  wire [13:0] _GEN_6870 = 14'h1ad6 == index ? 14'h35 : _GEN_6869;
  wire [13:0] _GEN_6871 = 14'h1ad7 == index ? 14'h35 : _GEN_6870;
  wire [13:0] _GEN_6872 = 14'h1ad8 == index ? 14'h35 : _GEN_6871;
  wire [13:0] _GEN_6873 = 14'h1ad9 == index ? 14'h35 : _GEN_6872;
  wire [13:0] _GEN_6874 = 14'h1ada == index ? 14'h35 : _GEN_6873;
  wire [13:0] _GEN_6875 = 14'h1adb == index ? 14'h35 : _GEN_6874;
  wire [13:0] _GEN_6876 = 14'h1adc == index ? 14'h35 : _GEN_6875;
  wire [13:0] _GEN_6877 = 14'h1add == index ? 14'h35 : _GEN_6876;
  wire [13:0] _GEN_6878 = 14'h1ade == index ? 14'h35 : _GEN_6877;
  wire [13:0] _GEN_6879 = 14'h1adf == index ? 14'h35 : _GEN_6878;
  wire [13:0] _GEN_6880 = 14'h1ae0 == index ? 14'h35 : _GEN_6879;
  wire [13:0] _GEN_6881 = 14'h1ae1 == index ? 14'h35 : _GEN_6880;
  wire [13:0] _GEN_6882 = 14'h1ae2 == index ? 14'h35 : _GEN_6881;
  wire [13:0] _GEN_6883 = 14'h1ae3 == index ? 14'h35 : _GEN_6882;
  wire [13:0] _GEN_6884 = 14'h1ae4 == index ? 14'h35 : _GEN_6883;
  wire [13:0] _GEN_6885 = 14'h1ae5 == index ? 14'h35 : _GEN_6884;
  wire [13:0] _GEN_6886 = 14'h1ae6 == index ? 14'h35 : _GEN_6885;
  wire [13:0] _GEN_6887 = 14'h1ae7 == index ? 14'h35 : _GEN_6886;
  wire [13:0] _GEN_6888 = 14'h1ae8 == index ? 14'h35 : _GEN_6887;
  wire [13:0] _GEN_6889 = 14'h1ae9 == index ? 14'h35 : _GEN_6888;
  wire [13:0] _GEN_6890 = 14'h1aea == index ? 14'h35 : _GEN_6889;
  wire [13:0] _GEN_6891 = 14'h1aeb == index ? 14'h35 : _GEN_6890;
  wire [13:0] _GEN_6892 = 14'h1aec == index ? 14'h35 : _GEN_6891;
  wire [13:0] _GEN_6893 = 14'h1aed == index ? 14'h35 : _GEN_6892;
  wire [13:0] _GEN_6894 = 14'h1aee == index ? 14'h35 : _GEN_6893;
  wire [13:0] _GEN_6895 = 14'h1aef == index ? 14'h35 : _GEN_6894;
  wire [13:0] _GEN_6896 = 14'h1af0 == index ? 14'h35 : _GEN_6895;
  wire [13:0] _GEN_6897 = 14'h1af1 == index ? 14'h35 : _GEN_6896;
  wire [13:0] _GEN_6898 = 14'h1af2 == index ? 14'h35 : _GEN_6897;
  wire [13:0] _GEN_6899 = 14'h1af3 == index ? 14'h35 : _GEN_6898;
  wire [13:0] _GEN_6900 = 14'h1af4 == index ? 14'h35 : _GEN_6899;
  wire [13:0] _GEN_6901 = 14'h1af5 == index ? 14'h35 : _GEN_6900;
  wire [13:0] _GEN_6902 = 14'h1af6 == index ? 14'h35 : _GEN_6901;
  wire [13:0] _GEN_6903 = 14'h1af7 == index ? 14'h35 : _GEN_6902;
  wire [13:0] _GEN_6904 = 14'h1af8 == index ? 14'h35 : _GEN_6903;
  wire [13:0] _GEN_6905 = 14'h1af9 == index ? 14'h35 : _GEN_6904;
  wire [13:0] _GEN_6906 = 14'h1afa == index ? 14'h35 : _GEN_6905;
  wire [13:0] _GEN_6907 = 14'h1afb == index ? 14'h35 : _GEN_6906;
  wire [13:0] _GEN_6908 = 14'h1afc == index ? 14'h35 : _GEN_6907;
  wire [13:0] _GEN_6909 = 14'h1afd == index ? 14'h35 : _GEN_6908;
  wire [13:0] _GEN_6910 = 14'h1afe == index ? 14'h35 : _GEN_6909;
  wire [13:0] _GEN_6911 = 14'h1aff == index ? 14'h35 : _GEN_6910;
  wire [13:0] _GEN_6912 = 14'h1b00 == index ? 14'h0 : _GEN_6911;
  wire [13:0] _GEN_6913 = 14'h1b01 == index ? 14'h1b00 : _GEN_6912;
  wire [13:0] _GEN_6914 = 14'h1b02 == index ? 14'hd80 : _GEN_6913;
  wire [13:0] _GEN_6915 = 14'h1b03 == index ? 14'h900 : _GEN_6914;
  wire [13:0] _GEN_6916 = 14'h1b04 == index ? 14'h682 : _GEN_6915;
  wire [13:0] _GEN_6917 = 14'h1b05 == index ? 14'h504 : _GEN_6916;
  wire [13:0] _GEN_6918 = 14'h1b06 == index ? 14'h480 : _GEN_6917;
  wire [13:0] _GEN_6919 = 14'h1b07 == index ? 14'h385 : _GEN_6918;
  wire [13:0] _GEN_6920 = 14'h1b08 == index ? 14'h306 : _GEN_6919;
  wire [13:0] _GEN_6921 = 14'h1b09 == index ? 14'h300 : _GEN_6920;
  wire [13:0] _GEN_6922 = 14'h1b0a == index ? 14'h284 : _GEN_6921;
  wire [13:0] _GEN_6923 = 14'h1b0b == index ? 14'h20a : _GEN_6922;
  wire [13:0] _GEN_6924 = 14'h1b0c == index ? 14'h206 : _GEN_6923;
  wire [13:0] _GEN_6925 = 14'h1b0d == index ? 14'h202 : _GEN_6924;
  wire [13:0] _GEN_6926 = 14'h1b0e == index ? 14'h18c : _GEN_6925;
  wire [13:0] _GEN_6927 = 14'h1b0f == index ? 14'h189 : _GEN_6926;
  wire [13:0] _GEN_6928 = 14'h1b10 == index ? 14'h186 : _GEN_6927;
  wire [13:0] _GEN_6929 = 14'h1b11 == index ? 14'h183 : _GEN_6928;
  wire [13:0] _GEN_6930 = 14'h1b12 == index ? 14'h180 : _GEN_6929;
  wire [13:0] _GEN_6931 = 14'h1b13 == index ? 14'h110 : _GEN_6930;
  wire [13:0] _GEN_6932 = 14'h1b14 == index ? 14'h10e : _GEN_6931;
  wire [13:0] _GEN_6933 = 14'h1b15 == index ? 14'h10c : _GEN_6932;
  wire [13:0] _GEN_6934 = 14'h1b16 == index ? 14'h10a : _GEN_6933;
  wire [13:0] _GEN_6935 = 14'h1b17 == index ? 14'h108 : _GEN_6934;
  wire [13:0] _GEN_6936 = 14'h1b18 == index ? 14'h106 : _GEN_6935;
  wire [13:0] _GEN_6937 = 14'h1b19 == index ? 14'h104 : _GEN_6936;
  wire [13:0] _GEN_6938 = 14'h1b1a == index ? 14'h102 : _GEN_6937;
  wire [13:0] _GEN_6939 = 14'h1b1b == index ? 14'h100 : _GEN_6938;
  wire [13:0] _GEN_6940 = 14'h1b1c == index ? 14'h9a : _GEN_6939;
  wire [13:0] _GEN_6941 = 14'h1b1d == index ? 14'h99 : _GEN_6940;
  wire [13:0] _GEN_6942 = 14'h1b1e == index ? 14'h98 : _GEN_6941;
  wire [13:0] _GEN_6943 = 14'h1b1f == index ? 14'h97 : _GEN_6942;
  wire [13:0] _GEN_6944 = 14'h1b20 == index ? 14'h96 : _GEN_6943;
  wire [13:0] _GEN_6945 = 14'h1b21 == index ? 14'h95 : _GEN_6944;
  wire [13:0] _GEN_6946 = 14'h1b22 == index ? 14'h94 : _GEN_6945;
  wire [13:0] _GEN_6947 = 14'h1b23 == index ? 14'h93 : _GEN_6946;
  wire [13:0] _GEN_6948 = 14'h1b24 == index ? 14'h92 : _GEN_6947;
  wire [13:0] _GEN_6949 = 14'h1b25 == index ? 14'h91 : _GEN_6948;
  wire [13:0] _GEN_6950 = 14'h1b26 == index ? 14'h90 : _GEN_6949;
  wire [13:0] _GEN_6951 = 14'h1b27 == index ? 14'h8f : _GEN_6950;
  wire [13:0] _GEN_6952 = 14'h1b28 == index ? 14'h8e : _GEN_6951;
  wire [13:0] _GEN_6953 = 14'h1b29 == index ? 14'h8d : _GEN_6952;
  wire [13:0] _GEN_6954 = 14'h1b2a == index ? 14'h8c : _GEN_6953;
  wire [13:0] _GEN_6955 = 14'h1b2b == index ? 14'h8b : _GEN_6954;
  wire [13:0] _GEN_6956 = 14'h1b2c == index ? 14'h8a : _GEN_6955;
  wire [13:0] _GEN_6957 = 14'h1b2d == index ? 14'h89 : _GEN_6956;
  wire [13:0] _GEN_6958 = 14'h1b2e == index ? 14'h88 : _GEN_6957;
  wire [13:0] _GEN_6959 = 14'h1b2f == index ? 14'h87 : _GEN_6958;
  wire [13:0] _GEN_6960 = 14'h1b30 == index ? 14'h86 : _GEN_6959;
  wire [13:0] _GEN_6961 = 14'h1b31 == index ? 14'h85 : _GEN_6960;
  wire [13:0] _GEN_6962 = 14'h1b32 == index ? 14'h84 : _GEN_6961;
  wire [13:0] _GEN_6963 = 14'h1b33 == index ? 14'h83 : _GEN_6962;
  wire [13:0] _GEN_6964 = 14'h1b34 == index ? 14'h82 : _GEN_6963;
  wire [13:0] _GEN_6965 = 14'h1b35 == index ? 14'h81 : _GEN_6964;
  wire [13:0] _GEN_6966 = 14'h1b36 == index ? 14'h80 : _GEN_6965;
  wire [13:0] _GEN_6967 = 14'h1b37 == index ? 14'h36 : _GEN_6966;
  wire [13:0] _GEN_6968 = 14'h1b38 == index ? 14'h36 : _GEN_6967;
  wire [13:0] _GEN_6969 = 14'h1b39 == index ? 14'h36 : _GEN_6968;
  wire [13:0] _GEN_6970 = 14'h1b3a == index ? 14'h36 : _GEN_6969;
  wire [13:0] _GEN_6971 = 14'h1b3b == index ? 14'h36 : _GEN_6970;
  wire [13:0] _GEN_6972 = 14'h1b3c == index ? 14'h36 : _GEN_6971;
  wire [13:0] _GEN_6973 = 14'h1b3d == index ? 14'h36 : _GEN_6972;
  wire [13:0] _GEN_6974 = 14'h1b3e == index ? 14'h36 : _GEN_6973;
  wire [13:0] _GEN_6975 = 14'h1b3f == index ? 14'h36 : _GEN_6974;
  wire [13:0] _GEN_6976 = 14'h1b40 == index ? 14'h36 : _GEN_6975;
  wire [13:0] _GEN_6977 = 14'h1b41 == index ? 14'h36 : _GEN_6976;
  wire [13:0] _GEN_6978 = 14'h1b42 == index ? 14'h36 : _GEN_6977;
  wire [13:0] _GEN_6979 = 14'h1b43 == index ? 14'h36 : _GEN_6978;
  wire [13:0] _GEN_6980 = 14'h1b44 == index ? 14'h36 : _GEN_6979;
  wire [13:0] _GEN_6981 = 14'h1b45 == index ? 14'h36 : _GEN_6980;
  wire [13:0] _GEN_6982 = 14'h1b46 == index ? 14'h36 : _GEN_6981;
  wire [13:0] _GEN_6983 = 14'h1b47 == index ? 14'h36 : _GEN_6982;
  wire [13:0] _GEN_6984 = 14'h1b48 == index ? 14'h36 : _GEN_6983;
  wire [13:0] _GEN_6985 = 14'h1b49 == index ? 14'h36 : _GEN_6984;
  wire [13:0] _GEN_6986 = 14'h1b4a == index ? 14'h36 : _GEN_6985;
  wire [13:0] _GEN_6987 = 14'h1b4b == index ? 14'h36 : _GEN_6986;
  wire [13:0] _GEN_6988 = 14'h1b4c == index ? 14'h36 : _GEN_6987;
  wire [13:0] _GEN_6989 = 14'h1b4d == index ? 14'h36 : _GEN_6988;
  wire [13:0] _GEN_6990 = 14'h1b4e == index ? 14'h36 : _GEN_6989;
  wire [13:0] _GEN_6991 = 14'h1b4f == index ? 14'h36 : _GEN_6990;
  wire [13:0] _GEN_6992 = 14'h1b50 == index ? 14'h36 : _GEN_6991;
  wire [13:0] _GEN_6993 = 14'h1b51 == index ? 14'h36 : _GEN_6992;
  wire [13:0] _GEN_6994 = 14'h1b52 == index ? 14'h36 : _GEN_6993;
  wire [13:0] _GEN_6995 = 14'h1b53 == index ? 14'h36 : _GEN_6994;
  wire [13:0] _GEN_6996 = 14'h1b54 == index ? 14'h36 : _GEN_6995;
  wire [13:0] _GEN_6997 = 14'h1b55 == index ? 14'h36 : _GEN_6996;
  wire [13:0] _GEN_6998 = 14'h1b56 == index ? 14'h36 : _GEN_6997;
  wire [13:0] _GEN_6999 = 14'h1b57 == index ? 14'h36 : _GEN_6998;
  wire [13:0] _GEN_7000 = 14'h1b58 == index ? 14'h36 : _GEN_6999;
  wire [13:0] _GEN_7001 = 14'h1b59 == index ? 14'h36 : _GEN_7000;
  wire [13:0] _GEN_7002 = 14'h1b5a == index ? 14'h36 : _GEN_7001;
  wire [13:0] _GEN_7003 = 14'h1b5b == index ? 14'h36 : _GEN_7002;
  wire [13:0] _GEN_7004 = 14'h1b5c == index ? 14'h36 : _GEN_7003;
  wire [13:0] _GEN_7005 = 14'h1b5d == index ? 14'h36 : _GEN_7004;
  wire [13:0] _GEN_7006 = 14'h1b5e == index ? 14'h36 : _GEN_7005;
  wire [13:0] _GEN_7007 = 14'h1b5f == index ? 14'h36 : _GEN_7006;
  wire [13:0] _GEN_7008 = 14'h1b60 == index ? 14'h36 : _GEN_7007;
  wire [13:0] _GEN_7009 = 14'h1b61 == index ? 14'h36 : _GEN_7008;
  wire [13:0] _GEN_7010 = 14'h1b62 == index ? 14'h36 : _GEN_7009;
  wire [13:0] _GEN_7011 = 14'h1b63 == index ? 14'h36 : _GEN_7010;
  wire [13:0] _GEN_7012 = 14'h1b64 == index ? 14'h36 : _GEN_7011;
  wire [13:0] _GEN_7013 = 14'h1b65 == index ? 14'h36 : _GEN_7012;
  wire [13:0] _GEN_7014 = 14'h1b66 == index ? 14'h36 : _GEN_7013;
  wire [13:0] _GEN_7015 = 14'h1b67 == index ? 14'h36 : _GEN_7014;
  wire [13:0] _GEN_7016 = 14'h1b68 == index ? 14'h36 : _GEN_7015;
  wire [13:0] _GEN_7017 = 14'h1b69 == index ? 14'h36 : _GEN_7016;
  wire [13:0] _GEN_7018 = 14'h1b6a == index ? 14'h36 : _GEN_7017;
  wire [13:0] _GEN_7019 = 14'h1b6b == index ? 14'h36 : _GEN_7018;
  wire [13:0] _GEN_7020 = 14'h1b6c == index ? 14'h36 : _GEN_7019;
  wire [13:0] _GEN_7021 = 14'h1b6d == index ? 14'h36 : _GEN_7020;
  wire [13:0] _GEN_7022 = 14'h1b6e == index ? 14'h36 : _GEN_7021;
  wire [13:0] _GEN_7023 = 14'h1b6f == index ? 14'h36 : _GEN_7022;
  wire [13:0] _GEN_7024 = 14'h1b70 == index ? 14'h36 : _GEN_7023;
  wire [13:0] _GEN_7025 = 14'h1b71 == index ? 14'h36 : _GEN_7024;
  wire [13:0] _GEN_7026 = 14'h1b72 == index ? 14'h36 : _GEN_7025;
  wire [13:0] _GEN_7027 = 14'h1b73 == index ? 14'h36 : _GEN_7026;
  wire [13:0] _GEN_7028 = 14'h1b74 == index ? 14'h36 : _GEN_7027;
  wire [13:0] _GEN_7029 = 14'h1b75 == index ? 14'h36 : _GEN_7028;
  wire [13:0] _GEN_7030 = 14'h1b76 == index ? 14'h36 : _GEN_7029;
  wire [13:0] _GEN_7031 = 14'h1b77 == index ? 14'h36 : _GEN_7030;
  wire [13:0] _GEN_7032 = 14'h1b78 == index ? 14'h36 : _GEN_7031;
  wire [13:0] _GEN_7033 = 14'h1b79 == index ? 14'h36 : _GEN_7032;
  wire [13:0] _GEN_7034 = 14'h1b7a == index ? 14'h36 : _GEN_7033;
  wire [13:0] _GEN_7035 = 14'h1b7b == index ? 14'h36 : _GEN_7034;
  wire [13:0] _GEN_7036 = 14'h1b7c == index ? 14'h36 : _GEN_7035;
  wire [13:0] _GEN_7037 = 14'h1b7d == index ? 14'h36 : _GEN_7036;
  wire [13:0] _GEN_7038 = 14'h1b7e == index ? 14'h36 : _GEN_7037;
  wire [13:0] _GEN_7039 = 14'h1b7f == index ? 14'h36 : _GEN_7038;
  wire [13:0] _GEN_7040 = 14'h1b80 == index ? 14'h0 : _GEN_7039;
  wire [13:0] _GEN_7041 = 14'h1b81 == index ? 14'h1b80 : _GEN_7040;
  wire [13:0] _GEN_7042 = 14'h1b82 == index ? 14'hd81 : _GEN_7041;
  wire [13:0] _GEN_7043 = 14'h1b83 == index ? 14'h901 : _GEN_7042;
  wire [13:0] _GEN_7044 = 14'h1b84 == index ? 14'h683 : _GEN_7043;
  wire [13:0] _GEN_7045 = 14'h1b85 == index ? 14'h580 : _GEN_7044;
  wire [13:0] _GEN_7046 = 14'h1b86 == index ? 14'h481 : _GEN_7045;
  wire [13:0] _GEN_7047 = 14'h1b87 == index ? 14'h386 : _GEN_7046;
  wire [13:0] _GEN_7048 = 14'h1b88 == index ? 14'h307 : _GEN_7047;
  wire [13:0] _GEN_7049 = 14'h1b89 == index ? 14'h301 : _GEN_7048;
  wire [13:0] _GEN_7050 = 14'h1b8a == index ? 14'h285 : _GEN_7049;
  wire [13:0] _GEN_7051 = 14'h1b8b == index ? 14'h280 : _GEN_7050;
  wire [13:0] _GEN_7052 = 14'h1b8c == index ? 14'h207 : _GEN_7051;
  wire [13:0] _GEN_7053 = 14'h1b8d == index ? 14'h203 : _GEN_7052;
  wire [13:0] _GEN_7054 = 14'h1b8e == index ? 14'h18d : _GEN_7053;
  wire [13:0] _GEN_7055 = 14'h1b8f == index ? 14'h18a : _GEN_7054;
  wire [13:0] _GEN_7056 = 14'h1b90 == index ? 14'h187 : _GEN_7055;
  wire [13:0] _GEN_7057 = 14'h1b91 == index ? 14'h184 : _GEN_7056;
  wire [13:0] _GEN_7058 = 14'h1b92 == index ? 14'h181 : _GEN_7057;
  wire [13:0] _GEN_7059 = 14'h1b93 == index ? 14'h111 : _GEN_7058;
  wire [13:0] _GEN_7060 = 14'h1b94 == index ? 14'h10f : _GEN_7059;
  wire [13:0] _GEN_7061 = 14'h1b95 == index ? 14'h10d : _GEN_7060;
  wire [13:0] _GEN_7062 = 14'h1b96 == index ? 14'h10b : _GEN_7061;
  wire [13:0] _GEN_7063 = 14'h1b97 == index ? 14'h109 : _GEN_7062;
  wire [13:0] _GEN_7064 = 14'h1b98 == index ? 14'h107 : _GEN_7063;
  wire [13:0] _GEN_7065 = 14'h1b99 == index ? 14'h105 : _GEN_7064;
  wire [13:0] _GEN_7066 = 14'h1b9a == index ? 14'h103 : _GEN_7065;
  wire [13:0] _GEN_7067 = 14'h1b9b == index ? 14'h101 : _GEN_7066;
  wire [13:0] _GEN_7068 = 14'h1b9c == index ? 14'h9b : _GEN_7067;
  wire [13:0] _GEN_7069 = 14'h1b9d == index ? 14'h9a : _GEN_7068;
  wire [13:0] _GEN_7070 = 14'h1b9e == index ? 14'h99 : _GEN_7069;
  wire [13:0] _GEN_7071 = 14'h1b9f == index ? 14'h98 : _GEN_7070;
  wire [13:0] _GEN_7072 = 14'h1ba0 == index ? 14'h97 : _GEN_7071;
  wire [13:0] _GEN_7073 = 14'h1ba1 == index ? 14'h96 : _GEN_7072;
  wire [13:0] _GEN_7074 = 14'h1ba2 == index ? 14'h95 : _GEN_7073;
  wire [13:0] _GEN_7075 = 14'h1ba3 == index ? 14'h94 : _GEN_7074;
  wire [13:0] _GEN_7076 = 14'h1ba4 == index ? 14'h93 : _GEN_7075;
  wire [13:0] _GEN_7077 = 14'h1ba5 == index ? 14'h92 : _GEN_7076;
  wire [13:0] _GEN_7078 = 14'h1ba6 == index ? 14'h91 : _GEN_7077;
  wire [13:0] _GEN_7079 = 14'h1ba7 == index ? 14'h90 : _GEN_7078;
  wire [13:0] _GEN_7080 = 14'h1ba8 == index ? 14'h8f : _GEN_7079;
  wire [13:0] _GEN_7081 = 14'h1ba9 == index ? 14'h8e : _GEN_7080;
  wire [13:0] _GEN_7082 = 14'h1baa == index ? 14'h8d : _GEN_7081;
  wire [13:0] _GEN_7083 = 14'h1bab == index ? 14'h8c : _GEN_7082;
  wire [13:0] _GEN_7084 = 14'h1bac == index ? 14'h8b : _GEN_7083;
  wire [13:0] _GEN_7085 = 14'h1bad == index ? 14'h8a : _GEN_7084;
  wire [13:0] _GEN_7086 = 14'h1bae == index ? 14'h89 : _GEN_7085;
  wire [13:0] _GEN_7087 = 14'h1baf == index ? 14'h88 : _GEN_7086;
  wire [13:0] _GEN_7088 = 14'h1bb0 == index ? 14'h87 : _GEN_7087;
  wire [13:0] _GEN_7089 = 14'h1bb1 == index ? 14'h86 : _GEN_7088;
  wire [13:0] _GEN_7090 = 14'h1bb2 == index ? 14'h85 : _GEN_7089;
  wire [13:0] _GEN_7091 = 14'h1bb3 == index ? 14'h84 : _GEN_7090;
  wire [13:0] _GEN_7092 = 14'h1bb4 == index ? 14'h83 : _GEN_7091;
  wire [13:0] _GEN_7093 = 14'h1bb5 == index ? 14'h82 : _GEN_7092;
  wire [13:0] _GEN_7094 = 14'h1bb6 == index ? 14'h81 : _GEN_7093;
  wire [13:0] _GEN_7095 = 14'h1bb7 == index ? 14'h80 : _GEN_7094;
  wire [13:0] _GEN_7096 = 14'h1bb8 == index ? 14'h37 : _GEN_7095;
  wire [13:0] _GEN_7097 = 14'h1bb9 == index ? 14'h37 : _GEN_7096;
  wire [13:0] _GEN_7098 = 14'h1bba == index ? 14'h37 : _GEN_7097;
  wire [13:0] _GEN_7099 = 14'h1bbb == index ? 14'h37 : _GEN_7098;
  wire [13:0] _GEN_7100 = 14'h1bbc == index ? 14'h37 : _GEN_7099;
  wire [13:0] _GEN_7101 = 14'h1bbd == index ? 14'h37 : _GEN_7100;
  wire [13:0] _GEN_7102 = 14'h1bbe == index ? 14'h37 : _GEN_7101;
  wire [13:0] _GEN_7103 = 14'h1bbf == index ? 14'h37 : _GEN_7102;
  wire [13:0] _GEN_7104 = 14'h1bc0 == index ? 14'h37 : _GEN_7103;
  wire [13:0] _GEN_7105 = 14'h1bc1 == index ? 14'h37 : _GEN_7104;
  wire [13:0] _GEN_7106 = 14'h1bc2 == index ? 14'h37 : _GEN_7105;
  wire [13:0] _GEN_7107 = 14'h1bc3 == index ? 14'h37 : _GEN_7106;
  wire [13:0] _GEN_7108 = 14'h1bc4 == index ? 14'h37 : _GEN_7107;
  wire [13:0] _GEN_7109 = 14'h1bc5 == index ? 14'h37 : _GEN_7108;
  wire [13:0] _GEN_7110 = 14'h1bc6 == index ? 14'h37 : _GEN_7109;
  wire [13:0] _GEN_7111 = 14'h1bc7 == index ? 14'h37 : _GEN_7110;
  wire [13:0] _GEN_7112 = 14'h1bc8 == index ? 14'h37 : _GEN_7111;
  wire [13:0] _GEN_7113 = 14'h1bc9 == index ? 14'h37 : _GEN_7112;
  wire [13:0] _GEN_7114 = 14'h1bca == index ? 14'h37 : _GEN_7113;
  wire [13:0] _GEN_7115 = 14'h1bcb == index ? 14'h37 : _GEN_7114;
  wire [13:0] _GEN_7116 = 14'h1bcc == index ? 14'h37 : _GEN_7115;
  wire [13:0] _GEN_7117 = 14'h1bcd == index ? 14'h37 : _GEN_7116;
  wire [13:0] _GEN_7118 = 14'h1bce == index ? 14'h37 : _GEN_7117;
  wire [13:0] _GEN_7119 = 14'h1bcf == index ? 14'h37 : _GEN_7118;
  wire [13:0] _GEN_7120 = 14'h1bd0 == index ? 14'h37 : _GEN_7119;
  wire [13:0] _GEN_7121 = 14'h1bd1 == index ? 14'h37 : _GEN_7120;
  wire [13:0] _GEN_7122 = 14'h1bd2 == index ? 14'h37 : _GEN_7121;
  wire [13:0] _GEN_7123 = 14'h1bd3 == index ? 14'h37 : _GEN_7122;
  wire [13:0] _GEN_7124 = 14'h1bd4 == index ? 14'h37 : _GEN_7123;
  wire [13:0] _GEN_7125 = 14'h1bd5 == index ? 14'h37 : _GEN_7124;
  wire [13:0] _GEN_7126 = 14'h1bd6 == index ? 14'h37 : _GEN_7125;
  wire [13:0] _GEN_7127 = 14'h1bd7 == index ? 14'h37 : _GEN_7126;
  wire [13:0] _GEN_7128 = 14'h1bd8 == index ? 14'h37 : _GEN_7127;
  wire [13:0] _GEN_7129 = 14'h1bd9 == index ? 14'h37 : _GEN_7128;
  wire [13:0] _GEN_7130 = 14'h1bda == index ? 14'h37 : _GEN_7129;
  wire [13:0] _GEN_7131 = 14'h1bdb == index ? 14'h37 : _GEN_7130;
  wire [13:0] _GEN_7132 = 14'h1bdc == index ? 14'h37 : _GEN_7131;
  wire [13:0] _GEN_7133 = 14'h1bdd == index ? 14'h37 : _GEN_7132;
  wire [13:0] _GEN_7134 = 14'h1bde == index ? 14'h37 : _GEN_7133;
  wire [13:0] _GEN_7135 = 14'h1bdf == index ? 14'h37 : _GEN_7134;
  wire [13:0] _GEN_7136 = 14'h1be0 == index ? 14'h37 : _GEN_7135;
  wire [13:0] _GEN_7137 = 14'h1be1 == index ? 14'h37 : _GEN_7136;
  wire [13:0] _GEN_7138 = 14'h1be2 == index ? 14'h37 : _GEN_7137;
  wire [13:0] _GEN_7139 = 14'h1be3 == index ? 14'h37 : _GEN_7138;
  wire [13:0] _GEN_7140 = 14'h1be4 == index ? 14'h37 : _GEN_7139;
  wire [13:0] _GEN_7141 = 14'h1be5 == index ? 14'h37 : _GEN_7140;
  wire [13:0] _GEN_7142 = 14'h1be6 == index ? 14'h37 : _GEN_7141;
  wire [13:0] _GEN_7143 = 14'h1be7 == index ? 14'h37 : _GEN_7142;
  wire [13:0] _GEN_7144 = 14'h1be8 == index ? 14'h37 : _GEN_7143;
  wire [13:0] _GEN_7145 = 14'h1be9 == index ? 14'h37 : _GEN_7144;
  wire [13:0] _GEN_7146 = 14'h1bea == index ? 14'h37 : _GEN_7145;
  wire [13:0] _GEN_7147 = 14'h1beb == index ? 14'h37 : _GEN_7146;
  wire [13:0] _GEN_7148 = 14'h1bec == index ? 14'h37 : _GEN_7147;
  wire [13:0] _GEN_7149 = 14'h1bed == index ? 14'h37 : _GEN_7148;
  wire [13:0] _GEN_7150 = 14'h1bee == index ? 14'h37 : _GEN_7149;
  wire [13:0] _GEN_7151 = 14'h1bef == index ? 14'h37 : _GEN_7150;
  wire [13:0] _GEN_7152 = 14'h1bf0 == index ? 14'h37 : _GEN_7151;
  wire [13:0] _GEN_7153 = 14'h1bf1 == index ? 14'h37 : _GEN_7152;
  wire [13:0] _GEN_7154 = 14'h1bf2 == index ? 14'h37 : _GEN_7153;
  wire [13:0] _GEN_7155 = 14'h1bf3 == index ? 14'h37 : _GEN_7154;
  wire [13:0] _GEN_7156 = 14'h1bf4 == index ? 14'h37 : _GEN_7155;
  wire [13:0] _GEN_7157 = 14'h1bf5 == index ? 14'h37 : _GEN_7156;
  wire [13:0] _GEN_7158 = 14'h1bf6 == index ? 14'h37 : _GEN_7157;
  wire [13:0] _GEN_7159 = 14'h1bf7 == index ? 14'h37 : _GEN_7158;
  wire [13:0] _GEN_7160 = 14'h1bf8 == index ? 14'h37 : _GEN_7159;
  wire [13:0] _GEN_7161 = 14'h1bf9 == index ? 14'h37 : _GEN_7160;
  wire [13:0] _GEN_7162 = 14'h1bfa == index ? 14'h37 : _GEN_7161;
  wire [13:0] _GEN_7163 = 14'h1bfb == index ? 14'h37 : _GEN_7162;
  wire [13:0] _GEN_7164 = 14'h1bfc == index ? 14'h37 : _GEN_7163;
  wire [13:0] _GEN_7165 = 14'h1bfd == index ? 14'h37 : _GEN_7164;
  wire [13:0] _GEN_7166 = 14'h1bfe == index ? 14'h37 : _GEN_7165;
  wire [13:0] _GEN_7167 = 14'h1bff == index ? 14'h37 : _GEN_7166;
  wire [13:0] _GEN_7168 = 14'h1c00 == index ? 14'h0 : _GEN_7167;
  wire [13:0] _GEN_7169 = 14'h1c01 == index ? 14'h1c00 : _GEN_7168;
  wire [13:0] _GEN_7170 = 14'h1c02 == index ? 14'he00 : _GEN_7169;
  wire [13:0] _GEN_7171 = 14'h1c03 == index ? 14'h902 : _GEN_7170;
  wire [13:0] _GEN_7172 = 14'h1c04 == index ? 14'h700 : _GEN_7171;
  wire [13:0] _GEN_7173 = 14'h1c05 == index ? 14'h581 : _GEN_7172;
  wire [13:0] _GEN_7174 = 14'h1c06 == index ? 14'h482 : _GEN_7173;
  wire [13:0] _GEN_7175 = 14'h1c07 == index ? 14'h400 : _GEN_7174;
  wire [13:0] _GEN_7176 = 14'h1c08 == index ? 14'h380 : _GEN_7175;
  wire [13:0] _GEN_7177 = 14'h1c09 == index ? 14'h302 : _GEN_7176;
  wire [13:0] _GEN_7178 = 14'h1c0a == index ? 14'h286 : _GEN_7177;
  wire [13:0] _GEN_7179 = 14'h1c0b == index ? 14'h281 : _GEN_7178;
  wire [13:0] _GEN_7180 = 14'h1c0c == index ? 14'h208 : _GEN_7179;
  wire [13:0] _GEN_7181 = 14'h1c0d == index ? 14'h204 : _GEN_7180;
  wire [13:0] _GEN_7182 = 14'h1c0e == index ? 14'h200 : _GEN_7181;
  wire [13:0] _GEN_7183 = 14'h1c0f == index ? 14'h18b : _GEN_7182;
  wire [13:0] _GEN_7184 = 14'h1c10 == index ? 14'h188 : _GEN_7183;
  wire [13:0] _GEN_7185 = 14'h1c11 == index ? 14'h185 : _GEN_7184;
  wire [13:0] _GEN_7186 = 14'h1c12 == index ? 14'h182 : _GEN_7185;
  wire [13:0] _GEN_7187 = 14'h1c13 == index ? 14'h112 : _GEN_7186;
  wire [13:0] _GEN_7188 = 14'h1c14 == index ? 14'h110 : _GEN_7187;
  wire [13:0] _GEN_7189 = 14'h1c15 == index ? 14'h10e : _GEN_7188;
  wire [13:0] _GEN_7190 = 14'h1c16 == index ? 14'h10c : _GEN_7189;
  wire [13:0] _GEN_7191 = 14'h1c17 == index ? 14'h10a : _GEN_7190;
  wire [13:0] _GEN_7192 = 14'h1c18 == index ? 14'h108 : _GEN_7191;
  wire [13:0] _GEN_7193 = 14'h1c19 == index ? 14'h106 : _GEN_7192;
  wire [13:0] _GEN_7194 = 14'h1c1a == index ? 14'h104 : _GEN_7193;
  wire [13:0] _GEN_7195 = 14'h1c1b == index ? 14'h102 : _GEN_7194;
  wire [13:0] _GEN_7196 = 14'h1c1c == index ? 14'h100 : _GEN_7195;
  wire [13:0] _GEN_7197 = 14'h1c1d == index ? 14'h9b : _GEN_7196;
  wire [13:0] _GEN_7198 = 14'h1c1e == index ? 14'h9a : _GEN_7197;
  wire [13:0] _GEN_7199 = 14'h1c1f == index ? 14'h99 : _GEN_7198;
  wire [13:0] _GEN_7200 = 14'h1c20 == index ? 14'h98 : _GEN_7199;
  wire [13:0] _GEN_7201 = 14'h1c21 == index ? 14'h97 : _GEN_7200;
  wire [13:0] _GEN_7202 = 14'h1c22 == index ? 14'h96 : _GEN_7201;
  wire [13:0] _GEN_7203 = 14'h1c23 == index ? 14'h95 : _GEN_7202;
  wire [13:0] _GEN_7204 = 14'h1c24 == index ? 14'h94 : _GEN_7203;
  wire [13:0] _GEN_7205 = 14'h1c25 == index ? 14'h93 : _GEN_7204;
  wire [13:0] _GEN_7206 = 14'h1c26 == index ? 14'h92 : _GEN_7205;
  wire [13:0] _GEN_7207 = 14'h1c27 == index ? 14'h91 : _GEN_7206;
  wire [13:0] _GEN_7208 = 14'h1c28 == index ? 14'h90 : _GEN_7207;
  wire [13:0] _GEN_7209 = 14'h1c29 == index ? 14'h8f : _GEN_7208;
  wire [13:0] _GEN_7210 = 14'h1c2a == index ? 14'h8e : _GEN_7209;
  wire [13:0] _GEN_7211 = 14'h1c2b == index ? 14'h8d : _GEN_7210;
  wire [13:0] _GEN_7212 = 14'h1c2c == index ? 14'h8c : _GEN_7211;
  wire [13:0] _GEN_7213 = 14'h1c2d == index ? 14'h8b : _GEN_7212;
  wire [13:0] _GEN_7214 = 14'h1c2e == index ? 14'h8a : _GEN_7213;
  wire [13:0] _GEN_7215 = 14'h1c2f == index ? 14'h89 : _GEN_7214;
  wire [13:0] _GEN_7216 = 14'h1c30 == index ? 14'h88 : _GEN_7215;
  wire [13:0] _GEN_7217 = 14'h1c31 == index ? 14'h87 : _GEN_7216;
  wire [13:0] _GEN_7218 = 14'h1c32 == index ? 14'h86 : _GEN_7217;
  wire [13:0] _GEN_7219 = 14'h1c33 == index ? 14'h85 : _GEN_7218;
  wire [13:0] _GEN_7220 = 14'h1c34 == index ? 14'h84 : _GEN_7219;
  wire [13:0] _GEN_7221 = 14'h1c35 == index ? 14'h83 : _GEN_7220;
  wire [13:0] _GEN_7222 = 14'h1c36 == index ? 14'h82 : _GEN_7221;
  wire [13:0] _GEN_7223 = 14'h1c37 == index ? 14'h81 : _GEN_7222;
  wire [13:0] _GEN_7224 = 14'h1c38 == index ? 14'h80 : _GEN_7223;
  wire [13:0] _GEN_7225 = 14'h1c39 == index ? 14'h38 : _GEN_7224;
  wire [13:0] _GEN_7226 = 14'h1c3a == index ? 14'h38 : _GEN_7225;
  wire [13:0] _GEN_7227 = 14'h1c3b == index ? 14'h38 : _GEN_7226;
  wire [13:0] _GEN_7228 = 14'h1c3c == index ? 14'h38 : _GEN_7227;
  wire [13:0] _GEN_7229 = 14'h1c3d == index ? 14'h38 : _GEN_7228;
  wire [13:0] _GEN_7230 = 14'h1c3e == index ? 14'h38 : _GEN_7229;
  wire [13:0] _GEN_7231 = 14'h1c3f == index ? 14'h38 : _GEN_7230;
  wire [13:0] _GEN_7232 = 14'h1c40 == index ? 14'h38 : _GEN_7231;
  wire [13:0] _GEN_7233 = 14'h1c41 == index ? 14'h38 : _GEN_7232;
  wire [13:0] _GEN_7234 = 14'h1c42 == index ? 14'h38 : _GEN_7233;
  wire [13:0] _GEN_7235 = 14'h1c43 == index ? 14'h38 : _GEN_7234;
  wire [13:0] _GEN_7236 = 14'h1c44 == index ? 14'h38 : _GEN_7235;
  wire [13:0] _GEN_7237 = 14'h1c45 == index ? 14'h38 : _GEN_7236;
  wire [13:0] _GEN_7238 = 14'h1c46 == index ? 14'h38 : _GEN_7237;
  wire [13:0] _GEN_7239 = 14'h1c47 == index ? 14'h38 : _GEN_7238;
  wire [13:0] _GEN_7240 = 14'h1c48 == index ? 14'h38 : _GEN_7239;
  wire [13:0] _GEN_7241 = 14'h1c49 == index ? 14'h38 : _GEN_7240;
  wire [13:0] _GEN_7242 = 14'h1c4a == index ? 14'h38 : _GEN_7241;
  wire [13:0] _GEN_7243 = 14'h1c4b == index ? 14'h38 : _GEN_7242;
  wire [13:0] _GEN_7244 = 14'h1c4c == index ? 14'h38 : _GEN_7243;
  wire [13:0] _GEN_7245 = 14'h1c4d == index ? 14'h38 : _GEN_7244;
  wire [13:0] _GEN_7246 = 14'h1c4e == index ? 14'h38 : _GEN_7245;
  wire [13:0] _GEN_7247 = 14'h1c4f == index ? 14'h38 : _GEN_7246;
  wire [13:0] _GEN_7248 = 14'h1c50 == index ? 14'h38 : _GEN_7247;
  wire [13:0] _GEN_7249 = 14'h1c51 == index ? 14'h38 : _GEN_7248;
  wire [13:0] _GEN_7250 = 14'h1c52 == index ? 14'h38 : _GEN_7249;
  wire [13:0] _GEN_7251 = 14'h1c53 == index ? 14'h38 : _GEN_7250;
  wire [13:0] _GEN_7252 = 14'h1c54 == index ? 14'h38 : _GEN_7251;
  wire [13:0] _GEN_7253 = 14'h1c55 == index ? 14'h38 : _GEN_7252;
  wire [13:0] _GEN_7254 = 14'h1c56 == index ? 14'h38 : _GEN_7253;
  wire [13:0] _GEN_7255 = 14'h1c57 == index ? 14'h38 : _GEN_7254;
  wire [13:0] _GEN_7256 = 14'h1c58 == index ? 14'h38 : _GEN_7255;
  wire [13:0] _GEN_7257 = 14'h1c59 == index ? 14'h38 : _GEN_7256;
  wire [13:0] _GEN_7258 = 14'h1c5a == index ? 14'h38 : _GEN_7257;
  wire [13:0] _GEN_7259 = 14'h1c5b == index ? 14'h38 : _GEN_7258;
  wire [13:0] _GEN_7260 = 14'h1c5c == index ? 14'h38 : _GEN_7259;
  wire [13:0] _GEN_7261 = 14'h1c5d == index ? 14'h38 : _GEN_7260;
  wire [13:0] _GEN_7262 = 14'h1c5e == index ? 14'h38 : _GEN_7261;
  wire [13:0] _GEN_7263 = 14'h1c5f == index ? 14'h38 : _GEN_7262;
  wire [13:0] _GEN_7264 = 14'h1c60 == index ? 14'h38 : _GEN_7263;
  wire [13:0] _GEN_7265 = 14'h1c61 == index ? 14'h38 : _GEN_7264;
  wire [13:0] _GEN_7266 = 14'h1c62 == index ? 14'h38 : _GEN_7265;
  wire [13:0] _GEN_7267 = 14'h1c63 == index ? 14'h38 : _GEN_7266;
  wire [13:0] _GEN_7268 = 14'h1c64 == index ? 14'h38 : _GEN_7267;
  wire [13:0] _GEN_7269 = 14'h1c65 == index ? 14'h38 : _GEN_7268;
  wire [13:0] _GEN_7270 = 14'h1c66 == index ? 14'h38 : _GEN_7269;
  wire [13:0] _GEN_7271 = 14'h1c67 == index ? 14'h38 : _GEN_7270;
  wire [13:0] _GEN_7272 = 14'h1c68 == index ? 14'h38 : _GEN_7271;
  wire [13:0] _GEN_7273 = 14'h1c69 == index ? 14'h38 : _GEN_7272;
  wire [13:0] _GEN_7274 = 14'h1c6a == index ? 14'h38 : _GEN_7273;
  wire [13:0] _GEN_7275 = 14'h1c6b == index ? 14'h38 : _GEN_7274;
  wire [13:0] _GEN_7276 = 14'h1c6c == index ? 14'h38 : _GEN_7275;
  wire [13:0] _GEN_7277 = 14'h1c6d == index ? 14'h38 : _GEN_7276;
  wire [13:0] _GEN_7278 = 14'h1c6e == index ? 14'h38 : _GEN_7277;
  wire [13:0] _GEN_7279 = 14'h1c6f == index ? 14'h38 : _GEN_7278;
  wire [13:0] _GEN_7280 = 14'h1c70 == index ? 14'h38 : _GEN_7279;
  wire [13:0] _GEN_7281 = 14'h1c71 == index ? 14'h38 : _GEN_7280;
  wire [13:0] _GEN_7282 = 14'h1c72 == index ? 14'h38 : _GEN_7281;
  wire [13:0] _GEN_7283 = 14'h1c73 == index ? 14'h38 : _GEN_7282;
  wire [13:0] _GEN_7284 = 14'h1c74 == index ? 14'h38 : _GEN_7283;
  wire [13:0] _GEN_7285 = 14'h1c75 == index ? 14'h38 : _GEN_7284;
  wire [13:0] _GEN_7286 = 14'h1c76 == index ? 14'h38 : _GEN_7285;
  wire [13:0] _GEN_7287 = 14'h1c77 == index ? 14'h38 : _GEN_7286;
  wire [13:0] _GEN_7288 = 14'h1c78 == index ? 14'h38 : _GEN_7287;
  wire [13:0] _GEN_7289 = 14'h1c79 == index ? 14'h38 : _GEN_7288;
  wire [13:0] _GEN_7290 = 14'h1c7a == index ? 14'h38 : _GEN_7289;
  wire [13:0] _GEN_7291 = 14'h1c7b == index ? 14'h38 : _GEN_7290;
  wire [13:0] _GEN_7292 = 14'h1c7c == index ? 14'h38 : _GEN_7291;
  wire [13:0] _GEN_7293 = 14'h1c7d == index ? 14'h38 : _GEN_7292;
  wire [13:0] _GEN_7294 = 14'h1c7e == index ? 14'h38 : _GEN_7293;
  wire [13:0] _GEN_7295 = 14'h1c7f == index ? 14'h38 : _GEN_7294;
  wire [13:0] _GEN_7296 = 14'h1c80 == index ? 14'h0 : _GEN_7295;
  wire [13:0] _GEN_7297 = 14'h1c81 == index ? 14'h1c80 : _GEN_7296;
  wire [13:0] _GEN_7298 = 14'h1c82 == index ? 14'he01 : _GEN_7297;
  wire [13:0] _GEN_7299 = 14'h1c83 == index ? 14'h980 : _GEN_7298;
  wire [13:0] _GEN_7300 = 14'h1c84 == index ? 14'h701 : _GEN_7299;
  wire [13:0] _GEN_7301 = 14'h1c85 == index ? 14'h582 : _GEN_7300;
  wire [13:0] _GEN_7302 = 14'h1c86 == index ? 14'h483 : _GEN_7301;
  wire [13:0] _GEN_7303 = 14'h1c87 == index ? 14'h401 : _GEN_7302;
  wire [13:0] _GEN_7304 = 14'h1c88 == index ? 14'h381 : _GEN_7303;
  wire [13:0] _GEN_7305 = 14'h1c89 == index ? 14'h303 : _GEN_7304;
  wire [13:0] _GEN_7306 = 14'h1c8a == index ? 14'h287 : _GEN_7305;
  wire [13:0] _GEN_7307 = 14'h1c8b == index ? 14'h282 : _GEN_7306;
  wire [13:0] _GEN_7308 = 14'h1c8c == index ? 14'h209 : _GEN_7307;
  wire [13:0] _GEN_7309 = 14'h1c8d == index ? 14'h205 : _GEN_7308;
  wire [13:0] _GEN_7310 = 14'h1c8e == index ? 14'h201 : _GEN_7309;
  wire [13:0] _GEN_7311 = 14'h1c8f == index ? 14'h18c : _GEN_7310;
  wire [13:0] _GEN_7312 = 14'h1c90 == index ? 14'h189 : _GEN_7311;
  wire [13:0] _GEN_7313 = 14'h1c91 == index ? 14'h186 : _GEN_7312;
  wire [13:0] _GEN_7314 = 14'h1c92 == index ? 14'h183 : _GEN_7313;
  wire [13:0] _GEN_7315 = 14'h1c93 == index ? 14'h180 : _GEN_7314;
  wire [13:0] _GEN_7316 = 14'h1c94 == index ? 14'h111 : _GEN_7315;
  wire [13:0] _GEN_7317 = 14'h1c95 == index ? 14'h10f : _GEN_7316;
  wire [13:0] _GEN_7318 = 14'h1c96 == index ? 14'h10d : _GEN_7317;
  wire [13:0] _GEN_7319 = 14'h1c97 == index ? 14'h10b : _GEN_7318;
  wire [13:0] _GEN_7320 = 14'h1c98 == index ? 14'h109 : _GEN_7319;
  wire [13:0] _GEN_7321 = 14'h1c99 == index ? 14'h107 : _GEN_7320;
  wire [13:0] _GEN_7322 = 14'h1c9a == index ? 14'h105 : _GEN_7321;
  wire [13:0] _GEN_7323 = 14'h1c9b == index ? 14'h103 : _GEN_7322;
  wire [13:0] _GEN_7324 = 14'h1c9c == index ? 14'h101 : _GEN_7323;
  wire [13:0] _GEN_7325 = 14'h1c9d == index ? 14'h9c : _GEN_7324;
  wire [13:0] _GEN_7326 = 14'h1c9e == index ? 14'h9b : _GEN_7325;
  wire [13:0] _GEN_7327 = 14'h1c9f == index ? 14'h9a : _GEN_7326;
  wire [13:0] _GEN_7328 = 14'h1ca0 == index ? 14'h99 : _GEN_7327;
  wire [13:0] _GEN_7329 = 14'h1ca1 == index ? 14'h98 : _GEN_7328;
  wire [13:0] _GEN_7330 = 14'h1ca2 == index ? 14'h97 : _GEN_7329;
  wire [13:0] _GEN_7331 = 14'h1ca3 == index ? 14'h96 : _GEN_7330;
  wire [13:0] _GEN_7332 = 14'h1ca4 == index ? 14'h95 : _GEN_7331;
  wire [13:0] _GEN_7333 = 14'h1ca5 == index ? 14'h94 : _GEN_7332;
  wire [13:0] _GEN_7334 = 14'h1ca6 == index ? 14'h93 : _GEN_7333;
  wire [13:0] _GEN_7335 = 14'h1ca7 == index ? 14'h92 : _GEN_7334;
  wire [13:0] _GEN_7336 = 14'h1ca8 == index ? 14'h91 : _GEN_7335;
  wire [13:0] _GEN_7337 = 14'h1ca9 == index ? 14'h90 : _GEN_7336;
  wire [13:0] _GEN_7338 = 14'h1caa == index ? 14'h8f : _GEN_7337;
  wire [13:0] _GEN_7339 = 14'h1cab == index ? 14'h8e : _GEN_7338;
  wire [13:0] _GEN_7340 = 14'h1cac == index ? 14'h8d : _GEN_7339;
  wire [13:0] _GEN_7341 = 14'h1cad == index ? 14'h8c : _GEN_7340;
  wire [13:0] _GEN_7342 = 14'h1cae == index ? 14'h8b : _GEN_7341;
  wire [13:0] _GEN_7343 = 14'h1caf == index ? 14'h8a : _GEN_7342;
  wire [13:0] _GEN_7344 = 14'h1cb0 == index ? 14'h89 : _GEN_7343;
  wire [13:0] _GEN_7345 = 14'h1cb1 == index ? 14'h88 : _GEN_7344;
  wire [13:0] _GEN_7346 = 14'h1cb2 == index ? 14'h87 : _GEN_7345;
  wire [13:0] _GEN_7347 = 14'h1cb3 == index ? 14'h86 : _GEN_7346;
  wire [13:0] _GEN_7348 = 14'h1cb4 == index ? 14'h85 : _GEN_7347;
  wire [13:0] _GEN_7349 = 14'h1cb5 == index ? 14'h84 : _GEN_7348;
  wire [13:0] _GEN_7350 = 14'h1cb6 == index ? 14'h83 : _GEN_7349;
  wire [13:0] _GEN_7351 = 14'h1cb7 == index ? 14'h82 : _GEN_7350;
  wire [13:0] _GEN_7352 = 14'h1cb8 == index ? 14'h81 : _GEN_7351;
  wire [13:0] _GEN_7353 = 14'h1cb9 == index ? 14'h80 : _GEN_7352;
  wire [13:0] _GEN_7354 = 14'h1cba == index ? 14'h39 : _GEN_7353;
  wire [13:0] _GEN_7355 = 14'h1cbb == index ? 14'h39 : _GEN_7354;
  wire [13:0] _GEN_7356 = 14'h1cbc == index ? 14'h39 : _GEN_7355;
  wire [13:0] _GEN_7357 = 14'h1cbd == index ? 14'h39 : _GEN_7356;
  wire [13:0] _GEN_7358 = 14'h1cbe == index ? 14'h39 : _GEN_7357;
  wire [13:0] _GEN_7359 = 14'h1cbf == index ? 14'h39 : _GEN_7358;
  wire [13:0] _GEN_7360 = 14'h1cc0 == index ? 14'h39 : _GEN_7359;
  wire [13:0] _GEN_7361 = 14'h1cc1 == index ? 14'h39 : _GEN_7360;
  wire [13:0] _GEN_7362 = 14'h1cc2 == index ? 14'h39 : _GEN_7361;
  wire [13:0] _GEN_7363 = 14'h1cc3 == index ? 14'h39 : _GEN_7362;
  wire [13:0] _GEN_7364 = 14'h1cc4 == index ? 14'h39 : _GEN_7363;
  wire [13:0] _GEN_7365 = 14'h1cc5 == index ? 14'h39 : _GEN_7364;
  wire [13:0] _GEN_7366 = 14'h1cc6 == index ? 14'h39 : _GEN_7365;
  wire [13:0] _GEN_7367 = 14'h1cc7 == index ? 14'h39 : _GEN_7366;
  wire [13:0] _GEN_7368 = 14'h1cc8 == index ? 14'h39 : _GEN_7367;
  wire [13:0] _GEN_7369 = 14'h1cc9 == index ? 14'h39 : _GEN_7368;
  wire [13:0] _GEN_7370 = 14'h1cca == index ? 14'h39 : _GEN_7369;
  wire [13:0] _GEN_7371 = 14'h1ccb == index ? 14'h39 : _GEN_7370;
  wire [13:0] _GEN_7372 = 14'h1ccc == index ? 14'h39 : _GEN_7371;
  wire [13:0] _GEN_7373 = 14'h1ccd == index ? 14'h39 : _GEN_7372;
  wire [13:0] _GEN_7374 = 14'h1cce == index ? 14'h39 : _GEN_7373;
  wire [13:0] _GEN_7375 = 14'h1ccf == index ? 14'h39 : _GEN_7374;
  wire [13:0] _GEN_7376 = 14'h1cd0 == index ? 14'h39 : _GEN_7375;
  wire [13:0] _GEN_7377 = 14'h1cd1 == index ? 14'h39 : _GEN_7376;
  wire [13:0] _GEN_7378 = 14'h1cd2 == index ? 14'h39 : _GEN_7377;
  wire [13:0] _GEN_7379 = 14'h1cd3 == index ? 14'h39 : _GEN_7378;
  wire [13:0] _GEN_7380 = 14'h1cd4 == index ? 14'h39 : _GEN_7379;
  wire [13:0] _GEN_7381 = 14'h1cd5 == index ? 14'h39 : _GEN_7380;
  wire [13:0] _GEN_7382 = 14'h1cd6 == index ? 14'h39 : _GEN_7381;
  wire [13:0] _GEN_7383 = 14'h1cd7 == index ? 14'h39 : _GEN_7382;
  wire [13:0] _GEN_7384 = 14'h1cd8 == index ? 14'h39 : _GEN_7383;
  wire [13:0] _GEN_7385 = 14'h1cd9 == index ? 14'h39 : _GEN_7384;
  wire [13:0] _GEN_7386 = 14'h1cda == index ? 14'h39 : _GEN_7385;
  wire [13:0] _GEN_7387 = 14'h1cdb == index ? 14'h39 : _GEN_7386;
  wire [13:0] _GEN_7388 = 14'h1cdc == index ? 14'h39 : _GEN_7387;
  wire [13:0] _GEN_7389 = 14'h1cdd == index ? 14'h39 : _GEN_7388;
  wire [13:0] _GEN_7390 = 14'h1cde == index ? 14'h39 : _GEN_7389;
  wire [13:0] _GEN_7391 = 14'h1cdf == index ? 14'h39 : _GEN_7390;
  wire [13:0] _GEN_7392 = 14'h1ce0 == index ? 14'h39 : _GEN_7391;
  wire [13:0] _GEN_7393 = 14'h1ce1 == index ? 14'h39 : _GEN_7392;
  wire [13:0] _GEN_7394 = 14'h1ce2 == index ? 14'h39 : _GEN_7393;
  wire [13:0] _GEN_7395 = 14'h1ce3 == index ? 14'h39 : _GEN_7394;
  wire [13:0] _GEN_7396 = 14'h1ce4 == index ? 14'h39 : _GEN_7395;
  wire [13:0] _GEN_7397 = 14'h1ce5 == index ? 14'h39 : _GEN_7396;
  wire [13:0] _GEN_7398 = 14'h1ce6 == index ? 14'h39 : _GEN_7397;
  wire [13:0] _GEN_7399 = 14'h1ce7 == index ? 14'h39 : _GEN_7398;
  wire [13:0] _GEN_7400 = 14'h1ce8 == index ? 14'h39 : _GEN_7399;
  wire [13:0] _GEN_7401 = 14'h1ce9 == index ? 14'h39 : _GEN_7400;
  wire [13:0] _GEN_7402 = 14'h1cea == index ? 14'h39 : _GEN_7401;
  wire [13:0] _GEN_7403 = 14'h1ceb == index ? 14'h39 : _GEN_7402;
  wire [13:0] _GEN_7404 = 14'h1cec == index ? 14'h39 : _GEN_7403;
  wire [13:0] _GEN_7405 = 14'h1ced == index ? 14'h39 : _GEN_7404;
  wire [13:0] _GEN_7406 = 14'h1cee == index ? 14'h39 : _GEN_7405;
  wire [13:0] _GEN_7407 = 14'h1cef == index ? 14'h39 : _GEN_7406;
  wire [13:0] _GEN_7408 = 14'h1cf0 == index ? 14'h39 : _GEN_7407;
  wire [13:0] _GEN_7409 = 14'h1cf1 == index ? 14'h39 : _GEN_7408;
  wire [13:0] _GEN_7410 = 14'h1cf2 == index ? 14'h39 : _GEN_7409;
  wire [13:0] _GEN_7411 = 14'h1cf3 == index ? 14'h39 : _GEN_7410;
  wire [13:0] _GEN_7412 = 14'h1cf4 == index ? 14'h39 : _GEN_7411;
  wire [13:0] _GEN_7413 = 14'h1cf5 == index ? 14'h39 : _GEN_7412;
  wire [13:0] _GEN_7414 = 14'h1cf6 == index ? 14'h39 : _GEN_7413;
  wire [13:0] _GEN_7415 = 14'h1cf7 == index ? 14'h39 : _GEN_7414;
  wire [13:0] _GEN_7416 = 14'h1cf8 == index ? 14'h39 : _GEN_7415;
  wire [13:0] _GEN_7417 = 14'h1cf9 == index ? 14'h39 : _GEN_7416;
  wire [13:0] _GEN_7418 = 14'h1cfa == index ? 14'h39 : _GEN_7417;
  wire [13:0] _GEN_7419 = 14'h1cfb == index ? 14'h39 : _GEN_7418;
  wire [13:0] _GEN_7420 = 14'h1cfc == index ? 14'h39 : _GEN_7419;
  wire [13:0] _GEN_7421 = 14'h1cfd == index ? 14'h39 : _GEN_7420;
  wire [13:0] _GEN_7422 = 14'h1cfe == index ? 14'h39 : _GEN_7421;
  wire [13:0] _GEN_7423 = 14'h1cff == index ? 14'h39 : _GEN_7422;
  wire [13:0] _GEN_7424 = 14'h1d00 == index ? 14'h0 : _GEN_7423;
  wire [13:0] _GEN_7425 = 14'h1d01 == index ? 14'h1d00 : _GEN_7424;
  wire [13:0] _GEN_7426 = 14'h1d02 == index ? 14'he80 : _GEN_7425;
  wire [13:0] _GEN_7427 = 14'h1d03 == index ? 14'h981 : _GEN_7426;
  wire [13:0] _GEN_7428 = 14'h1d04 == index ? 14'h702 : _GEN_7427;
  wire [13:0] _GEN_7429 = 14'h1d05 == index ? 14'h583 : _GEN_7428;
  wire [13:0] _GEN_7430 = 14'h1d06 == index ? 14'h484 : _GEN_7429;
  wire [13:0] _GEN_7431 = 14'h1d07 == index ? 14'h402 : _GEN_7430;
  wire [13:0] _GEN_7432 = 14'h1d08 == index ? 14'h382 : _GEN_7431;
  wire [13:0] _GEN_7433 = 14'h1d09 == index ? 14'h304 : _GEN_7432;
  wire [13:0] _GEN_7434 = 14'h1d0a == index ? 14'h288 : _GEN_7433;
  wire [13:0] _GEN_7435 = 14'h1d0b == index ? 14'h283 : _GEN_7434;
  wire [13:0] _GEN_7436 = 14'h1d0c == index ? 14'h20a : _GEN_7435;
  wire [13:0] _GEN_7437 = 14'h1d0d == index ? 14'h206 : _GEN_7436;
  wire [13:0] _GEN_7438 = 14'h1d0e == index ? 14'h202 : _GEN_7437;
  wire [13:0] _GEN_7439 = 14'h1d0f == index ? 14'h18d : _GEN_7438;
  wire [13:0] _GEN_7440 = 14'h1d10 == index ? 14'h18a : _GEN_7439;
  wire [13:0] _GEN_7441 = 14'h1d11 == index ? 14'h187 : _GEN_7440;
  wire [13:0] _GEN_7442 = 14'h1d12 == index ? 14'h184 : _GEN_7441;
  wire [13:0] _GEN_7443 = 14'h1d13 == index ? 14'h181 : _GEN_7442;
  wire [13:0] _GEN_7444 = 14'h1d14 == index ? 14'h112 : _GEN_7443;
  wire [13:0] _GEN_7445 = 14'h1d15 == index ? 14'h110 : _GEN_7444;
  wire [13:0] _GEN_7446 = 14'h1d16 == index ? 14'h10e : _GEN_7445;
  wire [13:0] _GEN_7447 = 14'h1d17 == index ? 14'h10c : _GEN_7446;
  wire [13:0] _GEN_7448 = 14'h1d18 == index ? 14'h10a : _GEN_7447;
  wire [13:0] _GEN_7449 = 14'h1d19 == index ? 14'h108 : _GEN_7448;
  wire [13:0] _GEN_7450 = 14'h1d1a == index ? 14'h106 : _GEN_7449;
  wire [13:0] _GEN_7451 = 14'h1d1b == index ? 14'h104 : _GEN_7450;
  wire [13:0] _GEN_7452 = 14'h1d1c == index ? 14'h102 : _GEN_7451;
  wire [13:0] _GEN_7453 = 14'h1d1d == index ? 14'h100 : _GEN_7452;
  wire [13:0] _GEN_7454 = 14'h1d1e == index ? 14'h9c : _GEN_7453;
  wire [13:0] _GEN_7455 = 14'h1d1f == index ? 14'h9b : _GEN_7454;
  wire [13:0] _GEN_7456 = 14'h1d20 == index ? 14'h9a : _GEN_7455;
  wire [13:0] _GEN_7457 = 14'h1d21 == index ? 14'h99 : _GEN_7456;
  wire [13:0] _GEN_7458 = 14'h1d22 == index ? 14'h98 : _GEN_7457;
  wire [13:0] _GEN_7459 = 14'h1d23 == index ? 14'h97 : _GEN_7458;
  wire [13:0] _GEN_7460 = 14'h1d24 == index ? 14'h96 : _GEN_7459;
  wire [13:0] _GEN_7461 = 14'h1d25 == index ? 14'h95 : _GEN_7460;
  wire [13:0] _GEN_7462 = 14'h1d26 == index ? 14'h94 : _GEN_7461;
  wire [13:0] _GEN_7463 = 14'h1d27 == index ? 14'h93 : _GEN_7462;
  wire [13:0] _GEN_7464 = 14'h1d28 == index ? 14'h92 : _GEN_7463;
  wire [13:0] _GEN_7465 = 14'h1d29 == index ? 14'h91 : _GEN_7464;
  wire [13:0] _GEN_7466 = 14'h1d2a == index ? 14'h90 : _GEN_7465;
  wire [13:0] _GEN_7467 = 14'h1d2b == index ? 14'h8f : _GEN_7466;
  wire [13:0] _GEN_7468 = 14'h1d2c == index ? 14'h8e : _GEN_7467;
  wire [13:0] _GEN_7469 = 14'h1d2d == index ? 14'h8d : _GEN_7468;
  wire [13:0] _GEN_7470 = 14'h1d2e == index ? 14'h8c : _GEN_7469;
  wire [13:0] _GEN_7471 = 14'h1d2f == index ? 14'h8b : _GEN_7470;
  wire [13:0] _GEN_7472 = 14'h1d30 == index ? 14'h8a : _GEN_7471;
  wire [13:0] _GEN_7473 = 14'h1d31 == index ? 14'h89 : _GEN_7472;
  wire [13:0] _GEN_7474 = 14'h1d32 == index ? 14'h88 : _GEN_7473;
  wire [13:0] _GEN_7475 = 14'h1d33 == index ? 14'h87 : _GEN_7474;
  wire [13:0] _GEN_7476 = 14'h1d34 == index ? 14'h86 : _GEN_7475;
  wire [13:0] _GEN_7477 = 14'h1d35 == index ? 14'h85 : _GEN_7476;
  wire [13:0] _GEN_7478 = 14'h1d36 == index ? 14'h84 : _GEN_7477;
  wire [13:0] _GEN_7479 = 14'h1d37 == index ? 14'h83 : _GEN_7478;
  wire [13:0] _GEN_7480 = 14'h1d38 == index ? 14'h82 : _GEN_7479;
  wire [13:0] _GEN_7481 = 14'h1d39 == index ? 14'h81 : _GEN_7480;
  wire [13:0] _GEN_7482 = 14'h1d3a == index ? 14'h80 : _GEN_7481;
  wire [13:0] _GEN_7483 = 14'h1d3b == index ? 14'h3a : _GEN_7482;
  wire [13:0] _GEN_7484 = 14'h1d3c == index ? 14'h3a : _GEN_7483;
  wire [13:0] _GEN_7485 = 14'h1d3d == index ? 14'h3a : _GEN_7484;
  wire [13:0] _GEN_7486 = 14'h1d3e == index ? 14'h3a : _GEN_7485;
  wire [13:0] _GEN_7487 = 14'h1d3f == index ? 14'h3a : _GEN_7486;
  wire [13:0] _GEN_7488 = 14'h1d40 == index ? 14'h3a : _GEN_7487;
  wire [13:0] _GEN_7489 = 14'h1d41 == index ? 14'h3a : _GEN_7488;
  wire [13:0] _GEN_7490 = 14'h1d42 == index ? 14'h3a : _GEN_7489;
  wire [13:0] _GEN_7491 = 14'h1d43 == index ? 14'h3a : _GEN_7490;
  wire [13:0] _GEN_7492 = 14'h1d44 == index ? 14'h3a : _GEN_7491;
  wire [13:0] _GEN_7493 = 14'h1d45 == index ? 14'h3a : _GEN_7492;
  wire [13:0] _GEN_7494 = 14'h1d46 == index ? 14'h3a : _GEN_7493;
  wire [13:0] _GEN_7495 = 14'h1d47 == index ? 14'h3a : _GEN_7494;
  wire [13:0] _GEN_7496 = 14'h1d48 == index ? 14'h3a : _GEN_7495;
  wire [13:0] _GEN_7497 = 14'h1d49 == index ? 14'h3a : _GEN_7496;
  wire [13:0] _GEN_7498 = 14'h1d4a == index ? 14'h3a : _GEN_7497;
  wire [13:0] _GEN_7499 = 14'h1d4b == index ? 14'h3a : _GEN_7498;
  wire [13:0] _GEN_7500 = 14'h1d4c == index ? 14'h3a : _GEN_7499;
  wire [13:0] _GEN_7501 = 14'h1d4d == index ? 14'h3a : _GEN_7500;
  wire [13:0] _GEN_7502 = 14'h1d4e == index ? 14'h3a : _GEN_7501;
  wire [13:0] _GEN_7503 = 14'h1d4f == index ? 14'h3a : _GEN_7502;
  wire [13:0] _GEN_7504 = 14'h1d50 == index ? 14'h3a : _GEN_7503;
  wire [13:0] _GEN_7505 = 14'h1d51 == index ? 14'h3a : _GEN_7504;
  wire [13:0] _GEN_7506 = 14'h1d52 == index ? 14'h3a : _GEN_7505;
  wire [13:0] _GEN_7507 = 14'h1d53 == index ? 14'h3a : _GEN_7506;
  wire [13:0] _GEN_7508 = 14'h1d54 == index ? 14'h3a : _GEN_7507;
  wire [13:0] _GEN_7509 = 14'h1d55 == index ? 14'h3a : _GEN_7508;
  wire [13:0] _GEN_7510 = 14'h1d56 == index ? 14'h3a : _GEN_7509;
  wire [13:0] _GEN_7511 = 14'h1d57 == index ? 14'h3a : _GEN_7510;
  wire [13:0] _GEN_7512 = 14'h1d58 == index ? 14'h3a : _GEN_7511;
  wire [13:0] _GEN_7513 = 14'h1d59 == index ? 14'h3a : _GEN_7512;
  wire [13:0] _GEN_7514 = 14'h1d5a == index ? 14'h3a : _GEN_7513;
  wire [13:0] _GEN_7515 = 14'h1d5b == index ? 14'h3a : _GEN_7514;
  wire [13:0] _GEN_7516 = 14'h1d5c == index ? 14'h3a : _GEN_7515;
  wire [13:0] _GEN_7517 = 14'h1d5d == index ? 14'h3a : _GEN_7516;
  wire [13:0] _GEN_7518 = 14'h1d5e == index ? 14'h3a : _GEN_7517;
  wire [13:0] _GEN_7519 = 14'h1d5f == index ? 14'h3a : _GEN_7518;
  wire [13:0] _GEN_7520 = 14'h1d60 == index ? 14'h3a : _GEN_7519;
  wire [13:0] _GEN_7521 = 14'h1d61 == index ? 14'h3a : _GEN_7520;
  wire [13:0] _GEN_7522 = 14'h1d62 == index ? 14'h3a : _GEN_7521;
  wire [13:0] _GEN_7523 = 14'h1d63 == index ? 14'h3a : _GEN_7522;
  wire [13:0] _GEN_7524 = 14'h1d64 == index ? 14'h3a : _GEN_7523;
  wire [13:0] _GEN_7525 = 14'h1d65 == index ? 14'h3a : _GEN_7524;
  wire [13:0] _GEN_7526 = 14'h1d66 == index ? 14'h3a : _GEN_7525;
  wire [13:0] _GEN_7527 = 14'h1d67 == index ? 14'h3a : _GEN_7526;
  wire [13:0] _GEN_7528 = 14'h1d68 == index ? 14'h3a : _GEN_7527;
  wire [13:0] _GEN_7529 = 14'h1d69 == index ? 14'h3a : _GEN_7528;
  wire [13:0] _GEN_7530 = 14'h1d6a == index ? 14'h3a : _GEN_7529;
  wire [13:0] _GEN_7531 = 14'h1d6b == index ? 14'h3a : _GEN_7530;
  wire [13:0] _GEN_7532 = 14'h1d6c == index ? 14'h3a : _GEN_7531;
  wire [13:0] _GEN_7533 = 14'h1d6d == index ? 14'h3a : _GEN_7532;
  wire [13:0] _GEN_7534 = 14'h1d6e == index ? 14'h3a : _GEN_7533;
  wire [13:0] _GEN_7535 = 14'h1d6f == index ? 14'h3a : _GEN_7534;
  wire [13:0] _GEN_7536 = 14'h1d70 == index ? 14'h3a : _GEN_7535;
  wire [13:0] _GEN_7537 = 14'h1d71 == index ? 14'h3a : _GEN_7536;
  wire [13:0] _GEN_7538 = 14'h1d72 == index ? 14'h3a : _GEN_7537;
  wire [13:0] _GEN_7539 = 14'h1d73 == index ? 14'h3a : _GEN_7538;
  wire [13:0] _GEN_7540 = 14'h1d74 == index ? 14'h3a : _GEN_7539;
  wire [13:0] _GEN_7541 = 14'h1d75 == index ? 14'h3a : _GEN_7540;
  wire [13:0] _GEN_7542 = 14'h1d76 == index ? 14'h3a : _GEN_7541;
  wire [13:0] _GEN_7543 = 14'h1d77 == index ? 14'h3a : _GEN_7542;
  wire [13:0] _GEN_7544 = 14'h1d78 == index ? 14'h3a : _GEN_7543;
  wire [13:0] _GEN_7545 = 14'h1d79 == index ? 14'h3a : _GEN_7544;
  wire [13:0] _GEN_7546 = 14'h1d7a == index ? 14'h3a : _GEN_7545;
  wire [13:0] _GEN_7547 = 14'h1d7b == index ? 14'h3a : _GEN_7546;
  wire [13:0] _GEN_7548 = 14'h1d7c == index ? 14'h3a : _GEN_7547;
  wire [13:0] _GEN_7549 = 14'h1d7d == index ? 14'h3a : _GEN_7548;
  wire [13:0] _GEN_7550 = 14'h1d7e == index ? 14'h3a : _GEN_7549;
  wire [13:0] _GEN_7551 = 14'h1d7f == index ? 14'h3a : _GEN_7550;
  wire [13:0] _GEN_7552 = 14'h1d80 == index ? 14'h0 : _GEN_7551;
  wire [13:0] _GEN_7553 = 14'h1d81 == index ? 14'h1d80 : _GEN_7552;
  wire [13:0] _GEN_7554 = 14'h1d82 == index ? 14'he81 : _GEN_7553;
  wire [13:0] _GEN_7555 = 14'h1d83 == index ? 14'h982 : _GEN_7554;
  wire [13:0] _GEN_7556 = 14'h1d84 == index ? 14'h703 : _GEN_7555;
  wire [13:0] _GEN_7557 = 14'h1d85 == index ? 14'h584 : _GEN_7556;
  wire [13:0] _GEN_7558 = 14'h1d86 == index ? 14'h485 : _GEN_7557;
  wire [13:0] _GEN_7559 = 14'h1d87 == index ? 14'h403 : _GEN_7558;
  wire [13:0] _GEN_7560 = 14'h1d88 == index ? 14'h383 : _GEN_7559;
  wire [13:0] _GEN_7561 = 14'h1d89 == index ? 14'h305 : _GEN_7560;
  wire [13:0] _GEN_7562 = 14'h1d8a == index ? 14'h289 : _GEN_7561;
  wire [13:0] _GEN_7563 = 14'h1d8b == index ? 14'h284 : _GEN_7562;
  wire [13:0] _GEN_7564 = 14'h1d8c == index ? 14'h20b : _GEN_7563;
  wire [13:0] _GEN_7565 = 14'h1d8d == index ? 14'h207 : _GEN_7564;
  wire [13:0] _GEN_7566 = 14'h1d8e == index ? 14'h203 : _GEN_7565;
  wire [13:0] _GEN_7567 = 14'h1d8f == index ? 14'h18e : _GEN_7566;
  wire [13:0] _GEN_7568 = 14'h1d90 == index ? 14'h18b : _GEN_7567;
  wire [13:0] _GEN_7569 = 14'h1d91 == index ? 14'h188 : _GEN_7568;
  wire [13:0] _GEN_7570 = 14'h1d92 == index ? 14'h185 : _GEN_7569;
  wire [13:0] _GEN_7571 = 14'h1d93 == index ? 14'h182 : _GEN_7570;
  wire [13:0] _GEN_7572 = 14'h1d94 == index ? 14'h113 : _GEN_7571;
  wire [13:0] _GEN_7573 = 14'h1d95 == index ? 14'h111 : _GEN_7572;
  wire [13:0] _GEN_7574 = 14'h1d96 == index ? 14'h10f : _GEN_7573;
  wire [13:0] _GEN_7575 = 14'h1d97 == index ? 14'h10d : _GEN_7574;
  wire [13:0] _GEN_7576 = 14'h1d98 == index ? 14'h10b : _GEN_7575;
  wire [13:0] _GEN_7577 = 14'h1d99 == index ? 14'h109 : _GEN_7576;
  wire [13:0] _GEN_7578 = 14'h1d9a == index ? 14'h107 : _GEN_7577;
  wire [13:0] _GEN_7579 = 14'h1d9b == index ? 14'h105 : _GEN_7578;
  wire [13:0] _GEN_7580 = 14'h1d9c == index ? 14'h103 : _GEN_7579;
  wire [13:0] _GEN_7581 = 14'h1d9d == index ? 14'h101 : _GEN_7580;
  wire [13:0] _GEN_7582 = 14'h1d9e == index ? 14'h9d : _GEN_7581;
  wire [13:0] _GEN_7583 = 14'h1d9f == index ? 14'h9c : _GEN_7582;
  wire [13:0] _GEN_7584 = 14'h1da0 == index ? 14'h9b : _GEN_7583;
  wire [13:0] _GEN_7585 = 14'h1da1 == index ? 14'h9a : _GEN_7584;
  wire [13:0] _GEN_7586 = 14'h1da2 == index ? 14'h99 : _GEN_7585;
  wire [13:0] _GEN_7587 = 14'h1da3 == index ? 14'h98 : _GEN_7586;
  wire [13:0] _GEN_7588 = 14'h1da4 == index ? 14'h97 : _GEN_7587;
  wire [13:0] _GEN_7589 = 14'h1da5 == index ? 14'h96 : _GEN_7588;
  wire [13:0] _GEN_7590 = 14'h1da6 == index ? 14'h95 : _GEN_7589;
  wire [13:0] _GEN_7591 = 14'h1da7 == index ? 14'h94 : _GEN_7590;
  wire [13:0] _GEN_7592 = 14'h1da8 == index ? 14'h93 : _GEN_7591;
  wire [13:0] _GEN_7593 = 14'h1da9 == index ? 14'h92 : _GEN_7592;
  wire [13:0] _GEN_7594 = 14'h1daa == index ? 14'h91 : _GEN_7593;
  wire [13:0] _GEN_7595 = 14'h1dab == index ? 14'h90 : _GEN_7594;
  wire [13:0] _GEN_7596 = 14'h1dac == index ? 14'h8f : _GEN_7595;
  wire [13:0] _GEN_7597 = 14'h1dad == index ? 14'h8e : _GEN_7596;
  wire [13:0] _GEN_7598 = 14'h1dae == index ? 14'h8d : _GEN_7597;
  wire [13:0] _GEN_7599 = 14'h1daf == index ? 14'h8c : _GEN_7598;
  wire [13:0] _GEN_7600 = 14'h1db0 == index ? 14'h8b : _GEN_7599;
  wire [13:0] _GEN_7601 = 14'h1db1 == index ? 14'h8a : _GEN_7600;
  wire [13:0] _GEN_7602 = 14'h1db2 == index ? 14'h89 : _GEN_7601;
  wire [13:0] _GEN_7603 = 14'h1db3 == index ? 14'h88 : _GEN_7602;
  wire [13:0] _GEN_7604 = 14'h1db4 == index ? 14'h87 : _GEN_7603;
  wire [13:0] _GEN_7605 = 14'h1db5 == index ? 14'h86 : _GEN_7604;
  wire [13:0] _GEN_7606 = 14'h1db6 == index ? 14'h85 : _GEN_7605;
  wire [13:0] _GEN_7607 = 14'h1db7 == index ? 14'h84 : _GEN_7606;
  wire [13:0] _GEN_7608 = 14'h1db8 == index ? 14'h83 : _GEN_7607;
  wire [13:0] _GEN_7609 = 14'h1db9 == index ? 14'h82 : _GEN_7608;
  wire [13:0] _GEN_7610 = 14'h1dba == index ? 14'h81 : _GEN_7609;
  wire [13:0] _GEN_7611 = 14'h1dbb == index ? 14'h80 : _GEN_7610;
  wire [13:0] _GEN_7612 = 14'h1dbc == index ? 14'h3b : _GEN_7611;
  wire [13:0] _GEN_7613 = 14'h1dbd == index ? 14'h3b : _GEN_7612;
  wire [13:0] _GEN_7614 = 14'h1dbe == index ? 14'h3b : _GEN_7613;
  wire [13:0] _GEN_7615 = 14'h1dbf == index ? 14'h3b : _GEN_7614;
  wire [13:0] _GEN_7616 = 14'h1dc0 == index ? 14'h3b : _GEN_7615;
  wire [13:0] _GEN_7617 = 14'h1dc1 == index ? 14'h3b : _GEN_7616;
  wire [13:0] _GEN_7618 = 14'h1dc2 == index ? 14'h3b : _GEN_7617;
  wire [13:0] _GEN_7619 = 14'h1dc3 == index ? 14'h3b : _GEN_7618;
  wire [13:0] _GEN_7620 = 14'h1dc4 == index ? 14'h3b : _GEN_7619;
  wire [13:0] _GEN_7621 = 14'h1dc5 == index ? 14'h3b : _GEN_7620;
  wire [13:0] _GEN_7622 = 14'h1dc6 == index ? 14'h3b : _GEN_7621;
  wire [13:0] _GEN_7623 = 14'h1dc7 == index ? 14'h3b : _GEN_7622;
  wire [13:0] _GEN_7624 = 14'h1dc8 == index ? 14'h3b : _GEN_7623;
  wire [13:0] _GEN_7625 = 14'h1dc9 == index ? 14'h3b : _GEN_7624;
  wire [13:0] _GEN_7626 = 14'h1dca == index ? 14'h3b : _GEN_7625;
  wire [13:0] _GEN_7627 = 14'h1dcb == index ? 14'h3b : _GEN_7626;
  wire [13:0] _GEN_7628 = 14'h1dcc == index ? 14'h3b : _GEN_7627;
  wire [13:0] _GEN_7629 = 14'h1dcd == index ? 14'h3b : _GEN_7628;
  wire [13:0] _GEN_7630 = 14'h1dce == index ? 14'h3b : _GEN_7629;
  wire [13:0] _GEN_7631 = 14'h1dcf == index ? 14'h3b : _GEN_7630;
  wire [13:0] _GEN_7632 = 14'h1dd0 == index ? 14'h3b : _GEN_7631;
  wire [13:0] _GEN_7633 = 14'h1dd1 == index ? 14'h3b : _GEN_7632;
  wire [13:0] _GEN_7634 = 14'h1dd2 == index ? 14'h3b : _GEN_7633;
  wire [13:0] _GEN_7635 = 14'h1dd3 == index ? 14'h3b : _GEN_7634;
  wire [13:0] _GEN_7636 = 14'h1dd4 == index ? 14'h3b : _GEN_7635;
  wire [13:0] _GEN_7637 = 14'h1dd5 == index ? 14'h3b : _GEN_7636;
  wire [13:0] _GEN_7638 = 14'h1dd6 == index ? 14'h3b : _GEN_7637;
  wire [13:0] _GEN_7639 = 14'h1dd7 == index ? 14'h3b : _GEN_7638;
  wire [13:0] _GEN_7640 = 14'h1dd8 == index ? 14'h3b : _GEN_7639;
  wire [13:0] _GEN_7641 = 14'h1dd9 == index ? 14'h3b : _GEN_7640;
  wire [13:0] _GEN_7642 = 14'h1dda == index ? 14'h3b : _GEN_7641;
  wire [13:0] _GEN_7643 = 14'h1ddb == index ? 14'h3b : _GEN_7642;
  wire [13:0] _GEN_7644 = 14'h1ddc == index ? 14'h3b : _GEN_7643;
  wire [13:0] _GEN_7645 = 14'h1ddd == index ? 14'h3b : _GEN_7644;
  wire [13:0] _GEN_7646 = 14'h1dde == index ? 14'h3b : _GEN_7645;
  wire [13:0] _GEN_7647 = 14'h1ddf == index ? 14'h3b : _GEN_7646;
  wire [13:0] _GEN_7648 = 14'h1de0 == index ? 14'h3b : _GEN_7647;
  wire [13:0] _GEN_7649 = 14'h1de1 == index ? 14'h3b : _GEN_7648;
  wire [13:0] _GEN_7650 = 14'h1de2 == index ? 14'h3b : _GEN_7649;
  wire [13:0] _GEN_7651 = 14'h1de3 == index ? 14'h3b : _GEN_7650;
  wire [13:0] _GEN_7652 = 14'h1de4 == index ? 14'h3b : _GEN_7651;
  wire [13:0] _GEN_7653 = 14'h1de5 == index ? 14'h3b : _GEN_7652;
  wire [13:0] _GEN_7654 = 14'h1de6 == index ? 14'h3b : _GEN_7653;
  wire [13:0] _GEN_7655 = 14'h1de7 == index ? 14'h3b : _GEN_7654;
  wire [13:0] _GEN_7656 = 14'h1de8 == index ? 14'h3b : _GEN_7655;
  wire [13:0] _GEN_7657 = 14'h1de9 == index ? 14'h3b : _GEN_7656;
  wire [13:0] _GEN_7658 = 14'h1dea == index ? 14'h3b : _GEN_7657;
  wire [13:0] _GEN_7659 = 14'h1deb == index ? 14'h3b : _GEN_7658;
  wire [13:0] _GEN_7660 = 14'h1dec == index ? 14'h3b : _GEN_7659;
  wire [13:0] _GEN_7661 = 14'h1ded == index ? 14'h3b : _GEN_7660;
  wire [13:0] _GEN_7662 = 14'h1dee == index ? 14'h3b : _GEN_7661;
  wire [13:0] _GEN_7663 = 14'h1def == index ? 14'h3b : _GEN_7662;
  wire [13:0] _GEN_7664 = 14'h1df0 == index ? 14'h3b : _GEN_7663;
  wire [13:0] _GEN_7665 = 14'h1df1 == index ? 14'h3b : _GEN_7664;
  wire [13:0] _GEN_7666 = 14'h1df2 == index ? 14'h3b : _GEN_7665;
  wire [13:0] _GEN_7667 = 14'h1df3 == index ? 14'h3b : _GEN_7666;
  wire [13:0] _GEN_7668 = 14'h1df4 == index ? 14'h3b : _GEN_7667;
  wire [13:0] _GEN_7669 = 14'h1df5 == index ? 14'h3b : _GEN_7668;
  wire [13:0] _GEN_7670 = 14'h1df6 == index ? 14'h3b : _GEN_7669;
  wire [13:0] _GEN_7671 = 14'h1df7 == index ? 14'h3b : _GEN_7670;
  wire [13:0] _GEN_7672 = 14'h1df8 == index ? 14'h3b : _GEN_7671;
  wire [13:0] _GEN_7673 = 14'h1df9 == index ? 14'h3b : _GEN_7672;
  wire [13:0] _GEN_7674 = 14'h1dfa == index ? 14'h3b : _GEN_7673;
  wire [13:0] _GEN_7675 = 14'h1dfb == index ? 14'h3b : _GEN_7674;
  wire [13:0] _GEN_7676 = 14'h1dfc == index ? 14'h3b : _GEN_7675;
  wire [13:0] _GEN_7677 = 14'h1dfd == index ? 14'h3b : _GEN_7676;
  wire [13:0] _GEN_7678 = 14'h1dfe == index ? 14'h3b : _GEN_7677;
  wire [13:0] _GEN_7679 = 14'h1dff == index ? 14'h3b : _GEN_7678;
  wire [13:0] _GEN_7680 = 14'h1e00 == index ? 14'h0 : _GEN_7679;
  wire [13:0] _GEN_7681 = 14'h1e01 == index ? 14'h1e00 : _GEN_7680;
  wire [13:0] _GEN_7682 = 14'h1e02 == index ? 14'hf00 : _GEN_7681;
  wire [13:0] _GEN_7683 = 14'h1e03 == index ? 14'ha00 : _GEN_7682;
  wire [13:0] _GEN_7684 = 14'h1e04 == index ? 14'h780 : _GEN_7683;
  wire [13:0] _GEN_7685 = 14'h1e05 == index ? 14'h600 : _GEN_7684;
  wire [13:0] _GEN_7686 = 14'h1e06 == index ? 14'h500 : _GEN_7685;
  wire [13:0] _GEN_7687 = 14'h1e07 == index ? 14'h404 : _GEN_7686;
  wire [13:0] _GEN_7688 = 14'h1e08 == index ? 14'h384 : _GEN_7687;
  wire [13:0] _GEN_7689 = 14'h1e09 == index ? 14'h306 : _GEN_7688;
  wire [13:0] _GEN_7690 = 14'h1e0a == index ? 14'h300 : _GEN_7689;
  wire [13:0] _GEN_7691 = 14'h1e0b == index ? 14'h285 : _GEN_7690;
  wire [13:0] _GEN_7692 = 14'h1e0c == index ? 14'h280 : _GEN_7691;
  wire [13:0] _GEN_7693 = 14'h1e0d == index ? 14'h208 : _GEN_7692;
  wire [13:0] _GEN_7694 = 14'h1e0e == index ? 14'h204 : _GEN_7693;
  wire [13:0] _GEN_7695 = 14'h1e0f == index ? 14'h200 : _GEN_7694;
  wire [13:0] _GEN_7696 = 14'h1e10 == index ? 14'h18c : _GEN_7695;
  wire [13:0] _GEN_7697 = 14'h1e11 == index ? 14'h189 : _GEN_7696;
  wire [13:0] _GEN_7698 = 14'h1e12 == index ? 14'h186 : _GEN_7697;
  wire [13:0] _GEN_7699 = 14'h1e13 == index ? 14'h183 : _GEN_7698;
  wire [13:0] _GEN_7700 = 14'h1e14 == index ? 14'h180 : _GEN_7699;
  wire [13:0] _GEN_7701 = 14'h1e15 == index ? 14'h112 : _GEN_7700;
  wire [13:0] _GEN_7702 = 14'h1e16 == index ? 14'h110 : _GEN_7701;
  wire [13:0] _GEN_7703 = 14'h1e17 == index ? 14'h10e : _GEN_7702;
  wire [13:0] _GEN_7704 = 14'h1e18 == index ? 14'h10c : _GEN_7703;
  wire [13:0] _GEN_7705 = 14'h1e19 == index ? 14'h10a : _GEN_7704;
  wire [13:0] _GEN_7706 = 14'h1e1a == index ? 14'h108 : _GEN_7705;
  wire [13:0] _GEN_7707 = 14'h1e1b == index ? 14'h106 : _GEN_7706;
  wire [13:0] _GEN_7708 = 14'h1e1c == index ? 14'h104 : _GEN_7707;
  wire [13:0] _GEN_7709 = 14'h1e1d == index ? 14'h102 : _GEN_7708;
  wire [13:0] _GEN_7710 = 14'h1e1e == index ? 14'h100 : _GEN_7709;
  wire [13:0] _GEN_7711 = 14'h1e1f == index ? 14'h9d : _GEN_7710;
  wire [13:0] _GEN_7712 = 14'h1e20 == index ? 14'h9c : _GEN_7711;
  wire [13:0] _GEN_7713 = 14'h1e21 == index ? 14'h9b : _GEN_7712;
  wire [13:0] _GEN_7714 = 14'h1e22 == index ? 14'h9a : _GEN_7713;
  wire [13:0] _GEN_7715 = 14'h1e23 == index ? 14'h99 : _GEN_7714;
  wire [13:0] _GEN_7716 = 14'h1e24 == index ? 14'h98 : _GEN_7715;
  wire [13:0] _GEN_7717 = 14'h1e25 == index ? 14'h97 : _GEN_7716;
  wire [13:0] _GEN_7718 = 14'h1e26 == index ? 14'h96 : _GEN_7717;
  wire [13:0] _GEN_7719 = 14'h1e27 == index ? 14'h95 : _GEN_7718;
  wire [13:0] _GEN_7720 = 14'h1e28 == index ? 14'h94 : _GEN_7719;
  wire [13:0] _GEN_7721 = 14'h1e29 == index ? 14'h93 : _GEN_7720;
  wire [13:0] _GEN_7722 = 14'h1e2a == index ? 14'h92 : _GEN_7721;
  wire [13:0] _GEN_7723 = 14'h1e2b == index ? 14'h91 : _GEN_7722;
  wire [13:0] _GEN_7724 = 14'h1e2c == index ? 14'h90 : _GEN_7723;
  wire [13:0] _GEN_7725 = 14'h1e2d == index ? 14'h8f : _GEN_7724;
  wire [13:0] _GEN_7726 = 14'h1e2e == index ? 14'h8e : _GEN_7725;
  wire [13:0] _GEN_7727 = 14'h1e2f == index ? 14'h8d : _GEN_7726;
  wire [13:0] _GEN_7728 = 14'h1e30 == index ? 14'h8c : _GEN_7727;
  wire [13:0] _GEN_7729 = 14'h1e31 == index ? 14'h8b : _GEN_7728;
  wire [13:0] _GEN_7730 = 14'h1e32 == index ? 14'h8a : _GEN_7729;
  wire [13:0] _GEN_7731 = 14'h1e33 == index ? 14'h89 : _GEN_7730;
  wire [13:0] _GEN_7732 = 14'h1e34 == index ? 14'h88 : _GEN_7731;
  wire [13:0] _GEN_7733 = 14'h1e35 == index ? 14'h87 : _GEN_7732;
  wire [13:0] _GEN_7734 = 14'h1e36 == index ? 14'h86 : _GEN_7733;
  wire [13:0] _GEN_7735 = 14'h1e37 == index ? 14'h85 : _GEN_7734;
  wire [13:0] _GEN_7736 = 14'h1e38 == index ? 14'h84 : _GEN_7735;
  wire [13:0] _GEN_7737 = 14'h1e39 == index ? 14'h83 : _GEN_7736;
  wire [13:0] _GEN_7738 = 14'h1e3a == index ? 14'h82 : _GEN_7737;
  wire [13:0] _GEN_7739 = 14'h1e3b == index ? 14'h81 : _GEN_7738;
  wire [13:0] _GEN_7740 = 14'h1e3c == index ? 14'h80 : _GEN_7739;
  wire [13:0] _GEN_7741 = 14'h1e3d == index ? 14'h3c : _GEN_7740;
  wire [13:0] _GEN_7742 = 14'h1e3e == index ? 14'h3c : _GEN_7741;
  wire [13:0] _GEN_7743 = 14'h1e3f == index ? 14'h3c : _GEN_7742;
  wire [13:0] _GEN_7744 = 14'h1e40 == index ? 14'h3c : _GEN_7743;
  wire [13:0] _GEN_7745 = 14'h1e41 == index ? 14'h3c : _GEN_7744;
  wire [13:0] _GEN_7746 = 14'h1e42 == index ? 14'h3c : _GEN_7745;
  wire [13:0] _GEN_7747 = 14'h1e43 == index ? 14'h3c : _GEN_7746;
  wire [13:0] _GEN_7748 = 14'h1e44 == index ? 14'h3c : _GEN_7747;
  wire [13:0] _GEN_7749 = 14'h1e45 == index ? 14'h3c : _GEN_7748;
  wire [13:0] _GEN_7750 = 14'h1e46 == index ? 14'h3c : _GEN_7749;
  wire [13:0] _GEN_7751 = 14'h1e47 == index ? 14'h3c : _GEN_7750;
  wire [13:0] _GEN_7752 = 14'h1e48 == index ? 14'h3c : _GEN_7751;
  wire [13:0] _GEN_7753 = 14'h1e49 == index ? 14'h3c : _GEN_7752;
  wire [13:0] _GEN_7754 = 14'h1e4a == index ? 14'h3c : _GEN_7753;
  wire [13:0] _GEN_7755 = 14'h1e4b == index ? 14'h3c : _GEN_7754;
  wire [13:0] _GEN_7756 = 14'h1e4c == index ? 14'h3c : _GEN_7755;
  wire [13:0] _GEN_7757 = 14'h1e4d == index ? 14'h3c : _GEN_7756;
  wire [13:0] _GEN_7758 = 14'h1e4e == index ? 14'h3c : _GEN_7757;
  wire [13:0] _GEN_7759 = 14'h1e4f == index ? 14'h3c : _GEN_7758;
  wire [13:0] _GEN_7760 = 14'h1e50 == index ? 14'h3c : _GEN_7759;
  wire [13:0] _GEN_7761 = 14'h1e51 == index ? 14'h3c : _GEN_7760;
  wire [13:0] _GEN_7762 = 14'h1e52 == index ? 14'h3c : _GEN_7761;
  wire [13:0] _GEN_7763 = 14'h1e53 == index ? 14'h3c : _GEN_7762;
  wire [13:0] _GEN_7764 = 14'h1e54 == index ? 14'h3c : _GEN_7763;
  wire [13:0] _GEN_7765 = 14'h1e55 == index ? 14'h3c : _GEN_7764;
  wire [13:0] _GEN_7766 = 14'h1e56 == index ? 14'h3c : _GEN_7765;
  wire [13:0] _GEN_7767 = 14'h1e57 == index ? 14'h3c : _GEN_7766;
  wire [13:0] _GEN_7768 = 14'h1e58 == index ? 14'h3c : _GEN_7767;
  wire [13:0] _GEN_7769 = 14'h1e59 == index ? 14'h3c : _GEN_7768;
  wire [13:0] _GEN_7770 = 14'h1e5a == index ? 14'h3c : _GEN_7769;
  wire [13:0] _GEN_7771 = 14'h1e5b == index ? 14'h3c : _GEN_7770;
  wire [13:0] _GEN_7772 = 14'h1e5c == index ? 14'h3c : _GEN_7771;
  wire [13:0] _GEN_7773 = 14'h1e5d == index ? 14'h3c : _GEN_7772;
  wire [13:0] _GEN_7774 = 14'h1e5e == index ? 14'h3c : _GEN_7773;
  wire [13:0] _GEN_7775 = 14'h1e5f == index ? 14'h3c : _GEN_7774;
  wire [13:0] _GEN_7776 = 14'h1e60 == index ? 14'h3c : _GEN_7775;
  wire [13:0] _GEN_7777 = 14'h1e61 == index ? 14'h3c : _GEN_7776;
  wire [13:0] _GEN_7778 = 14'h1e62 == index ? 14'h3c : _GEN_7777;
  wire [13:0] _GEN_7779 = 14'h1e63 == index ? 14'h3c : _GEN_7778;
  wire [13:0] _GEN_7780 = 14'h1e64 == index ? 14'h3c : _GEN_7779;
  wire [13:0] _GEN_7781 = 14'h1e65 == index ? 14'h3c : _GEN_7780;
  wire [13:0] _GEN_7782 = 14'h1e66 == index ? 14'h3c : _GEN_7781;
  wire [13:0] _GEN_7783 = 14'h1e67 == index ? 14'h3c : _GEN_7782;
  wire [13:0] _GEN_7784 = 14'h1e68 == index ? 14'h3c : _GEN_7783;
  wire [13:0] _GEN_7785 = 14'h1e69 == index ? 14'h3c : _GEN_7784;
  wire [13:0] _GEN_7786 = 14'h1e6a == index ? 14'h3c : _GEN_7785;
  wire [13:0] _GEN_7787 = 14'h1e6b == index ? 14'h3c : _GEN_7786;
  wire [13:0] _GEN_7788 = 14'h1e6c == index ? 14'h3c : _GEN_7787;
  wire [13:0] _GEN_7789 = 14'h1e6d == index ? 14'h3c : _GEN_7788;
  wire [13:0] _GEN_7790 = 14'h1e6e == index ? 14'h3c : _GEN_7789;
  wire [13:0] _GEN_7791 = 14'h1e6f == index ? 14'h3c : _GEN_7790;
  wire [13:0] _GEN_7792 = 14'h1e70 == index ? 14'h3c : _GEN_7791;
  wire [13:0] _GEN_7793 = 14'h1e71 == index ? 14'h3c : _GEN_7792;
  wire [13:0] _GEN_7794 = 14'h1e72 == index ? 14'h3c : _GEN_7793;
  wire [13:0] _GEN_7795 = 14'h1e73 == index ? 14'h3c : _GEN_7794;
  wire [13:0] _GEN_7796 = 14'h1e74 == index ? 14'h3c : _GEN_7795;
  wire [13:0] _GEN_7797 = 14'h1e75 == index ? 14'h3c : _GEN_7796;
  wire [13:0] _GEN_7798 = 14'h1e76 == index ? 14'h3c : _GEN_7797;
  wire [13:0] _GEN_7799 = 14'h1e77 == index ? 14'h3c : _GEN_7798;
  wire [13:0] _GEN_7800 = 14'h1e78 == index ? 14'h3c : _GEN_7799;
  wire [13:0] _GEN_7801 = 14'h1e79 == index ? 14'h3c : _GEN_7800;
  wire [13:0] _GEN_7802 = 14'h1e7a == index ? 14'h3c : _GEN_7801;
  wire [13:0] _GEN_7803 = 14'h1e7b == index ? 14'h3c : _GEN_7802;
  wire [13:0] _GEN_7804 = 14'h1e7c == index ? 14'h3c : _GEN_7803;
  wire [13:0] _GEN_7805 = 14'h1e7d == index ? 14'h3c : _GEN_7804;
  wire [13:0] _GEN_7806 = 14'h1e7e == index ? 14'h3c : _GEN_7805;
  wire [13:0] _GEN_7807 = 14'h1e7f == index ? 14'h3c : _GEN_7806;
  wire [13:0] _GEN_7808 = 14'h1e80 == index ? 14'h0 : _GEN_7807;
  wire [13:0] _GEN_7809 = 14'h1e81 == index ? 14'h1e80 : _GEN_7808;
  wire [13:0] _GEN_7810 = 14'h1e82 == index ? 14'hf01 : _GEN_7809;
  wire [13:0] _GEN_7811 = 14'h1e83 == index ? 14'ha01 : _GEN_7810;
  wire [13:0] _GEN_7812 = 14'h1e84 == index ? 14'h781 : _GEN_7811;
  wire [13:0] _GEN_7813 = 14'h1e85 == index ? 14'h601 : _GEN_7812;
  wire [13:0] _GEN_7814 = 14'h1e86 == index ? 14'h501 : _GEN_7813;
  wire [13:0] _GEN_7815 = 14'h1e87 == index ? 14'h405 : _GEN_7814;
  wire [13:0] _GEN_7816 = 14'h1e88 == index ? 14'h385 : _GEN_7815;
  wire [13:0] _GEN_7817 = 14'h1e89 == index ? 14'h307 : _GEN_7816;
  wire [13:0] _GEN_7818 = 14'h1e8a == index ? 14'h301 : _GEN_7817;
  wire [13:0] _GEN_7819 = 14'h1e8b == index ? 14'h286 : _GEN_7818;
  wire [13:0] _GEN_7820 = 14'h1e8c == index ? 14'h281 : _GEN_7819;
  wire [13:0] _GEN_7821 = 14'h1e8d == index ? 14'h209 : _GEN_7820;
  wire [13:0] _GEN_7822 = 14'h1e8e == index ? 14'h205 : _GEN_7821;
  wire [13:0] _GEN_7823 = 14'h1e8f == index ? 14'h201 : _GEN_7822;
  wire [13:0] _GEN_7824 = 14'h1e90 == index ? 14'h18d : _GEN_7823;
  wire [13:0] _GEN_7825 = 14'h1e91 == index ? 14'h18a : _GEN_7824;
  wire [13:0] _GEN_7826 = 14'h1e92 == index ? 14'h187 : _GEN_7825;
  wire [13:0] _GEN_7827 = 14'h1e93 == index ? 14'h184 : _GEN_7826;
  wire [13:0] _GEN_7828 = 14'h1e94 == index ? 14'h181 : _GEN_7827;
  wire [13:0] _GEN_7829 = 14'h1e95 == index ? 14'h113 : _GEN_7828;
  wire [13:0] _GEN_7830 = 14'h1e96 == index ? 14'h111 : _GEN_7829;
  wire [13:0] _GEN_7831 = 14'h1e97 == index ? 14'h10f : _GEN_7830;
  wire [13:0] _GEN_7832 = 14'h1e98 == index ? 14'h10d : _GEN_7831;
  wire [13:0] _GEN_7833 = 14'h1e99 == index ? 14'h10b : _GEN_7832;
  wire [13:0] _GEN_7834 = 14'h1e9a == index ? 14'h109 : _GEN_7833;
  wire [13:0] _GEN_7835 = 14'h1e9b == index ? 14'h107 : _GEN_7834;
  wire [13:0] _GEN_7836 = 14'h1e9c == index ? 14'h105 : _GEN_7835;
  wire [13:0] _GEN_7837 = 14'h1e9d == index ? 14'h103 : _GEN_7836;
  wire [13:0] _GEN_7838 = 14'h1e9e == index ? 14'h101 : _GEN_7837;
  wire [13:0] _GEN_7839 = 14'h1e9f == index ? 14'h9e : _GEN_7838;
  wire [13:0] _GEN_7840 = 14'h1ea0 == index ? 14'h9d : _GEN_7839;
  wire [13:0] _GEN_7841 = 14'h1ea1 == index ? 14'h9c : _GEN_7840;
  wire [13:0] _GEN_7842 = 14'h1ea2 == index ? 14'h9b : _GEN_7841;
  wire [13:0] _GEN_7843 = 14'h1ea3 == index ? 14'h9a : _GEN_7842;
  wire [13:0] _GEN_7844 = 14'h1ea4 == index ? 14'h99 : _GEN_7843;
  wire [13:0] _GEN_7845 = 14'h1ea5 == index ? 14'h98 : _GEN_7844;
  wire [13:0] _GEN_7846 = 14'h1ea6 == index ? 14'h97 : _GEN_7845;
  wire [13:0] _GEN_7847 = 14'h1ea7 == index ? 14'h96 : _GEN_7846;
  wire [13:0] _GEN_7848 = 14'h1ea8 == index ? 14'h95 : _GEN_7847;
  wire [13:0] _GEN_7849 = 14'h1ea9 == index ? 14'h94 : _GEN_7848;
  wire [13:0] _GEN_7850 = 14'h1eaa == index ? 14'h93 : _GEN_7849;
  wire [13:0] _GEN_7851 = 14'h1eab == index ? 14'h92 : _GEN_7850;
  wire [13:0] _GEN_7852 = 14'h1eac == index ? 14'h91 : _GEN_7851;
  wire [13:0] _GEN_7853 = 14'h1ead == index ? 14'h90 : _GEN_7852;
  wire [13:0] _GEN_7854 = 14'h1eae == index ? 14'h8f : _GEN_7853;
  wire [13:0] _GEN_7855 = 14'h1eaf == index ? 14'h8e : _GEN_7854;
  wire [13:0] _GEN_7856 = 14'h1eb0 == index ? 14'h8d : _GEN_7855;
  wire [13:0] _GEN_7857 = 14'h1eb1 == index ? 14'h8c : _GEN_7856;
  wire [13:0] _GEN_7858 = 14'h1eb2 == index ? 14'h8b : _GEN_7857;
  wire [13:0] _GEN_7859 = 14'h1eb3 == index ? 14'h8a : _GEN_7858;
  wire [13:0] _GEN_7860 = 14'h1eb4 == index ? 14'h89 : _GEN_7859;
  wire [13:0] _GEN_7861 = 14'h1eb5 == index ? 14'h88 : _GEN_7860;
  wire [13:0] _GEN_7862 = 14'h1eb6 == index ? 14'h87 : _GEN_7861;
  wire [13:0] _GEN_7863 = 14'h1eb7 == index ? 14'h86 : _GEN_7862;
  wire [13:0] _GEN_7864 = 14'h1eb8 == index ? 14'h85 : _GEN_7863;
  wire [13:0] _GEN_7865 = 14'h1eb9 == index ? 14'h84 : _GEN_7864;
  wire [13:0] _GEN_7866 = 14'h1eba == index ? 14'h83 : _GEN_7865;
  wire [13:0] _GEN_7867 = 14'h1ebb == index ? 14'h82 : _GEN_7866;
  wire [13:0] _GEN_7868 = 14'h1ebc == index ? 14'h81 : _GEN_7867;
  wire [13:0] _GEN_7869 = 14'h1ebd == index ? 14'h80 : _GEN_7868;
  wire [13:0] _GEN_7870 = 14'h1ebe == index ? 14'h3d : _GEN_7869;
  wire [13:0] _GEN_7871 = 14'h1ebf == index ? 14'h3d : _GEN_7870;
  wire [13:0] _GEN_7872 = 14'h1ec0 == index ? 14'h3d : _GEN_7871;
  wire [13:0] _GEN_7873 = 14'h1ec1 == index ? 14'h3d : _GEN_7872;
  wire [13:0] _GEN_7874 = 14'h1ec2 == index ? 14'h3d : _GEN_7873;
  wire [13:0] _GEN_7875 = 14'h1ec3 == index ? 14'h3d : _GEN_7874;
  wire [13:0] _GEN_7876 = 14'h1ec4 == index ? 14'h3d : _GEN_7875;
  wire [13:0] _GEN_7877 = 14'h1ec5 == index ? 14'h3d : _GEN_7876;
  wire [13:0] _GEN_7878 = 14'h1ec6 == index ? 14'h3d : _GEN_7877;
  wire [13:0] _GEN_7879 = 14'h1ec7 == index ? 14'h3d : _GEN_7878;
  wire [13:0] _GEN_7880 = 14'h1ec8 == index ? 14'h3d : _GEN_7879;
  wire [13:0] _GEN_7881 = 14'h1ec9 == index ? 14'h3d : _GEN_7880;
  wire [13:0] _GEN_7882 = 14'h1eca == index ? 14'h3d : _GEN_7881;
  wire [13:0] _GEN_7883 = 14'h1ecb == index ? 14'h3d : _GEN_7882;
  wire [13:0] _GEN_7884 = 14'h1ecc == index ? 14'h3d : _GEN_7883;
  wire [13:0] _GEN_7885 = 14'h1ecd == index ? 14'h3d : _GEN_7884;
  wire [13:0] _GEN_7886 = 14'h1ece == index ? 14'h3d : _GEN_7885;
  wire [13:0] _GEN_7887 = 14'h1ecf == index ? 14'h3d : _GEN_7886;
  wire [13:0] _GEN_7888 = 14'h1ed0 == index ? 14'h3d : _GEN_7887;
  wire [13:0] _GEN_7889 = 14'h1ed1 == index ? 14'h3d : _GEN_7888;
  wire [13:0] _GEN_7890 = 14'h1ed2 == index ? 14'h3d : _GEN_7889;
  wire [13:0] _GEN_7891 = 14'h1ed3 == index ? 14'h3d : _GEN_7890;
  wire [13:0] _GEN_7892 = 14'h1ed4 == index ? 14'h3d : _GEN_7891;
  wire [13:0] _GEN_7893 = 14'h1ed5 == index ? 14'h3d : _GEN_7892;
  wire [13:0] _GEN_7894 = 14'h1ed6 == index ? 14'h3d : _GEN_7893;
  wire [13:0] _GEN_7895 = 14'h1ed7 == index ? 14'h3d : _GEN_7894;
  wire [13:0] _GEN_7896 = 14'h1ed8 == index ? 14'h3d : _GEN_7895;
  wire [13:0] _GEN_7897 = 14'h1ed9 == index ? 14'h3d : _GEN_7896;
  wire [13:0] _GEN_7898 = 14'h1eda == index ? 14'h3d : _GEN_7897;
  wire [13:0] _GEN_7899 = 14'h1edb == index ? 14'h3d : _GEN_7898;
  wire [13:0] _GEN_7900 = 14'h1edc == index ? 14'h3d : _GEN_7899;
  wire [13:0] _GEN_7901 = 14'h1edd == index ? 14'h3d : _GEN_7900;
  wire [13:0] _GEN_7902 = 14'h1ede == index ? 14'h3d : _GEN_7901;
  wire [13:0] _GEN_7903 = 14'h1edf == index ? 14'h3d : _GEN_7902;
  wire [13:0] _GEN_7904 = 14'h1ee0 == index ? 14'h3d : _GEN_7903;
  wire [13:0] _GEN_7905 = 14'h1ee1 == index ? 14'h3d : _GEN_7904;
  wire [13:0] _GEN_7906 = 14'h1ee2 == index ? 14'h3d : _GEN_7905;
  wire [13:0] _GEN_7907 = 14'h1ee3 == index ? 14'h3d : _GEN_7906;
  wire [13:0] _GEN_7908 = 14'h1ee4 == index ? 14'h3d : _GEN_7907;
  wire [13:0] _GEN_7909 = 14'h1ee5 == index ? 14'h3d : _GEN_7908;
  wire [13:0] _GEN_7910 = 14'h1ee6 == index ? 14'h3d : _GEN_7909;
  wire [13:0] _GEN_7911 = 14'h1ee7 == index ? 14'h3d : _GEN_7910;
  wire [13:0] _GEN_7912 = 14'h1ee8 == index ? 14'h3d : _GEN_7911;
  wire [13:0] _GEN_7913 = 14'h1ee9 == index ? 14'h3d : _GEN_7912;
  wire [13:0] _GEN_7914 = 14'h1eea == index ? 14'h3d : _GEN_7913;
  wire [13:0] _GEN_7915 = 14'h1eeb == index ? 14'h3d : _GEN_7914;
  wire [13:0] _GEN_7916 = 14'h1eec == index ? 14'h3d : _GEN_7915;
  wire [13:0] _GEN_7917 = 14'h1eed == index ? 14'h3d : _GEN_7916;
  wire [13:0] _GEN_7918 = 14'h1eee == index ? 14'h3d : _GEN_7917;
  wire [13:0] _GEN_7919 = 14'h1eef == index ? 14'h3d : _GEN_7918;
  wire [13:0] _GEN_7920 = 14'h1ef0 == index ? 14'h3d : _GEN_7919;
  wire [13:0] _GEN_7921 = 14'h1ef1 == index ? 14'h3d : _GEN_7920;
  wire [13:0] _GEN_7922 = 14'h1ef2 == index ? 14'h3d : _GEN_7921;
  wire [13:0] _GEN_7923 = 14'h1ef3 == index ? 14'h3d : _GEN_7922;
  wire [13:0] _GEN_7924 = 14'h1ef4 == index ? 14'h3d : _GEN_7923;
  wire [13:0] _GEN_7925 = 14'h1ef5 == index ? 14'h3d : _GEN_7924;
  wire [13:0] _GEN_7926 = 14'h1ef6 == index ? 14'h3d : _GEN_7925;
  wire [13:0] _GEN_7927 = 14'h1ef7 == index ? 14'h3d : _GEN_7926;
  wire [13:0] _GEN_7928 = 14'h1ef8 == index ? 14'h3d : _GEN_7927;
  wire [13:0] _GEN_7929 = 14'h1ef9 == index ? 14'h3d : _GEN_7928;
  wire [13:0] _GEN_7930 = 14'h1efa == index ? 14'h3d : _GEN_7929;
  wire [13:0] _GEN_7931 = 14'h1efb == index ? 14'h3d : _GEN_7930;
  wire [13:0] _GEN_7932 = 14'h1efc == index ? 14'h3d : _GEN_7931;
  wire [13:0] _GEN_7933 = 14'h1efd == index ? 14'h3d : _GEN_7932;
  wire [13:0] _GEN_7934 = 14'h1efe == index ? 14'h3d : _GEN_7933;
  wire [13:0] _GEN_7935 = 14'h1eff == index ? 14'h3d : _GEN_7934;
  wire [13:0] _GEN_7936 = 14'h1f00 == index ? 14'h0 : _GEN_7935;
  wire [13:0] _GEN_7937 = 14'h1f01 == index ? 14'h1f00 : _GEN_7936;
  wire [13:0] _GEN_7938 = 14'h1f02 == index ? 14'hf80 : _GEN_7937;
  wire [13:0] _GEN_7939 = 14'h1f03 == index ? 14'ha02 : _GEN_7938;
  wire [13:0] _GEN_7940 = 14'h1f04 == index ? 14'h782 : _GEN_7939;
  wire [13:0] _GEN_7941 = 14'h1f05 == index ? 14'h602 : _GEN_7940;
  wire [13:0] _GEN_7942 = 14'h1f06 == index ? 14'h502 : _GEN_7941;
  wire [13:0] _GEN_7943 = 14'h1f07 == index ? 14'h406 : _GEN_7942;
  wire [13:0] _GEN_7944 = 14'h1f08 == index ? 14'h386 : _GEN_7943;
  wire [13:0] _GEN_7945 = 14'h1f09 == index ? 14'h308 : _GEN_7944;
  wire [13:0] _GEN_7946 = 14'h1f0a == index ? 14'h302 : _GEN_7945;
  wire [13:0] _GEN_7947 = 14'h1f0b == index ? 14'h287 : _GEN_7946;
  wire [13:0] _GEN_7948 = 14'h1f0c == index ? 14'h282 : _GEN_7947;
  wire [13:0] _GEN_7949 = 14'h1f0d == index ? 14'h20a : _GEN_7948;
  wire [13:0] _GEN_7950 = 14'h1f0e == index ? 14'h206 : _GEN_7949;
  wire [13:0] _GEN_7951 = 14'h1f0f == index ? 14'h202 : _GEN_7950;
  wire [13:0] _GEN_7952 = 14'h1f10 == index ? 14'h18e : _GEN_7951;
  wire [13:0] _GEN_7953 = 14'h1f11 == index ? 14'h18b : _GEN_7952;
  wire [13:0] _GEN_7954 = 14'h1f12 == index ? 14'h188 : _GEN_7953;
  wire [13:0] _GEN_7955 = 14'h1f13 == index ? 14'h185 : _GEN_7954;
  wire [13:0] _GEN_7956 = 14'h1f14 == index ? 14'h182 : _GEN_7955;
  wire [13:0] _GEN_7957 = 14'h1f15 == index ? 14'h114 : _GEN_7956;
  wire [13:0] _GEN_7958 = 14'h1f16 == index ? 14'h112 : _GEN_7957;
  wire [13:0] _GEN_7959 = 14'h1f17 == index ? 14'h110 : _GEN_7958;
  wire [13:0] _GEN_7960 = 14'h1f18 == index ? 14'h10e : _GEN_7959;
  wire [13:0] _GEN_7961 = 14'h1f19 == index ? 14'h10c : _GEN_7960;
  wire [13:0] _GEN_7962 = 14'h1f1a == index ? 14'h10a : _GEN_7961;
  wire [13:0] _GEN_7963 = 14'h1f1b == index ? 14'h108 : _GEN_7962;
  wire [13:0] _GEN_7964 = 14'h1f1c == index ? 14'h106 : _GEN_7963;
  wire [13:0] _GEN_7965 = 14'h1f1d == index ? 14'h104 : _GEN_7964;
  wire [13:0] _GEN_7966 = 14'h1f1e == index ? 14'h102 : _GEN_7965;
  wire [13:0] _GEN_7967 = 14'h1f1f == index ? 14'h100 : _GEN_7966;
  wire [13:0] _GEN_7968 = 14'h1f20 == index ? 14'h9e : _GEN_7967;
  wire [13:0] _GEN_7969 = 14'h1f21 == index ? 14'h9d : _GEN_7968;
  wire [13:0] _GEN_7970 = 14'h1f22 == index ? 14'h9c : _GEN_7969;
  wire [13:0] _GEN_7971 = 14'h1f23 == index ? 14'h9b : _GEN_7970;
  wire [13:0] _GEN_7972 = 14'h1f24 == index ? 14'h9a : _GEN_7971;
  wire [13:0] _GEN_7973 = 14'h1f25 == index ? 14'h99 : _GEN_7972;
  wire [13:0] _GEN_7974 = 14'h1f26 == index ? 14'h98 : _GEN_7973;
  wire [13:0] _GEN_7975 = 14'h1f27 == index ? 14'h97 : _GEN_7974;
  wire [13:0] _GEN_7976 = 14'h1f28 == index ? 14'h96 : _GEN_7975;
  wire [13:0] _GEN_7977 = 14'h1f29 == index ? 14'h95 : _GEN_7976;
  wire [13:0] _GEN_7978 = 14'h1f2a == index ? 14'h94 : _GEN_7977;
  wire [13:0] _GEN_7979 = 14'h1f2b == index ? 14'h93 : _GEN_7978;
  wire [13:0] _GEN_7980 = 14'h1f2c == index ? 14'h92 : _GEN_7979;
  wire [13:0] _GEN_7981 = 14'h1f2d == index ? 14'h91 : _GEN_7980;
  wire [13:0] _GEN_7982 = 14'h1f2e == index ? 14'h90 : _GEN_7981;
  wire [13:0] _GEN_7983 = 14'h1f2f == index ? 14'h8f : _GEN_7982;
  wire [13:0] _GEN_7984 = 14'h1f30 == index ? 14'h8e : _GEN_7983;
  wire [13:0] _GEN_7985 = 14'h1f31 == index ? 14'h8d : _GEN_7984;
  wire [13:0] _GEN_7986 = 14'h1f32 == index ? 14'h8c : _GEN_7985;
  wire [13:0] _GEN_7987 = 14'h1f33 == index ? 14'h8b : _GEN_7986;
  wire [13:0] _GEN_7988 = 14'h1f34 == index ? 14'h8a : _GEN_7987;
  wire [13:0] _GEN_7989 = 14'h1f35 == index ? 14'h89 : _GEN_7988;
  wire [13:0] _GEN_7990 = 14'h1f36 == index ? 14'h88 : _GEN_7989;
  wire [13:0] _GEN_7991 = 14'h1f37 == index ? 14'h87 : _GEN_7990;
  wire [13:0] _GEN_7992 = 14'h1f38 == index ? 14'h86 : _GEN_7991;
  wire [13:0] _GEN_7993 = 14'h1f39 == index ? 14'h85 : _GEN_7992;
  wire [13:0] _GEN_7994 = 14'h1f3a == index ? 14'h84 : _GEN_7993;
  wire [13:0] _GEN_7995 = 14'h1f3b == index ? 14'h83 : _GEN_7994;
  wire [13:0] _GEN_7996 = 14'h1f3c == index ? 14'h82 : _GEN_7995;
  wire [13:0] _GEN_7997 = 14'h1f3d == index ? 14'h81 : _GEN_7996;
  wire [13:0] _GEN_7998 = 14'h1f3e == index ? 14'h80 : _GEN_7997;
  wire [13:0] _GEN_7999 = 14'h1f3f == index ? 14'h3e : _GEN_7998;
  wire [13:0] _GEN_8000 = 14'h1f40 == index ? 14'h3e : _GEN_7999;
  wire [13:0] _GEN_8001 = 14'h1f41 == index ? 14'h3e : _GEN_8000;
  wire [13:0] _GEN_8002 = 14'h1f42 == index ? 14'h3e : _GEN_8001;
  wire [13:0] _GEN_8003 = 14'h1f43 == index ? 14'h3e : _GEN_8002;
  wire [13:0] _GEN_8004 = 14'h1f44 == index ? 14'h3e : _GEN_8003;
  wire [13:0] _GEN_8005 = 14'h1f45 == index ? 14'h3e : _GEN_8004;
  wire [13:0] _GEN_8006 = 14'h1f46 == index ? 14'h3e : _GEN_8005;
  wire [13:0] _GEN_8007 = 14'h1f47 == index ? 14'h3e : _GEN_8006;
  wire [13:0] _GEN_8008 = 14'h1f48 == index ? 14'h3e : _GEN_8007;
  wire [13:0] _GEN_8009 = 14'h1f49 == index ? 14'h3e : _GEN_8008;
  wire [13:0] _GEN_8010 = 14'h1f4a == index ? 14'h3e : _GEN_8009;
  wire [13:0] _GEN_8011 = 14'h1f4b == index ? 14'h3e : _GEN_8010;
  wire [13:0] _GEN_8012 = 14'h1f4c == index ? 14'h3e : _GEN_8011;
  wire [13:0] _GEN_8013 = 14'h1f4d == index ? 14'h3e : _GEN_8012;
  wire [13:0] _GEN_8014 = 14'h1f4e == index ? 14'h3e : _GEN_8013;
  wire [13:0] _GEN_8015 = 14'h1f4f == index ? 14'h3e : _GEN_8014;
  wire [13:0] _GEN_8016 = 14'h1f50 == index ? 14'h3e : _GEN_8015;
  wire [13:0] _GEN_8017 = 14'h1f51 == index ? 14'h3e : _GEN_8016;
  wire [13:0] _GEN_8018 = 14'h1f52 == index ? 14'h3e : _GEN_8017;
  wire [13:0] _GEN_8019 = 14'h1f53 == index ? 14'h3e : _GEN_8018;
  wire [13:0] _GEN_8020 = 14'h1f54 == index ? 14'h3e : _GEN_8019;
  wire [13:0] _GEN_8021 = 14'h1f55 == index ? 14'h3e : _GEN_8020;
  wire [13:0] _GEN_8022 = 14'h1f56 == index ? 14'h3e : _GEN_8021;
  wire [13:0] _GEN_8023 = 14'h1f57 == index ? 14'h3e : _GEN_8022;
  wire [13:0] _GEN_8024 = 14'h1f58 == index ? 14'h3e : _GEN_8023;
  wire [13:0] _GEN_8025 = 14'h1f59 == index ? 14'h3e : _GEN_8024;
  wire [13:0] _GEN_8026 = 14'h1f5a == index ? 14'h3e : _GEN_8025;
  wire [13:0] _GEN_8027 = 14'h1f5b == index ? 14'h3e : _GEN_8026;
  wire [13:0] _GEN_8028 = 14'h1f5c == index ? 14'h3e : _GEN_8027;
  wire [13:0] _GEN_8029 = 14'h1f5d == index ? 14'h3e : _GEN_8028;
  wire [13:0] _GEN_8030 = 14'h1f5e == index ? 14'h3e : _GEN_8029;
  wire [13:0] _GEN_8031 = 14'h1f5f == index ? 14'h3e : _GEN_8030;
  wire [13:0] _GEN_8032 = 14'h1f60 == index ? 14'h3e : _GEN_8031;
  wire [13:0] _GEN_8033 = 14'h1f61 == index ? 14'h3e : _GEN_8032;
  wire [13:0] _GEN_8034 = 14'h1f62 == index ? 14'h3e : _GEN_8033;
  wire [13:0] _GEN_8035 = 14'h1f63 == index ? 14'h3e : _GEN_8034;
  wire [13:0] _GEN_8036 = 14'h1f64 == index ? 14'h3e : _GEN_8035;
  wire [13:0] _GEN_8037 = 14'h1f65 == index ? 14'h3e : _GEN_8036;
  wire [13:0] _GEN_8038 = 14'h1f66 == index ? 14'h3e : _GEN_8037;
  wire [13:0] _GEN_8039 = 14'h1f67 == index ? 14'h3e : _GEN_8038;
  wire [13:0] _GEN_8040 = 14'h1f68 == index ? 14'h3e : _GEN_8039;
  wire [13:0] _GEN_8041 = 14'h1f69 == index ? 14'h3e : _GEN_8040;
  wire [13:0] _GEN_8042 = 14'h1f6a == index ? 14'h3e : _GEN_8041;
  wire [13:0] _GEN_8043 = 14'h1f6b == index ? 14'h3e : _GEN_8042;
  wire [13:0] _GEN_8044 = 14'h1f6c == index ? 14'h3e : _GEN_8043;
  wire [13:0] _GEN_8045 = 14'h1f6d == index ? 14'h3e : _GEN_8044;
  wire [13:0] _GEN_8046 = 14'h1f6e == index ? 14'h3e : _GEN_8045;
  wire [13:0] _GEN_8047 = 14'h1f6f == index ? 14'h3e : _GEN_8046;
  wire [13:0] _GEN_8048 = 14'h1f70 == index ? 14'h3e : _GEN_8047;
  wire [13:0] _GEN_8049 = 14'h1f71 == index ? 14'h3e : _GEN_8048;
  wire [13:0] _GEN_8050 = 14'h1f72 == index ? 14'h3e : _GEN_8049;
  wire [13:0] _GEN_8051 = 14'h1f73 == index ? 14'h3e : _GEN_8050;
  wire [13:0] _GEN_8052 = 14'h1f74 == index ? 14'h3e : _GEN_8051;
  wire [13:0] _GEN_8053 = 14'h1f75 == index ? 14'h3e : _GEN_8052;
  wire [13:0] _GEN_8054 = 14'h1f76 == index ? 14'h3e : _GEN_8053;
  wire [13:0] _GEN_8055 = 14'h1f77 == index ? 14'h3e : _GEN_8054;
  wire [13:0] _GEN_8056 = 14'h1f78 == index ? 14'h3e : _GEN_8055;
  wire [13:0] _GEN_8057 = 14'h1f79 == index ? 14'h3e : _GEN_8056;
  wire [13:0] _GEN_8058 = 14'h1f7a == index ? 14'h3e : _GEN_8057;
  wire [13:0] _GEN_8059 = 14'h1f7b == index ? 14'h3e : _GEN_8058;
  wire [13:0] _GEN_8060 = 14'h1f7c == index ? 14'h3e : _GEN_8059;
  wire [13:0] _GEN_8061 = 14'h1f7d == index ? 14'h3e : _GEN_8060;
  wire [13:0] _GEN_8062 = 14'h1f7e == index ? 14'h3e : _GEN_8061;
  wire [13:0] _GEN_8063 = 14'h1f7f == index ? 14'h3e : _GEN_8062;
  wire [13:0] _GEN_8064 = 14'h1f80 == index ? 14'h0 : _GEN_8063;
  wire [13:0] _GEN_8065 = 14'h1f81 == index ? 14'h1f80 : _GEN_8064;
  wire [13:0] _GEN_8066 = 14'h1f82 == index ? 14'hf81 : _GEN_8065;
  wire [13:0] _GEN_8067 = 14'h1f83 == index ? 14'ha80 : _GEN_8066;
  wire [13:0] _GEN_8068 = 14'h1f84 == index ? 14'h783 : _GEN_8067;
  wire [13:0] _GEN_8069 = 14'h1f85 == index ? 14'h603 : _GEN_8068;
  wire [13:0] _GEN_8070 = 14'h1f86 == index ? 14'h503 : _GEN_8069;
  wire [13:0] _GEN_8071 = 14'h1f87 == index ? 14'h480 : _GEN_8070;
  wire [13:0] _GEN_8072 = 14'h1f88 == index ? 14'h387 : _GEN_8071;
  wire [13:0] _GEN_8073 = 14'h1f89 == index ? 14'h380 : _GEN_8072;
  wire [13:0] _GEN_8074 = 14'h1f8a == index ? 14'h303 : _GEN_8073;
  wire [13:0] _GEN_8075 = 14'h1f8b == index ? 14'h288 : _GEN_8074;
  wire [13:0] _GEN_8076 = 14'h1f8c == index ? 14'h283 : _GEN_8075;
  wire [13:0] _GEN_8077 = 14'h1f8d == index ? 14'h20b : _GEN_8076;
  wire [13:0] _GEN_8078 = 14'h1f8e == index ? 14'h207 : _GEN_8077;
  wire [13:0] _GEN_8079 = 14'h1f8f == index ? 14'h203 : _GEN_8078;
  wire [13:0] _GEN_8080 = 14'h1f90 == index ? 14'h18f : _GEN_8079;
  wire [13:0] _GEN_8081 = 14'h1f91 == index ? 14'h18c : _GEN_8080;
  wire [13:0] _GEN_8082 = 14'h1f92 == index ? 14'h189 : _GEN_8081;
  wire [13:0] _GEN_8083 = 14'h1f93 == index ? 14'h186 : _GEN_8082;
  wire [13:0] _GEN_8084 = 14'h1f94 == index ? 14'h183 : _GEN_8083;
  wire [13:0] _GEN_8085 = 14'h1f95 == index ? 14'h180 : _GEN_8084;
  wire [13:0] _GEN_8086 = 14'h1f96 == index ? 14'h113 : _GEN_8085;
  wire [13:0] _GEN_8087 = 14'h1f97 == index ? 14'h111 : _GEN_8086;
  wire [13:0] _GEN_8088 = 14'h1f98 == index ? 14'h10f : _GEN_8087;
  wire [13:0] _GEN_8089 = 14'h1f99 == index ? 14'h10d : _GEN_8088;
  wire [13:0] _GEN_8090 = 14'h1f9a == index ? 14'h10b : _GEN_8089;
  wire [13:0] _GEN_8091 = 14'h1f9b == index ? 14'h109 : _GEN_8090;
  wire [13:0] _GEN_8092 = 14'h1f9c == index ? 14'h107 : _GEN_8091;
  wire [13:0] _GEN_8093 = 14'h1f9d == index ? 14'h105 : _GEN_8092;
  wire [13:0] _GEN_8094 = 14'h1f9e == index ? 14'h103 : _GEN_8093;
  wire [13:0] _GEN_8095 = 14'h1f9f == index ? 14'h101 : _GEN_8094;
  wire [13:0] _GEN_8096 = 14'h1fa0 == index ? 14'h9f : _GEN_8095;
  wire [13:0] _GEN_8097 = 14'h1fa1 == index ? 14'h9e : _GEN_8096;
  wire [13:0] _GEN_8098 = 14'h1fa2 == index ? 14'h9d : _GEN_8097;
  wire [13:0] _GEN_8099 = 14'h1fa3 == index ? 14'h9c : _GEN_8098;
  wire [13:0] _GEN_8100 = 14'h1fa4 == index ? 14'h9b : _GEN_8099;
  wire [13:0] _GEN_8101 = 14'h1fa5 == index ? 14'h9a : _GEN_8100;
  wire [13:0] _GEN_8102 = 14'h1fa6 == index ? 14'h99 : _GEN_8101;
  wire [13:0] _GEN_8103 = 14'h1fa7 == index ? 14'h98 : _GEN_8102;
  wire [13:0] _GEN_8104 = 14'h1fa8 == index ? 14'h97 : _GEN_8103;
  wire [13:0] _GEN_8105 = 14'h1fa9 == index ? 14'h96 : _GEN_8104;
  wire [13:0] _GEN_8106 = 14'h1faa == index ? 14'h95 : _GEN_8105;
  wire [13:0] _GEN_8107 = 14'h1fab == index ? 14'h94 : _GEN_8106;
  wire [13:0] _GEN_8108 = 14'h1fac == index ? 14'h93 : _GEN_8107;
  wire [13:0] _GEN_8109 = 14'h1fad == index ? 14'h92 : _GEN_8108;
  wire [13:0] _GEN_8110 = 14'h1fae == index ? 14'h91 : _GEN_8109;
  wire [13:0] _GEN_8111 = 14'h1faf == index ? 14'h90 : _GEN_8110;
  wire [13:0] _GEN_8112 = 14'h1fb0 == index ? 14'h8f : _GEN_8111;
  wire [13:0] _GEN_8113 = 14'h1fb1 == index ? 14'h8e : _GEN_8112;
  wire [13:0] _GEN_8114 = 14'h1fb2 == index ? 14'h8d : _GEN_8113;
  wire [13:0] _GEN_8115 = 14'h1fb3 == index ? 14'h8c : _GEN_8114;
  wire [13:0] _GEN_8116 = 14'h1fb4 == index ? 14'h8b : _GEN_8115;
  wire [13:0] _GEN_8117 = 14'h1fb5 == index ? 14'h8a : _GEN_8116;
  wire [13:0] _GEN_8118 = 14'h1fb6 == index ? 14'h89 : _GEN_8117;
  wire [13:0] _GEN_8119 = 14'h1fb7 == index ? 14'h88 : _GEN_8118;
  wire [13:0] _GEN_8120 = 14'h1fb8 == index ? 14'h87 : _GEN_8119;
  wire [13:0] _GEN_8121 = 14'h1fb9 == index ? 14'h86 : _GEN_8120;
  wire [13:0] _GEN_8122 = 14'h1fba == index ? 14'h85 : _GEN_8121;
  wire [13:0] _GEN_8123 = 14'h1fbb == index ? 14'h84 : _GEN_8122;
  wire [13:0] _GEN_8124 = 14'h1fbc == index ? 14'h83 : _GEN_8123;
  wire [13:0] _GEN_8125 = 14'h1fbd == index ? 14'h82 : _GEN_8124;
  wire [13:0] _GEN_8126 = 14'h1fbe == index ? 14'h81 : _GEN_8125;
  wire [13:0] _GEN_8127 = 14'h1fbf == index ? 14'h80 : _GEN_8126;
  wire [13:0] _GEN_8128 = 14'h1fc0 == index ? 14'h3f : _GEN_8127;
  wire [13:0] _GEN_8129 = 14'h1fc1 == index ? 14'h3f : _GEN_8128;
  wire [13:0] _GEN_8130 = 14'h1fc2 == index ? 14'h3f : _GEN_8129;
  wire [13:0] _GEN_8131 = 14'h1fc3 == index ? 14'h3f : _GEN_8130;
  wire [13:0] _GEN_8132 = 14'h1fc4 == index ? 14'h3f : _GEN_8131;
  wire [13:0] _GEN_8133 = 14'h1fc5 == index ? 14'h3f : _GEN_8132;
  wire [13:0] _GEN_8134 = 14'h1fc6 == index ? 14'h3f : _GEN_8133;
  wire [13:0] _GEN_8135 = 14'h1fc7 == index ? 14'h3f : _GEN_8134;
  wire [13:0] _GEN_8136 = 14'h1fc8 == index ? 14'h3f : _GEN_8135;
  wire [13:0] _GEN_8137 = 14'h1fc9 == index ? 14'h3f : _GEN_8136;
  wire [13:0] _GEN_8138 = 14'h1fca == index ? 14'h3f : _GEN_8137;
  wire [13:0] _GEN_8139 = 14'h1fcb == index ? 14'h3f : _GEN_8138;
  wire [13:0] _GEN_8140 = 14'h1fcc == index ? 14'h3f : _GEN_8139;
  wire [13:0] _GEN_8141 = 14'h1fcd == index ? 14'h3f : _GEN_8140;
  wire [13:0] _GEN_8142 = 14'h1fce == index ? 14'h3f : _GEN_8141;
  wire [13:0] _GEN_8143 = 14'h1fcf == index ? 14'h3f : _GEN_8142;
  wire [13:0] _GEN_8144 = 14'h1fd0 == index ? 14'h3f : _GEN_8143;
  wire [13:0] _GEN_8145 = 14'h1fd1 == index ? 14'h3f : _GEN_8144;
  wire [13:0] _GEN_8146 = 14'h1fd2 == index ? 14'h3f : _GEN_8145;
  wire [13:0] _GEN_8147 = 14'h1fd3 == index ? 14'h3f : _GEN_8146;
  wire [13:0] _GEN_8148 = 14'h1fd4 == index ? 14'h3f : _GEN_8147;
  wire [13:0] _GEN_8149 = 14'h1fd5 == index ? 14'h3f : _GEN_8148;
  wire [13:0] _GEN_8150 = 14'h1fd6 == index ? 14'h3f : _GEN_8149;
  wire [13:0] _GEN_8151 = 14'h1fd7 == index ? 14'h3f : _GEN_8150;
  wire [13:0] _GEN_8152 = 14'h1fd8 == index ? 14'h3f : _GEN_8151;
  wire [13:0] _GEN_8153 = 14'h1fd9 == index ? 14'h3f : _GEN_8152;
  wire [13:0] _GEN_8154 = 14'h1fda == index ? 14'h3f : _GEN_8153;
  wire [13:0] _GEN_8155 = 14'h1fdb == index ? 14'h3f : _GEN_8154;
  wire [13:0] _GEN_8156 = 14'h1fdc == index ? 14'h3f : _GEN_8155;
  wire [13:0] _GEN_8157 = 14'h1fdd == index ? 14'h3f : _GEN_8156;
  wire [13:0] _GEN_8158 = 14'h1fde == index ? 14'h3f : _GEN_8157;
  wire [13:0] _GEN_8159 = 14'h1fdf == index ? 14'h3f : _GEN_8158;
  wire [13:0] _GEN_8160 = 14'h1fe0 == index ? 14'h3f : _GEN_8159;
  wire [13:0] _GEN_8161 = 14'h1fe1 == index ? 14'h3f : _GEN_8160;
  wire [13:0] _GEN_8162 = 14'h1fe2 == index ? 14'h3f : _GEN_8161;
  wire [13:0] _GEN_8163 = 14'h1fe3 == index ? 14'h3f : _GEN_8162;
  wire [13:0] _GEN_8164 = 14'h1fe4 == index ? 14'h3f : _GEN_8163;
  wire [13:0] _GEN_8165 = 14'h1fe5 == index ? 14'h3f : _GEN_8164;
  wire [13:0] _GEN_8166 = 14'h1fe6 == index ? 14'h3f : _GEN_8165;
  wire [13:0] _GEN_8167 = 14'h1fe7 == index ? 14'h3f : _GEN_8166;
  wire [13:0] _GEN_8168 = 14'h1fe8 == index ? 14'h3f : _GEN_8167;
  wire [13:0] _GEN_8169 = 14'h1fe9 == index ? 14'h3f : _GEN_8168;
  wire [13:0] _GEN_8170 = 14'h1fea == index ? 14'h3f : _GEN_8169;
  wire [13:0] _GEN_8171 = 14'h1feb == index ? 14'h3f : _GEN_8170;
  wire [13:0] _GEN_8172 = 14'h1fec == index ? 14'h3f : _GEN_8171;
  wire [13:0] _GEN_8173 = 14'h1fed == index ? 14'h3f : _GEN_8172;
  wire [13:0] _GEN_8174 = 14'h1fee == index ? 14'h3f : _GEN_8173;
  wire [13:0] _GEN_8175 = 14'h1fef == index ? 14'h3f : _GEN_8174;
  wire [13:0] _GEN_8176 = 14'h1ff0 == index ? 14'h3f : _GEN_8175;
  wire [13:0] _GEN_8177 = 14'h1ff1 == index ? 14'h3f : _GEN_8176;
  wire [13:0] _GEN_8178 = 14'h1ff2 == index ? 14'h3f : _GEN_8177;
  wire [13:0] _GEN_8179 = 14'h1ff3 == index ? 14'h3f : _GEN_8178;
  wire [13:0] _GEN_8180 = 14'h1ff4 == index ? 14'h3f : _GEN_8179;
  wire [13:0] _GEN_8181 = 14'h1ff5 == index ? 14'h3f : _GEN_8180;
  wire [13:0] _GEN_8182 = 14'h1ff6 == index ? 14'h3f : _GEN_8181;
  wire [13:0] _GEN_8183 = 14'h1ff7 == index ? 14'h3f : _GEN_8182;
  wire [13:0] _GEN_8184 = 14'h1ff8 == index ? 14'h3f : _GEN_8183;
  wire [13:0] _GEN_8185 = 14'h1ff9 == index ? 14'h3f : _GEN_8184;
  wire [13:0] _GEN_8186 = 14'h1ffa == index ? 14'h3f : _GEN_8185;
  wire [13:0] _GEN_8187 = 14'h1ffb == index ? 14'h3f : _GEN_8186;
  wire [13:0] _GEN_8188 = 14'h1ffc == index ? 14'h3f : _GEN_8187;
  wire [13:0] _GEN_8189 = 14'h1ffd == index ? 14'h3f : _GEN_8188;
  wire [13:0] _GEN_8190 = 14'h1ffe == index ? 14'h3f : _GEN_8189;
  wire [13:0] _GEN_8191 = 14'h1fff == index ? 14'h3f : _GEN_8190;
  wire [13:0] _GEN_8192 = 14'h2000 == index ? 14'h0 : _GEN_8191;
  wire [13:0] _GEN_8193 = 14'h2001 == index ? 14'h2000 : _GEN_8192;
  wire [13:0] _GEN_8194 = 14'h2002 == index ? 14'h1000 : _GEN_8193;
  wire [13:0] _GEN_8195 = 14'h2003 == index ? 14'ha81 : _GEN_8194;
  wire [13:0] _GEN_8196 = 14'h2004 == index ? 14'h800 : _GEN_8195;
  wire [13:0] _GEN_8197 = 14'h2005 == index ? 14'h604 : _GEN_8196;
  wire [13:0] _GEN_8198 = 14'h2006 == index ? 14'h504 : _GEN_8197;
  wire [13:0] _GEN_8199 = 14'h2007 == index ? 14'h481 : _GEN_8198;
  wire [13:0] _GEN_8200 = 14'h2008 == index ? 14'h400 : _GEN_8199;
  wire [13:0] _GEN_8201 = 14'h2009 == index ? 14'h381 : _GEN_8200;
  wire [13:0] _GEN_8202 = 14'h200a == index ? 14'h304 : _GEN_8201;
  wire [13:0] _GEN_8203 = 14'h200b == index ? 14'h289 : _GEN_8202;
  wire [13:0] _GEN_8204 = 14'h200c == index ? 14'h284 : _GEN_8203;
  wire [13:0] _GEN_8205 = 14'h200d == index ? 14'h20c : _GEN_8204;
  wire [13:0] _GEN_8206 = 14'h200e == index ? 14'h208 : _GEN_8205;
  wire [13:0] _GEN_8207 = 14'h200f == index ? 14'h204 : _GEN_8206;
  wire [13:0] _GEN_8208 = 14'h2010 == index ? 14'h200 : _GEN_8207;
  wire [13:0] _GEN_8209 = 14'h2011 == index ? 14'h18d : _GEN_8208;
  wire [13:0] _GEN_8210 = 14'h2012 == index ? 14'h18a : _GEN_8209;
  wire [13:0] _GEN_8211 = 14'h2013 == index ? 14'h187 : _GEN_8210;
  wire [13:0] _GEN_8212 = 14'h2014 == index ? 14'h184 : _GEN_8211;
  wire [13:0] _GEN_8213 = 14'h2015 == index ? 14'h181 : _GEN_8212;
  wire [13:0] _GEN_8214 = 14'h2016 == index ? 14'h114 : _GEN_8213;
  wire [13:0] _GEN_8215 = 14'h2017 == index ? 14'h112 : _GEN_8214;
  wire [13:0] _GEN_8216 = 14'h2018 == index ? 14'h110 : _GEN_8215;
  wire [13:0] _GEN_8217 = 14'h2019 == index ? 14'h10e : _GEN_8216;
  wire [13:0] _GEN_8218 = 14'h201a == index ? 14'h10c : _GEN_8217;
  wire [13:0] _GEN_8219 = 14'h201b == index ? 14'h10a : _GEN_8218;
  wire [13:0] _GEN_8220 = 14'h201c == index ? 14'h108 : _GEN_8219;
  wire [13:0] _GEN_8221 = 14'h201d == index ? 14'h106 : _GEN_8220;
  wire [13:0] _GEN_8222 = 14'h201e == index ? 14'h104 : _GEN_8221;
  wire [13:0] _GEN_8223 = 14'h201f == index ? 14'h102 : _GEN_8222;
  wire [13:0] _GEN_8224 = 14'h2020 == index ? 14'h100 : _GEN_8223;
  wire [13:0] _GEN_8225 = 14'h2021 == index ? 14'h9f : _GEN_8224;
  wire [13:0] _GEN_8226 = 14'h2022 == index ? 14'h9e : _GEN_8225;
  wire [13:0] _GEN_8227 = 14'h2023 == index ? 14'h9d : _GEN_8226;
  wire [13:0] _GEN_8228 = 14'h2024 == index ? 14'h9c : _GEN_8227;
  wire [13:0] _GEN_8229 = 14'h2025 == index ? 14'h9b : _GEN_8228;
  wire [13:0] _GEN_8230 = 14'h2026 == index ? 14'h9a : _GEN_8229;
  wire [13:0] _GEN_8231 = 14'h2027 == index ? 14'h99 : _GEN_8230;
  wire [13:0] _GEN_8232 = 14'h2028 == index ? 14'h98 : _GEN_8231;
  wire [13:0] _GEN_8233 = 14'h2029 == index ? 14'h97 : _GEN_8232;
  wire [13:0] _GEN_8234 = 14'h202a == index ? 14'h96 : _GEN_8233;
  wire [13:0] _GEN_8235 = 14'h202b == index ? 14'h95 : _GEN_8234;
  wire [13:0] _GEN_8236 = 14'h202c == index ? 14'h94 : _GEN_8235;
  wire [13:0] _GEN_8237 = 14'h202d == index ? 14'h93 : _GEN_8236;
  wire [13:0] _GEN_8238 = 14'h202e == index ? 14'h92 : _GEN_8237;
  wire [13:0] _GEN_8239 = 14'h202f == index ? 14'h91 : _GEN_8238;
  wire [13:0] _GEN_8240 = 14'h2030 == index ? 14'h90 : _GEN_8239;
  wire [13:0] _GEN_8241 = 14'h2031 == index ? 14'h8f : _GEN_8240;
  wire [13:0] _GEN_8242 = 14'h2032 == index ? 14'h8e : _GEN_8241;
  wire [13:0] _GEN_8243 = 14'h2033 == index ? 14'h8d : _GEN_8242;
  wire [13:0] _GEN_8244 = 14'h2034 == index ? 14'h8c : _GEN_8243;
  wire [13:0] _GEN_8245 = 14'h2035 == index ? 14'h8b : _GEN_8244;
  wire [13:0] _GEN_8246 = 14'h2036 == index ? 14'h8a : _GEN_8245;
  wire [13:0] _GEN_8247 = 14'h2037 == index ? 14'h89 : _GEN_8246;
  wire [13:0] _GEN_8248 = 14'h2038 == index ? 14'h88 : _GEN_8247;
  wire [13:0] _GEN_8249 = 14'h2039 == index ? 14'h87 : _GEN_8248;
  wire [13:0] _GEN_8250 = 14'h203a == index ? 14'h86 : _GEN_8249;
  wire [13:0] _GEN_8251 = 14'h203b == index ? 14'h85 : _GEN_8250;
  wire [13:0] _GEN_8252 = 14'h203c == index ? 14'h84 : _GEN_8251;
  wire [13:0] _GEN_8253 = 14'h203d == index ? 14'h83 : _GEN_8252;
  wire [13:0] _GEN_8254 = 14'h203e == index ? 14'h82 : _GEN_8253;
  wire [13:0] _GEN_8255 = 14'h203f == index ? 14'h81 : _GEN_8254;
  wire [13:0] _GEN_8256 = 14'h2040 == index ? 14'h80 : _GEN_8255;
  wire [13:0] _GEN_8257 = 14'h2041 == index ? 14'h40 : _GEN_8256;
  wire [13:0] _GEN_8258 = 14'h2042 == index ? 14'h40 : _GEN_8257;
  wire [13:0] _GEN_8259 = 14'h2043 == index ? 14'h40 : _GEN_8258;
  wire [13:0] _GEN_8260 = 14'h2044 == index ? 14'h40 : _GEN_8259;
  wire [13:0] _GEN_8261 = 14'h2045 == index ? 14'h40 : _GEN_8260;
  wire [13:0] _GEN_8262 = 14'h2046 == index ? 14'h40 : _GEN_8261;
  wire [13:0] _GEN_8263 = 14'h2047 == index ? 14'h40 : _GEN_8262;
  wire [13:0] _GEN_8264 = 14'h2048 == index ? 14'h40 : _GEN_8263;
  wire [13:0] _GEN_8265 = 14'h2049 == index ? 14'h40 : _GEN_8264;
  wire [13:0] _GEN_8266 = 14'h204a == index ? 14'h40 : _GEN_8265;
  wire [13:0] _GEN_8267 = 14'h204b == index ? 14'h40 : _GEN_8266;
  wire [13:0] _GEN_8268 = 14'h204c == index ? 14'h40 : _GEN_8267;
  wire [13:0] _GEN_8269 = 14'h204d == index ? 14'h40 : _GEN_8268;
  wire [13:0] _GEN_8270 = 14'h204e == index ? 14'h40 : _GEN_8269;
  wire [13:0] _GEN_8271 = 14'h204f == index ? 14'h40 : _GEN_8270;
  wire [13:0] _GEN_8272 = 14'h2050 == index ? 14'h40 : _GEN_8271;
  wire [13:0] _GEN_8273 = 14'h2051 == index ? 14'h40 : _GEN_8272;
  wire [13:0] _GEN_8274 = 14'h2052 == index ? 14'h40 : _GEN_8273;
  wire [13:0] _GEN_8275 = 14'h2053 == index ? 14'h40 : _GEN_8274;
  wire [13:0] _GEN_8276 = 14'h2054 == index ? 14'h40 : _GEN_8275;
  wire [13:0] _GEN_8277 = 14'h2055 == index ? 14'h40 : _GEN_8276;
  wire [13:0] _GEN_8278 = 14'h2056 == index ? 14'h40 : _GEN_8277;
  wire [13:0] _GEN_8279 = 14'h2057 == index ? 14'h40 : _GEN_8278;
  wire [13:0] _GEN_8280 = 14'h2058 == index ? 14'h40 : _GEN_8279;
  wire [13:0] _GEN_8281 = 14'h2059 == index ? 14'h40 : _GEN_8280;
  wire [13:0] _GEN_8282 = 14'h205a == index ? 14'h40 : _GEN_8281;
  wire [13:0] _GEN_8283 = 14'h205b == index ? 14'h40 : _GEN_8282;
  wire [13:0] _GEN_8284 = 14'h205c == index ? 14'h40 : _GEN_8283;
  wire [13:0] _GEN_8285 = 14'h205d == index ? 14'h40 : _GEN_8284;
  wire [13:0] _GEN_8286 = 14'h205e == index ? 14'h40 : _GEN_8285;
  wire [13:0] _GEN_8287 = 14'h205f == index ? 14'h40 : _GEN_8286;
  wire [13:0] _GEN_8288 = 14'h2060 == index ? 14'h40 : _GEN_8287;
  wire [13:0] _GEN_8289 = 14'h2061 == index ? 14'h40 : _GEN_8288;
  wire [13:0] _GEN_8290 = 14'h2062 == index ? 14'h40 : _GEN_8289;
  wire [13:0] _GEN_8291 = 14'h2063 == index ? 14'h40 : _GEN_8290;
  wire [13:0] _GEN_8292 = 14'h2064 == index ? 14'h40 : _GEN_8291;
  wire [13:0] _GEN_8293 = 14'h2065 == index ? 14'h40 : _GEN_8292;
  wire [13:0] _GEN_8294 = 14'h2066 == index ? 14'h40 : _GEN_8293;
  wire [13:0] _GEN_8295 = 14'h2067 == index ? 14'h40 : _GEN_8294;
  wire [13:0] _GEN_8296 = 14'h2068 == index ? 14'h40 : _GEN_8295;
  wire [13:0] _GEN_8297 = 14'h2069 == index ? 14'h40 : _GEN_8296;
  wire [13:0] _GEN_8298 = 14'h206a == index ? 14'h40 : _GEN_8297;
  wire [13:0] _GEN_8299 = 14'h206b == index ? 14'h40 : _GEN_8298;
  wire [13:0] _GEN_8300 = 14'h206c == index ? 14'h40 : _GEN_8299;
  wire [13:0] _GEN_8301 = 14'h206d == index ? 14'h40 : _GEN_8300;
  wire [13:0] _GEN_8302 = 14'h206e == index ? 14'h40 : _GEN_8301;
  wire [13:0] _GEN_8303 = 14'h206f == index ? 14'h40 : _GEN_8302;
  wire [13:0] _GEN_8304 = 14'h2070 == index ? 14'h40 : _GEN_8303;
  wire [13:0] _GEN_8305 = 14'h2071 == index ? 14'h40 : _GEN_8304;
  wire [13:0] _GEN_8306 = 14'h2072 == index ? 14'h40 : _GEN_8305;
  wire [13:0] _GEN_8307 = 14'h2073 == index ? 14'h40 : _GEN_8306;
  wire [13:0] _GEN_8308 = 14'h2074 == index ? 14'h40 : _GEN_8307;
  wire [13:0] _GEN_8309 = 14'h2075 == index ? 14'h40 : _GEN_8308;
  wire [13:0] _GEN_8310 = 14'h2076 == index ? 14'h40 : _GEN_8309;
  wire [13:0] _GEN_8311 = 14'h2077 == index ? 14'h40 : _GEN_8310;
  wire [13:0] _GEN_8312 = 14'h2078 == index ? 14'h40 : _GEN_8311;
  wire [13:0] _GEN_8313 = 14'h2079 == index ? 14'h40 : _GEN_8312;
  wire [13:0] _GEN_8314 = 14'h207a == index ? 14'h40 : _GEN_8313;
  wire [13:0] _GEN_8315 = 14'h207b == index ? 14'h40 : _GEN_8314;
  wire [13:0] _GEN_8316 = 14'h207c == index ? 14'h40 : _GEN_8315;
  wire [13:0] _GEN_8317 = 14'h207d == index ? 14'h40 : _GEN_8316;
  wire [13:0] _GEN_8318 = 14'h207e == index ? 14'h40 : _GEN_8317;
  wire [13:0] _GEN_8319 = 14'h207f == index ? 14'h40 : _GEN_8318;
  wire [13:0] _GEN_8320 = 14'h2080 == index ? 14'h0 : _GEN_8319;
  wire [13:0] _GEN_8321 = 14'h2081 == index ? 14'h2080 : _GEN_8320;
  wire [13:0] _GEN_8322 = 14'h2082 == index ? 14'h1001 : _GEN_8321;
  wire [13:0] _GEN_8323 = 14'h2083 == index ? 14'ha82 : _GEN_8322;
  wire [13:0] _GEN_8324 = 14'h2084 == index ? 14'h801 : _GEN_8323;
  wire [13:0] _GEN_8325 = 14'h2085 == index ? 14'h680 : _GEN_8324;
  wire [13:0] _GEN_8326 = 14'h2086 == index ? 14'h505 : _GEN_8325;
  wire [13:0] _GEN_8327 = 14'h2087 == index ? 14'h482 : _GEN_8326;
  wire [13:0] _GEN_8328 = 14'h2088 == index ? 14'h401 : _GEN_8327;
  wire [13:0] _GEN_8329 = 14'h2089 == index ? 14'h382 : _GEN_8328;
  wire [13:0] _GEN_8330 = 14'h208a == index ? 14'h305 : _GEN_8329;
  wire [13:0] _GEN_8331 = 14'h208b == index ? 14'h28a : _GEN_8330;
  wire [13:0] _GEN_8332 = 14'h208c == index ? 14'h285 : _GEN_8331;
  wire [13:0] _GEN_8333 = 14'h208d == index ? 14'h280 : _GEN_8332;
  wire [13:0] _GEN_8334 = 14'h208e == index ? 14'h209 : _GEN_8333;
  wire [13:0] _GEN_8335 = 14'h208f == index ? 14'h205 : _GEN_8334;
  wire [13:0] _GEN_8336 = 14'h2090 == index ? 14'h201 : _GEN_8335;
  wire [13:0] _GEN_8337 = 14'h2091 == index ? 14'h18e : _GEN_8336;
  wire [13:0] _GEN_8338 = 14'h2092 == index ? 14'h18b : _GEN_8337;
  wire [13:0] _GEN_8339 = 14'h2093 == index ? 14'h188 : _GEN_8338;
  wire [13:0] _GEN_8340 = 14'h2094 == index ? 14'h185 : _GEN_8339;
  wire [13:0] _GEN_8341 = 14'h2095 == index ? 14'h182 : _GEN_8340;
  wire [13:0] _GEN_8342 = 14'h2096 == index ? 14'h115 : _GEN_8341;
  wire [13:0] _GEN_8343 = 14'h2097 == index ? 14'h113 : _GEN_8342;
  wire [13:0] _GEN_8344 = 14'h2098 == index ? 14'h111 : _GEN_8343;
  wire [13:0] _GEN_8345 = 14'h2099 == index ? 14'h10f : _GEN_8344;
  wire [13:0] _GEN_8346 = 14'h209a == index ? 14'h10d : _GEN_8345;
  wire [13:0] _GEN_8347 = 14'h209b == index ? 14'h10b : _GEN_8346;
  wire [13:0] _GEN_8348 = 14'h209c == index ? 14'h109 : _GEN_8347;
  wire [13:0] _GEN_8349 = 14'h209d == index ? 14'h107 : _GEN_8348;
  wire [13:0] _GEN_8350 = 14'h209e == index ? 14'h105 : _GEN_8349;
  wire [13:0] _GEN_8351 = 14'h209f == index ? 14'h103 : _GEN_8350;
  wire [13:0] _GEN_8352 = 14'h20a0 == index ? 14'h101 : _GEN_8351;
  wire [13:0] _GEN_8353 = 14'h20a1 == index ? 14'ha0 : _GEN_8352;
  wire [13:0] _GEN_8354 = 14'h20a2 == index ? 14'h9f : _GEN_8353;
  wire [13:0] _GEN_8355 = 14'h20a3 == index ? 14'h9e : _GEN_8354;
  wire [13:0] _GEN_8356 = 14'h20a4 == index ? 14'h9d : _GEN_8355;
  wire [13:0] _GEN_8357 = 14'h20a5 == index ? 14'h9c : _GEN_8356;
  wire [13:0] _GEN_8358 = 14'h20a6 == index ? 14'h9b : _GEN_8357;
  wire [13:0] _GEN_8359 = 14'h20a7 == index ? 14'h9a : _GEN_8358;
  wire [13:0] _GEN_8360 = 14'h20a8 == index ? 14'h99 : _GEN_8359;
  wire [13:0] _GEN_8361 = 14'h20a9 == index ? 14'h98 : _GEN_8360;
  wire [13:0] _GEN_8362 = 14'h20aa == index ? 14'h97 : _GEN_8361;
  wire [13:0] _GEN_8363 = 14'h20ab == index ? 14'h96 : _GEN_8362;
  wire [13:0] _GEN_8364 = 14'h20ac == index ? 14'h95 : _GEN_8363;
  wire [13:0] _GEN_8365 = 14'h20ad == index ? 14'h94 : _GEN_8364;
  wire [13:0] _GEN_8366 = 14'h20ae == index ? 14'h93 : _GEN_8365;
  wire [13:0] _GEN_8367 = 14'h20af == index ? 14'h92 : _GEN_8366;
  wire [13:0] _GEN_8368 = 14'h20b0 == index ? 14'h91 : _GEN_8367;
  wire [13:0] _GEN_8369 = 14'h20b1 == index ? 14'h90 : _GEN_8368;
  wire [13:0] _GEN_8370 = 14'h20b2 == index ? 14'h8f : _GEN_8369;
  wire [13:0] _GEN_8371 = 14'h20b3 == index ? 14'h8e : _GEN_8370;
  wire [13:0] _GEN_8372 = 14'h20b4 == index ? 14'h8d : _GEN_8371;
  wire [13:0] _GEN_8373 = 14'h20b5 == index ? 14'h8c : _GEN_8372;
  wire [13:0] _GEN_8374 = 14'h20b6 == index ? 14'h8b : _GEN_8373;
  wire [13:0] _GEN_8375 = 14'h20b7 == index ? 14'h8a : _GEN_8374;
  wire [13:0] _GEN_8376 = 14'h20b8 == index ? 14'h89 : _GEN_8375;
  wire [13:0] _GEN_8377 = 14'h20b9 == index ? 14'h88 : _GEN_8376;
  wire [13:0] _GEN_8378 = 14'h20ba == index ? 14'h87 : _GEN_8377;
  wire [13:0] _GEN_8379 = 14'h20bb == index ? 14'h86 : _GEN_8378;
  wire [13:0] _GEN_8380 = 14'h20bc == index ? 14'h85 : _GEN_8379;
  wire [13:0] _GEN_8381 = 14'h20bd == index ? 14'h84 : _GEN_8380;
  wire [13:0] _GEN_8382 = 14'h20be == index ? 14'h83 : _GEN_8381;
  wire [13:0] _GEN_8383 = 14'h20bf == index ? 14'h82 : _GEN_8382;
  wire [13:0] _GEN_8384 = 14'h20c0 == index ? 14'h81 : _GEN_8383;
  wire [13:0] _GEN_8385 = 14'h20c1 == index ? 14'h80 : _GEN_8384;
  wire [13:0] _GEN_8386 = 14'h20c2 == index ? 14'h41 : _GEN_8385;
  wire [13:0] _GEN_8387 = 14'h20c3 == index ? 14'h41 : _GEN_8386;
  wire [13:0] _GEN_8388 = 14'h20c4 == index ? 14'h41 : _GEN_8387;
  wire [13:0] _GEN_8389 = 14'h20c5 == index ? 14'h41 : _GEN_8388;
  wire [13:0] _GEN_8390 = 14'h20c6 == index ? 14'h41 : _GEN_8389;
  wire [13:0] _GEN_8391 = 14'h20c7 == index ? 14'h41 : _GEN_8390;
  wire [13:0] _GEN_8392 = 14'h20c8 == index ? 14'h41 : _GEN_8391;
  wire [13:0] _GEN_8393 = 14'h20c9 == index ? 14'h41 : _GEN_8392;
  wire [13:0] _GEN_8394 = 14'h20ca == index ? 14'h41 : _GEN_8393;
  wire [13:0] _GEN_8395 = 14'h20cb == index ? 14'h41 : _GEN_8394;
  wire [13:0] _GEN_8396 = 14'h20cc == index ? 14'h41 : _GEN_8395;
  wire [13:0] _GEN_8397 = 14'h20cd == index ? 14'h41 : _GEN_8396;
  wire [13:0] _GEN_8398 = 14'h20ce == index ? 14'h41 : _GEN_8397;
  wire [13:0] _GEN_8399 = 14'h20cf == index ? 14'h41 : _GEN_8398;
  wire [13:0] _GEN_8400 = 14'h20d0 == index ? 14'h41 : _GEN_8399;
  wire [13:0] _GEN_8401 = 14'h20d1 == index ? 14'h41 : _GEN_8400;
  wire [13:0] _GEN_8402 = 14'h20d2 == index ? 14'h41 : _GEN_8401;
  wire [13:0] _GEN_8403 = 14'h20d3 == index ? 14'h41 : _GEN_8402;
  wire [13:0] _GEN_8404 = 14'h20d4 == index ? 14'h41 : _GEN_8403;
  wire [13:0] _GEN_8405 = 14'h20d5 == index ? 14'h41 : _GEN_8404;
  wire [13:0] _GEN_8406 = 14'h20d6 == index ? 14'h41 : _GEN_8405;
  wire [13:0] _GEN_8407 = 14'h20d7 == index ? 14'h41 : _GEN_8406;
  wire [13:0] _GEN_8408 = 14'h20d8 == index ? 14'h41 : _GEN_8407;
  wire [13:0] _GEN_8409 = 14'h20d9 == index ? 14'h41 : _GEN_8408;
  wire [13:0] _GEN_8410 = 14'h20da == index ? 14'h41 : _GEN_8409;
  wire [13:0] _GEN_8411 = 14'h20db == index ? 14'h41 : _GEN_8410;
  wire [13:0] _GEN_8412 = 14'h20dc == index ? 14'h41 : _GEN_8411;
  wire [13:0] _GEN_8413 = 14'h20dd == index ? 14'h41 : _GEN_8412;
  wire [13:0] _GEN_8414 = 14'h20de == index ? 14'h41 : _GEN_8413;
  wire [13:0] _GEN_8415 = 14'h20df == index ? 14'h41 : _GEN_8414;
  wire [13:0] _GEN_8416 = 14'h20e0 == index ? 14'h41 : _GEN_8415;
  wire [13:0] _GEN_8417 = 14'h20e1 == index ? 14'h41 : _GEN_8416;
  wire [13:0] _GEN_8418 = 14'h20e2 == index ? 14'h41 : _GEN_8417;
  wire [13:0] _GEN_8419 = 14'h20e3 == index ? 14'h41 : _GEN_8418;
  wire [13:0] _GEN_8420 = 14'h20e4 == index ? 14'h41 : _GEN_8419;
  wire [13:0] _GEN_8421 = 14'h20e5 == index ? 14'h41 : _GEN_8420;
  wire [13:0] _GEN_8422 = 14'h20e6 == index ? 14'h41 : _GEN_8421;
  wire [13:0] _GEN_8423 = 14'h20e7 == index ? 14'h41 : _GEN_8422;
  wire [13:0] _GEN_8424 = 14'h20e8 == index ? 14'h41 : _GEN_8423;
  wire [13:0] _GEN_8425 = 14'h20e9 == index ? 14'h41 : _GEN_8424;
  wire [13:0] _GEN_8426 = 14'h20ea == index ? 14'h41 : _GEN_8425;
  wire [13:0] _GEN_8427 = 14'h20eb == index ? 14'h41 : _GEN_8426;
  wire [13:0] _GEN_8428 = 14'h20ec == index ? 14'h41 : _GEN_8427;
  wire [13:0] _GEN_8429 = 14'h20ed == index ? 14'h41 : _GEN_8428;
  wire [13:0] _GEN_8430 = 14'h20ee == index ? 14'h41 : _GEN_8429;
  wire [13:0] _GEN_8431 = 14'h20ef == index ? 14'h41 : _GEN_8430;
  wire [13:0] _GEN_8432 = 14'h20f0 == index ? 14'h41 : _GEN_8431;
  wire [13:0] _GEN_8433 = 14'h20f1 == index ? 14'h41 : _GEN_8432;
  wire [13:0] _GEN_8434 = 14'h20f2 == index ? 14'h41 : _GEN_8433;
  wire [13:0] _GEN_8435 = 14'h20f3 == index ? 14'h41 : _GEN_8434;
  wire [13:0] _GEN_8436 = 14'h20f4 == index ? 14'h41 : _GEN_8435;
  wire [13:0] _GEN_8437 = 14'h20f5 == index ? 14'h41 : _GEN_8436;
  wire [13:0] _GEN_8438 = 14'h20f6 == index ? 14'h41 : _GEN_8437;
  wire [13:0] _GEN_8439 = 14'h20f7 == index ? 14'h41 : _GEN_8438;
  wire [13:0] _GEN_8440 = 14'h20f8 == index ? 14'h41 : _GEN_8439;
  wire [13:0] _GEN_8441 = 14'h20f9 == index ? 14'h41 : _GEN_8440;
  wire [13:0] _GEN_8442 = 14'h20fa == index ? 14'h41 : _GEN_8441;
  wire [13:0] _GEN_8443 = 14'h20fb == index ? 14'h41 : _GEN_8442;
  wire [13:0] _GEN_8444 = 14'h20fc == index ? 14'h41 : _GEN_8443;
  wire [13:0] _GEN_8445 = 14'h20fd == index ? 14'h41 : _GEN_8444;
  wire [13:0] _GEN_8446 = 14'h20fe == index ? 14'h41 : _GEN_8445;
  wire [13:0] _GEN_8447 = 14'h20ff == index ? 14'h41 : _GEN_8446;
  wire [13:0] _GEN_8448 = 14'h2100 == index ? 14'h0 : _GEN_8447;
  wire [13:0] _GEN_8449 = 14'h2101 == index ? 14'h2100 : _GEN_8448;
  wire [13:0] _GEN_8450 = 14'h2102 == index ? 14'h1080 : _GEN_8449;
  wire [13:0] _GEN_8451 = 14'h2103 == index ? 14'hb00 : _GEN_8450;
  wire [13:0] _GEN_8452 = 14'h2104 == index ? 14'h802 : _GEN_8451;
  wire [13:0] _GEN_8453 = 14'h2105 == index ? 14'h681 : _GEN_8452;
  wire [13:0] _GEN_8454 = 14'h2106 == index ? 14'h580 : _GEN_8453;
  wire [13:0] _GEN_8455 = 14'h2107 == index ? 14'h483 : _GEN_8454;
  wire [13:0] _GEN_8456 = 14'h2108 == index ? 14'h402 : _GEN_8455;
  wire [13:0] _GEN_8457 = 14'h2109 == index ? 14'h383 : _GEN_8456;
  wire [13:0] _GEN_8458 = 14'h210a == index ? 14'h306 : _GEN_8457;
  wire [13:0] _GEN_8459 = 14'h210b == index ? 14'h300 : _GEN_8458;
  wire [13:0] _GEN_8460 = 14'h210c == index ? 14'h286 : _GEN_8459;
  wire [13:0] _GEN_8461 = 14'h210d == index ? 14'h281 : _GEN_8460;
  wire [13:0] _GEN_8462 = 14'h210e == index ? 14'h20a : _GEN_8461;
  wire [13:0] _GEN_8463 = 14'h210f == index ? 14'h206 : _GEN_8462;
  wire [13:0] _GEN_8464 = 14'h2110 == index ? 14'h202 : _GEN_8463;
  wire [13:0] _GEN_8465 = 14'h2111 == index ? 14'h18f : _GEN_8464;
  wire [13:0] _GEN_8466 = 14'h2112 == index ? 14'h18c : _GEN_8465;
  wire [13:0] _GEN_8467 = 14'h2113 == index ? 14'h189 : _GEN_8466;
  wire [13:0] _GEN_8468 = 14'h2114 == index ? 14'h186 : _GEN_8467;
  wire [13:0] _GEN_8469 = 14'h2115 == index ? 14'h183 : _GEN_8468;
  wire [13:0] _GEN_8470 = 14'h2116 == index ? 14'h180 : _GEN_8469;
  wire [13:0] _GEN_8471 = 14'h2117 == index ? 14'h114 : _GEN_8470;
  wire [13:0] _GEN_8472 = 14'h2118 == index ? 14'h112 : _GEN_8471;
  wire [13:0] _GEN_8473 = 14'h2119 == index ? 14'h110 : _GEN_8472;
  wire [13:0] _GEN_8474 = 14'h211a == index ? 14'h10e : _GEN_8473;
  wire [13:0] _GEN_8475 = 14'h211b == index ? 14'h10c : _GEN_8474;
  wire [13:0] _GEN_8476 = 14'h211c == index ? 14'h10a : _GEN_8475;
  wire [13:0] _GEN_8477 = 14'h211d == index ? 14'h108 : _GEN_8476;
  wire [13:0] _GEN_8478 = 14'h211e == index ? 14'h106 : _GEN_8477;
  wire [13:0] _GEN_8479 = 14'h211f == index ? 14'h104 : _GEN_8478;
  wire [13:0] _GEN_8480 = 14'h2120 == index ? 14'h102 : _GEN_8479;
  wire [13:0] _GEN_8481 = 14'h2121 == index ? 14'h100 : _GEN_8480;
  wire [13:0] _GEN_8482 = 14'h2122 == index ? 14'ha0 : _GEN_8481;
  wire [13:0] _GEN_8483 = 14'h2123 == index ? 14'h9f : _GEN_8482;
  wire [13:0] _GEN_8484 = 14'h2124 == index ? 14'h9e : _GEN_8483;
  wire [13:0] _GEN_8485 = 14'h2125 == index ? 14'h9d : _GEN_8484;
  wire [13:0] _GEN_8486 = 14'h2126 == index ? 14'h9c : _GEN_8485;
  wire [13:0] _GEN_8487 = 14'h2127 == index ? 14'h9b : _GEN_8486;
  wire [13:0] _GEN_8488 = 14'h2128 == index ? 14'h9a : _GEN_8487;
  wire [13:0] _GEN_8489 = 14'h2129 == index ? 14'h99 : _GEN_8488;
  wire [13:0] _GEN_8490 = 14'h212a == index ? 14'h98 : _GEN_8489;
  wire [13:0] _GEN_8491 = 14'h212b == index ? 14'h97 : _GEN_8490;
  wire [13:0] _GEN_8492 = 14'h212c == index ? 14'h96 : _GEN_8491;
  wire [13:0] _GEN_8493 = 14'h212d == index ? 14'h95 : _GEN_8492;
  wire [13:0] _GEN_8494 = 14'h212e == index ? 14'h94 : _GEN_8493;
  wire [13:0] _GEN_8495 = 14'h212f == index ? 14'h93 : _GEN_8494;
  wire [13:0] _GEN_8496 = 14'h2130 == index ? 14'h92 : _GEN_8495;
  wire [13:0] _GEN_8497 = 14'h2131 == index ? 14'h91 : _GEN_8496;
  wire [13:0] _GEN_8498 = 14'h2132 == index ? 14'h90 : _GEN_8497;
  wire [13:0] _GEN_8499 = 14'h2133 == index ? 14'h8f : _GEN_8498;
  wire [13:0] _GEN_8500 = 14'h2134 == index ? 14'h8e : _GEN_8499;
  wire [13:0] _GEN_8501 = 14'h2135 == index ? 14'h8d : _GEN_8500;
  wire [13:0] _GEN_8502 = 14'h2136 == index ? 14'h8c : _GEN_8501;
  wire [13:0] _GEN_8503 = 14'h2137 == index ? 14'h8b : _GEN_8502;
  wire [13:0] _GEN_8504 = 14'h2138 == index ? 14'h8a : _GEN_8503;
  wire [13:0] _GEN_8505 = 14'h2139 == index ? 14'h89 : _GEN_8504;
  wire [13:0] _GEN_8506 = 14'h213a == index ? 14'h88 : _GEN_8505;
  wire [13:0] _GEN_8507 = 14'h213b == index ? 14'h87 : _GEN_8506;
  wire [13:0] _GEN_8508 = 14'h213c == index ? 14'h86 : _GEN_8507;
  wire [13:0] _GEN_8509 = 14'h213d == index ? 14'h85 : _GEN_8508;
  wire [13:0] _GEN_8510 = 14'h213e == index ? 14'h84 : _GEN_8509;
  wire [13:0] _GEN_8511 = 14'h213f == index ? 14'h83 : _GEN_8510;
  wire [13:0] _GEN_8512 = 14'h2140 == index ? 14'h82 : _GEN_8511;
  wire [13:0] _GEN_8513 = 14'h2141 == index ? 14'h81 : _GEN_8512;
  wire [13:0] _GEN_8514 = 14'h2142 == index ? 14'h80 : _GEN_8513;
  wire [13:0] _GEN_8515 = 14'h2143 == index ? 14'h42 : _GEN_8514;
  wire [13:0] _GEN_8516 = 14'h2144 == index ? 14'h42 : _GEN_8515;
  wire [13:0] _GEN_8517 = 14'h2145 == index ? 14'h42 : _GEN_8516;
  wire [13:0] _GEN_8518 = 14'h2146 == index ? 14'h42 : _GEN_8517;
  wire [13:0] _GEN_8519 = 14'h2147 == index ? 14'h42 : _GEN_8518;
  wire [13:0] _GEN_8520 = 14'h2148 == index ? 14'h42 : _GEN_8519;
  wire [13:0] _GEN_8521 = 14'h2149 == index ? 14'h42 : _GEN_8520;
  wire [13:0] _GEN_8522 = 14'h214a == index ? 14'h42 : _GEN_8521;
  wire [13:0] _GEN_8523 = 14'h214b == index ? 14'h42 : _GEN_8522;
  wire [13:0] _GEN_8524 = 14'h214c == index ? 14'h42 : _GEN_8523;
  wire [13:0] _GEN_8525 = 14'h214d == index ? 14'h42 : _GEN_8524;
  wire [13:0] _GEN_8526 = 14'h214e == index ? 14'h42 : _GEN_8525;
  wire [13:0] _GEN_8527 = 14'h214f == index ? 14'h42 : _GEN_8526;
  wire [13:0] _GEN_8528 = 14'h2150 == index ? 14'h42 : _GEN_8527;
  wire [13:0] _GEN_8529 = 14'h2151 == index ? 14'h42 : _GEN_8528;
  wire [13:0] _GEN_8530 = 14'h2152 == index ? 14'h42 : _GEN_8529;
  wire [13:0] _GEN_8531 = 14'h2153 == index ? 14'h42 : _GEN_8530;
  wire [13:0] _GEN_8532 = 14'h2154 == index ? 14'h42 : _GEN_8531;
  wire [13:0] _GEN_8533 = 14'h2155 == index ? 14'h42 : _GEN_8532;
  wire [13:0] _GEN_8534 = 14'h2156 == index ? 14'h42 : _GEN_8533;
  wire [13:0] _GEN_8535 = 14'h2157 == index ? 14'h42 : _GEN_8534;
  wire [13:0] _GEN_8536 = 14'h2158 == index ? 14'h42 : _GEN_8535;
  wire [13:0] _GEN_8537 = 14'h2159 == index ? 14'h42 : _GEN_8536;
  wire [13:0] _GEN_8538 = 14'h215a == index ? 14'h42 : _GEN_8537;
  wire [13:0] _GEN_8539 = 14'h215b == index ? 14'h42 : _GEN_8538;
  wire [13:0] _GEN_8540 = 14'h215c == index ? 14'h42 : _GEN_8539;
  wire [13:0] _GEN_8541 = 14'h215d == index ? 14'h42 : _GEN_8540;
  wire [13:0] _GEN_8542 = 14'h215e == index ? 14'h42 : _GEN_8541;
  wire [13:0] _GEN_8543 = 14'h215f == index ? 14'h42 : _GEN_8542;
  wire [13:0] _GEN_8544 = 14'h2160 == index ? 14'h42 : _GEN_8543;
  wire [13:0] _GEN_8545 = 14'h2161 == index ? 14'h42 : _GEN_8544;
  wire [13:0] _GEN_8546 = 14'h2162 == index ? 14'h42 : _GEN_8545;
  wire [13:0] _GEN_8547 = 14'h2163 == index ? 14'h42 : _GEN_8546;
  wire [13:0] _GEN_8548 = 14'h2164 == index ? 14'h42 : _GEN_8547;
  wire [13:0] _GEN_8549 = 14'h2165 == index ? 14'h42 : _GEN_8548;
  wire [13:0] _GEN_8550 = 14'h2166 == index ? 14'h42 : _GEN_8549;
  wire [13:0] _GEN_8551 = 14'h2167 == index ? 14'h42 : _GEN_8550;
  wire [13:0] _GEN_8552 = 14'h2168 == index ? 14'h42 : _GEN_8551;
  wire [13:0] _GEN_8553 = 14'h2169 == index ? 14'h42 : _GEN_8552;
  wire [13:0] _GEN_8554 = 14'h216a == index ? 14'h42 : _GEN_8553;
  wire [13:0] _GEN_8555 = 14'h216b == index ? 14'h42 : _GEN_8554;
  wire [13:0] _GEN_8556 = 14'h216c == index ? 14'h42 : _GEN_8555;
  wire [13:0] _GEN_8557 = 14'h216d == index ? 14'h42 : _GEN_8556;
  wire [13:0] _GEN_8558 = 14'h216e == index ? 14'h42 : _GEN_8557;
  wire [13:0] _GEN_8559 = 14'h216f == index ? 14'h42 : _GEN_8558;
  wire [13:0] _GEN_8560 = 14'h2170 == index ? 14'h42 : _GEN_8559;
  wire [13:0] _GEN_8561 = 14'h2171 == index ? 14'h42 : _GEN_8560;
  wire [13:0] _GEN_8562 = 14'h2172 == index ? 14'h42 : _GEN_8561;
  wire [13:0] _GEN_8563 = 14'h2173 == index ? 14'h42 : _GEN_8562;
  wire [13:0] _GEN_8564 = 14'h2174 == index ? 14'h42 : _GEN_8563;
  wire [13:0] _GEN_8565 = 14'h2175 == index ? 14'h42 : _GEN_8564;
  wire [13:0] _GEN_8566 = 14'h2176 == index ? 14'h42 : _GEN_8565;
  wire [13:0] _GEN_8567 = 14'h2177 == index ? 14'h42 : _GEN_8566;
  wire [13:0] _GEN_8568 = 14'h2178 == index ? 14'h42 : _GEN_8567;
  wire [13:0] _GEN_8569 = 14'h2179 == index ? 14'h42 : _GEN_8568;
  wire [13:0] _GEN_8570 = 14'h217a == index ? 14'h42 : _GEN_8569;
  wire [13:0] _GEN_8571 = 14'h217b == index ? 14'h42 : _GEN_8570;
  wire [13:0] _GEN_8572 = 14'h217c == index ? 14'h42 : _GEN_8571;
  wire [13:0] _GEN_8573 = 14'h217d == index ? 14'h42 : _GEN_8572;
  wire [13:0] _GEN_8574 = 14'h217e == index ? 14'h42 : _GEN_8573;
  wire [13:0] _GEN_8575 = 14'h217f == index ? 14'h42 : _GEN_8574;
  wire [13:0] _GEN_8576 = 14'h2180 == index ? 14'h0 : _GEN_8575;
  wire [13:0] _GEN_8577 = 14'h2181 == index ? 14'h2180 : _GEN_8576;
  wire [13:0] _GEN_8578 = 14'h2182 == index ? 14'h1081 : _GEN_8577;
  wire [13:0] _GEN_8579 = 14'h2183 == index ? 14'hb01 : _GEN_8578;
  wire [13:0] _GEN_8580 = 14'h2184 == index ? 14'h803 : _GEN_8579;
  wire [13:0] _GEN_8581 = 14'h2185 == index ? 14'h682 : _GEN_8580;
  wire [13:0] _GEN_8582 = 14'h2186 == index ? 14'h581 : _GEN_8581;
  wire [13:0] _GEN_8583 = 14'h2187 == index ? 14'h484 : _GEN_8582;
  wire [13:0] _GEN_8584 = 14'h2188 == index ? 14'h403 : _GEN_8583;
  wire [13:0] _GEN_8585 = 14'h2189 == index ? 14'h384 : _GEN_8584;
  wire [13:0] _GEN_8586 = 14'h218a == index ? 14'h307 : _GEN_8585;
  wire [13:0] _GEN_8587 = 14'h218b == index ? 14'h301 : _GEN_8586;
  wire [13:0] _GEN_8588 = 14'h218c == index ? 14'h287 : _GEN_8587;
  wire [13:0] _GEN_8589 = 14'h218d == index ? 14'h282 : _GEN_8588;
  wire [13:0] _GEN_8590 = 14'h218e == index ? 14'h20b : _GEN_8589;
  wire [13:0] _GEN_8591 = 14'h218f == index ? 14'h207 : _GEN_8590;
  wire [13:0] _GEN_8592 = 14'h2190 == index ? 14'h203 : _GEN_8591;
  wire [13:0] _GEN_8593 = 14'h2191 == index ? 14'h190 : _GEN_8592;
  wire [13:0] _GEN_8594 = 14'h2192 == index ? 14'h18d : _GEN_8593;
  wire [13:0] _GEN_8595 = 14'h2193 == index ? 14'h18a : _GEN_8594;
  wire [13:0] _GEN_8596 = 14'h2194 == index ? 14'h187 : _GEN_8595;
  wire [13:0] _GEN_8597 = 14'h2195 == index ? 14'h184 : _GEN_8596;
  wire [13:0] _GEN_8598 = 14'h2196 == index ? 14'h181 : _GEN_8597;
  wire [13:0] _GEN_8599 = 14'h2197 == index ? 14'h115 : _GEN_8598;
  wire [13:0] _GEN_8600 = 14'h2198 == index ? 14'h113 : _GEN_8599;
  wire [13:0] _GEN_8601 = 14'h2199 == index ? 14'h111 : _GEN_8600;
  wire [13:0] _GEN_8602 = 14'h219a == index ? 14'h10f : _GEN_8601;
  wire [13:0] _GEN_8603 = 14'h219b == index ? 14'h10d : _GEN_8602;
  wire [13:0] _GEN_8604 = 14'h219c == index ? 14'h10b : _GEN_8603;
  wire [13:0] _GEN_8605 = 14'h219d == index ? 14'h109 : _GEN_8604;
  wire [13:0] _GEN_8606 = 14'h219e == index ? 14'h107 : _GEN_8605;
  wire [13:0] _GEN_8607 = 14'h219f == index ? 14'h105 : _GEN_8606;
  wire [13:0] _GEN_8608 = 14'h21a0 == index ? 14'h103 : _GEN_8607;
  wire [13:0] _GEN_8609 = 14'h21a1 == index ? 14'h101 : _GEN_8608;
  wire [13:0] _GEN_8610 = 14'h21a2 == index ? 14'ha1 : _GEN_8609;
  wire [13:0] _GEN_8611 = 14'h21a3 == index ? 14'ha0 : _GEN_8610;
  wire [13:0] _GEN_8612 = 14'h21a4 == index ? 14'h9f : _GEN_8611;
  wire [13:0] _GEN_8613 = 14'h21a5 == index ? 14'h9e : _GEN_8612;
  wire [13:0] _GEN_8614 = 14'h21a6 == index ? 14'h9d : _GEN_8613;
  wire [13:0] _GEN_8615 = 14'h21a7 == index ? 14'h9c : _GEN_8614;
  wire [13:0] _GEN_8616 = 14'h21a8 == index ? 14'h9b : _GEN_8615;
  wire [13:0] _GEN_8617 = 14'h21a9 == index ? 14'h9a : _GEN_8616;
  wire [13:0] _GEN_8618 = 14'h21aa == index ? 14'h99 : _GEN_8617;
  wire [13:0] _GEN_8619 = 14'h21ab == index ? 14'h98 : _GEN_8618;
  wire [13:0] _GEN_8620 = 14'h21ac == index ? 14'h97 : _GEN_8619;
  wire [13:0] _GEN_8621 = 14'h21ad == index ? 14'h96 : _GEN_8620;
  wire [13:0] _GEN_8622 = 14'h21ae == index ? 14'h95 : _GEN_8621;
  wire [13:0] _GEN_8623 = 14'h21af == index ? 14'h94 : _GEN_8622;
  wire [13:0] _GEN_8624 = 14'h21b0 == index ? 14'h93 : _GEN_8623;
  wire [13:0] _GEN_8625 = 14'h21b1 == index ? 14'h92 : _GEN_8624;
  wire [13:0] _GEN_8626 = 14'h21b2 == index ? 14'h91 : _GEN_8625;
  wire [13:0] _GEN_8627 = 14'h21b3 == index ? 14'h90 : _GEN_8626;
  wire [13:0] _GEN_8628 = 14'h21b4 == index ? 14'h8f : _GEN_8627;
  wire [13:0] _GEN_8629 = 14'h21b5 == index ? 14'h8e : _GEN_8628;
  wire [13:0] _GEN_8630 = 14'h21b6 == index ? 14'h8d : _GEN_8629;
  wire [13:0] _GEN_8631 = 14'h21b7 == index ? 14'h8c : _GEN_8630;
  wire [13:0] _GEN_8632 = 14'h21b8 == index ? 14'h8b : _GEN_8631;
  wire [13:0] _GEN_8633 = 14'h21b9 == index ? 14'h8a : _GEN_8632;
  wire [13:0] _GEN_8634 = 14'h21ba == index ? 14'h89 : _GEN_8633;
  wire [13:0] _GEN_8635 = 14'h21bb == index ? 14'h88 : _GEN_8634;
  wire [13:0] _GEN_8636 = 14'h21bc == index ? 14'h87 : _GEN_8635;
  wire [13:0] _GEN_8637 = 14'h21bd == index ? 14'h86 : _GEN_8636;
  wire [13:0] _GEN_8638 = 14'h21be == index ? 14'h85 : _GEN_8637;
  wire [13:0] _GEN_8639 = 14'h21bf == index ? 14'h84 : _GEN_8638;
  wire [13:0] _GEN_8640 = 14'h21c0 == index ? 14'h83 : _GEN_8639;
  wire [13:0] _GEN_8641 = 14'h21c1 == index ? 14'h82 : _GEN_8640;
  wire [13:0] _GEN_8642 = 14'h21c2 == index ? 14'h81 : _GEN_8641;
  wire [13:0] _GEN_8643 = 14'h21c3 == index ? 14'h80 : _GEN_8642;
  wire [13:0] _GEN_8644 = 14'h21c4 == index ? 14'h43 : _GEN_8643;
  wire [13:0] _GEN_8645 = 14'h21c5 == index ? 14'h43 : _GEN_8644;
  wire [13:0] _GEN_8646 = 14'h21c6 == index ? 14'h43 : _GEN_8645;
  wire [13:0] _GEN_8647 = 14'h21c7 == index ? 14'h43 : _GEN_8646;
  wire [13:0] _GEN_8648 = 14'h21c8 == index ? 14'h43 : _GEN_8647;
  wire [13:0] _GEN_8649 = 14'h21c9 == index ? 14'h43 : _GEN_8648;
  wire [13:0] _GEN_8650 = 14'h21ca == index ? 14'h43 : _GEN_8649;
  wire [13:0] _GEN_8651 = 14'h21cb == index ? 14'h43 : _GEN_8650;
  wire [13:0] _GEN_8652 = 14'h21cc == index ? 14'h43 : _GEN_8651;
  wire [13:0] _GEN_8653 = 14'h21cd == index ? 14'h43 : _GEN_8652;
  wire [13:0] _GEN_8654 = 14'h21ce == index ? 14'h43 : _GEN_8653;
  wire [13:0] _GEN_8655 = 14'h21cf == index ? 14'h43 : _GEN_8654;
  wire [13:0] _GEN_8656 = 14'h21d0 == index ? 14'h43 : _GEN_8655;
  wire [13:0] _GEN_8657 = 14'h21d1 == index ? 14'h43 : _GEN_8656;
  wire [13:0] _GEN_8658 = 14'h21d2 == index ? 14'h43 : _GEN_8657;
  wire [13:0] _GEN_8659 = 14'h21d3 == index ? 14'h43 : _GEN_8658;
  wire [13:0] _GEN_8660 = 14'h21d4 == index ? 14'h43 : _GEN_8659;
  wire [13:0] _GEN_8661 = 14'h21d5 == index ? 14'h43 : _GEN_8660;
  wire [13:0] _GEN_8662 = 14'h21d6 == index ? 14'h43 : _GEN_8661;
  wire [13:0] _GEN_8663 = 14'h21d7 == index ? 14'h43 : _GEN_8662;
  wire [13:0] _GEN_8664 = 14'h21d8 == index ? 14'h43 : _GEN_8663;
  wire [13:0] _GEN_8665 = 14'h21d9 == index ? 14'h43 : _GEN_8664;
  wire [13:0] _GEN_8666 = 14'h21da == index ? 14'h43 : _GEN_8665;
  wire [13:0] _GEN_8667 = 14'h21db == index ? 14'h43 : _GEN_8666;
  wire [13:0] _GEN_8668 = 14'h21dc == index ? 14'h43 : _GEN_8667;
  wire [13:0] _GEN_8669 = 14'h21dd == index ? 14'h43 : _GEN_8668;
  wire [13:0] _GEN_8670 = 14'h21de == index ? 14'h43 : _GEN_8669;
  wire [13:0] _GEN_8671 = 14'h21df == index ? 14'h43 : _GEN_8670;
  wire [13:0] _GEN_8672 = 14'h21e0 == index ? 14'h43 : _GEN_8671;
  wire [13:0] _GEN_8673 = 14'h21e1 == index ? 14'h43 : _GEN_8672;
  wire [13:0] _GEN_8674 = 14'h21e2 == index ? 14'h43 : _GEN_8673;
  wire [13:0] _GEN_8675 = 14'h21e3 == index ? 14'h43 : _GEN_8674;
  wire [13:0] _GEN_8676 = 14'h21e4 == index ? 14'h43 : _GEN_8675;
  wire [13:0] _GEN_8677 = 14'h21e5 == index ? 14'h43 : _GEN_8676;
  wire [13:0] _GEN_8678 = 14'h21e6 == index ? 14'h43 : _GEN_8677;
  wire [13:0] _GEN_8679 = 14'h21e7 == index ? 14'h43 : _GEN_8678;
  wire [13:0] _GEN_8680 = 14'h21e8 == index ? 14'h43 : _GEN_8679;
  wire [13:0] _GEN_8681 = 14'h21e9 == index ? 14'h43 : _GEN_8680;
  wire [13:0] _GEN_8682 = 14'h21ea == index ? 14'h43 : _GEN_8681;
  wire [13:0] _GEN_8683 = 14'h21eb == index ? 14'h43 : _GEN_8682;
  wire [13:0] _GEN_8684 = 14'h21ec == index ? 14'h43 : _GEN_8683;
  wire [13:0] _GEN_8685 = 14'h21ed == index ? 14'h43 : _GEN_8684;
  wire [13:0] _GEN_8686 = 14'h21ee == index ? 14'h43 : _GEN_8685;
  wire [13:0] _GEN_8687 = 14'h21ef == index ? 14'h43 : _GEN_8686;
  wire [13:0] _GEN_8688 = 14'h21f0 == index ? 14'h43 : _GEN_8687;
  wire [13:0] _GEN_8689 = 14'h21f1 == index ? 14'h43 : _GEN_8688;
  wire [13:0] _GEN_8690 = 14'h21f2 == index ? 14'h43 : _GEN_8689;
  wire [13:0] _GEN_8691 = 14'h21f3 == index ? 14'h43 : _GEN_8690;
  wire [13:0] _GEN_8692 = 14'h21f4 == index ? 14'h43 : _GEN_8691;
  wire [13:0] _GEN_8693 = 14'h21f5 == index ? 14'h43 : _GEN_8692;
  wire [13:0] _GEN_8694 = 14'h21f6 == index ? 14'h43 : _GEN_8693;
  wire [13:0] _GEN_8695 = 14'h21f7 == index ? 14'h43 : _GEN_8694;
  wire [13:0] _GEN_8696 = 14'h21f8 == index ? 14'h43 : _GEN_8695;
  wire [13:0] _GEN_8697 = 14'h21f9 == index ? 14'h43 : _GEN_8696;
  wire [13:0] _GEN_8698 = 14'h21fa == index ? 14'h43 : _GEN_8697;
  wire [13:0] _GEN_8699 = 14'h21fb == index ? 14'h43 : _GEN_8698;
  wire [13:0] _GEN_8700 = 14'h21fc == index ? 14'h43 : _GEN_8699;
  wire [13:0] _GEN_8701 = 14'h21fd == index ? 14'h43 : _GEN_8700;
  wire [13:0] _GEN_8702 = 14'h21fe == index ? 14'h43 : _GEN_8701;
  wire [13:0] _GEN_8703 = 14'h21ff == index ? 14'h43 : _GEN_8702;
  wire [13:0] _GEN_8704 = 14'h2200 == index ? 14'h0 : _GEN_8703;
  wire [13:0] _GEN_8705 = 14'h2201 == index ? 14'h2200 : _GEN_8704;
  wire [13:0] _GEN_8706 = 14'h2202 == index ? 14'h1100 : _GEN_8705;
  wire [13:0] _GEN_8707 = 14'h2203 == index ? 14'hb02 : _GEN_8706;
  wire [13:0] _GEN_8708 = 14'h2204 == index ? 14'h880 : _GEN_8707;
  wire [13:0] _GEN_8709 = 14'h2205 == index ? 14'h683 : _GEN_8708;
  wire [13:0] _GEN_8710 = 14'h2206 == index ? 14'h582 : _GEN_8709;
  wire [13:0] _GEN_8711 = 14'h2207 == index ? 14'h485 : _GEN_8710;
  wire [13:0] _GEN_8712 = 14'h2208 == index ? 14'h404 : _GEN_8711;
  wire [13:0] _GEN_8713 = 14'h2209 == index ? 14'h385 : _GEN_8712;
  wire [13:0] _GEN_8714 = 14'h220a == index ? 14'h308 : _GEN_8713;
  wire [13:0] _GEN_8715 = 14'h220b == index ? 14'h302 : _GEN_8714;
  wire [13:0] _GEN_8716 = 14'h220c == index ? 14'h288 : _GEN_8715;
  wire [13:0] _GEN_8717 = 14'h220d == index ? 14'h283 : _GEN_8716;
  wire [13:0] _GEN_8718 = 14'h220e == index ? 14'h20c : _GEN_8717;
  wire [13:0] _GEN_8719 = 14'h220f == index ? 14'h208 : _GEN_8718;
  wire [13:0] _GEN_8720 = 14'h2210 == index ? 14'h204 : _GEN_8719;
  wire [13:0] _GEN_8721 = 14'h2211 == index ? 14'h200 : _GEN_8720;
  wire [13:0] _GEN_8722 = 14'h2212 == index ? 14'h18e : _GEN_8721;
  wire [13:0] _GEN_8723 = 14'h2213 == index ? 14'h18b : _GEN_8722;
  wire [13:0] _GEN_8724 = 14'h2214 == index ? 14'h188 : _GEN_8723;
  wire [13:0] _GEN_8725 = 14'h2215 == index ? 14'h185 : _GEN_8724;
  wire [13:0] _GEN_8726 = 14'h2216 == index ? 14'h182 : _GEN_8725;
  wire [13:0] _GEN_8727 = 14'h2217 == index ? 14'h116 : _GEN_8726;
  wire [13:0] _GEN_8728 = 14'h2218 == index ? 14'h114 : _GEN_8727;
  wire [13:0] _GEN_8729 = 14'h2219 == index ? 14'h112 : _GEN_8728;
  wire [13:0] _GEN_8730 = 14'h221a == index ? 14'h110 : _GEN_8729;
  wire [13:0] _GEN_8731 = 14'h221b == index ? 14'h10e : _GEN_8730;
  wire [13:0] _GEN_8732 = 14'h221c == index ? 14'h10c : _GEN_8731;
  wire [13:0] _GEN_8733 = 14'h221d == index ? 14'h10a : _GEN_8732;
  wire [13:0] _GEN_8734 = 14'h221e == index ? 14'h108 : _GEN_8733;
  wire [13:0] _GEN_8735 = 14'h221f == index ? 14'h106 : _GEN_8734;
  wire [13:0] _GEN_8736 = 14'h2220 == index ? 14'h104 : _GEN_8735;
  wire [13:0] _GEN_8737 = 14'h2221 == index ? 14'h102 : _GEN_8736;
  wire [13:0] _GEN_8738 = 14'h2222 == index ? 14'h100 : _GEN_8737;
  wire [13:0] _GEN_8739 = 14'h2223 == index ? 14'ha1 : _GEN_8738;
  wire [13:0] _GEN_8740 = 14'h2224 == index ? 14'ha0 : _GEN_8739;
  wire [13:0] _GEN_8741 = 14'h2225 == index ? 14'h9f : _GEN_8740;
  wire [13:0] _GEN_8742 = 14'h2226 == index ? 14'h9e : _GEN_8741;
  wire [13:0] _GEN_8743 = 14'h2227 == index ? 14'h9d : _GEN_8742;
  wire [13:0] _GEN_8744 = 14'h2228 == index ? 14'h9c : _GEN_8743;
  wire [13:0] _GEN_8745 = 14'h2229 == index ? 14'h9b : _GEN_8744;
  wire [13:0] _GEN_8746 = 14'h222a == index ? 14'h9a : _GEN_8745;
  wire [13:0] _GEN_8747 = 14'h222b == index ? 14'h99 : _GEN_8746;
  wire [13:0] _GEN_8748 = 14'h222c == index ? 14'h98 : _GEN_8747;
  wire [13:0] _GEN_8749 = 14'h222d == index ? 14'h97 : _GEN_8748;
  wire [13:0] _GEN_8750 = 14'h222e == index ? 14'h96 : _GEN_8749;
  wire [13:0] _GEN_8751 = 14'h222f == index ? 14'h95 : _GEN_8750;
  wire [13:0] _GEN_8752 = 14'h2230 == index ? 14'h94 : _GEN_8751;
  wire [13:0] _GEN_8753 = 14'h2231 == index ? 14'h93 : _GEN_8752;
  wire [13:0] _GEN_8754 = 14'h2232 == index ? 14'h92 : _GEN_8753;
  wire [13:0] _GEN_8755 = 14'h2233 == index ? 14'h91 : _GEN_8754;
  wire [13:0] _GEN_8756 = 14'h2234 == index ? 14'h90 : _GEN_8755;
  wire [13:0] _GEN_8757 = 14'h2235 == index ? 14'h8f : _GEN_8756;
  wire [13:0] _GEN_8758 = 14'h2236 == index ? 14'h8e : _GEN_8757;
  wire [13:0] _GEN_8759 = 14'h2237 == index ? 14'h8d : _GEN_8758;
  wire [13:0] _GEN_8760 = 14'h2238 == index ? 14'h8c : _GEN_8759;
  wire [13:0] _GEN_8761 = 14'h2239 == index ? 14'h8b : _GEN_8760;
  wire [13:0] _GEN_8762 = 14'h223a == index ? 14'h8a : _GEN_8761;
  wire [13:0] _GEN_8763 = 14'h223b == index ? 14'h89 : _GEN_8762;
  wire [13:0] _GEN_8764 = 14'h223c == index ? 14'h88 : _GEN_8763;
  wire [13:0] _GEN_8765 = 14'h223d == index ? 14'h87 : _GEN_8764;
  wire [13:0] _GEN_8766 = 14'h223e == index ? 14'h86 : _GEN_8765;
  wire [13:0] _GEN_8767 = 14'h223f == index ? 14'h85 : _GEN_8766;
  wire [13:0] _GEN_8768 = 14'h2240 == index ? 14'h84 : _GEN_8767;
  wire [13:0] _GEN_8769 = 14'h2241 == index ? 14'h83 : _GEN_8768;
  wire [13:0] _GEN_8770 = 14'h2242 == index ? 14'h82 : _GEN_8769;
  wire [13:0] _GEN_8771 = 14'h2243 == index ? 14'h81 : _GEN_8770;
  wire [13:0] _GEN_8772 = 14'h2244 == index ? 14'h80 : _GEN_8771;
  wire [13:0] _GEN_8773 = 14'h2245 == index ? 14'h44 : _GEN_8772;
  wire [13:0] _GEN_8774 = 14'h2246 == index ? 14'h44 : _GEN_8773;
  wire [13:0] _GEN_8775 = 14'h2247 == index ? 14'h44 : _GEN_8774;
  wire [13:0] _GEN_8776 = 14'h2248 == index ? 14'h44 : _GEN_8775;
  wire [13:0] _GEN_8777 = 14'h2249 == index ? 14'h44 : _GEN_8776;
  wire [13:0] _GEN_8778 = 14'h224a == index ? 14'h44 : _GEN_8777;
  wire [13:0] _GEN_8779 = 14'h224b == index ? 14'h44 : _GEN_8778;
  wire [13:0] _GEN_8780 = 14'h224c == index ? 14'h44 : _GEN_8779;
  wire [13:0] _GEN_8781 = 14'h224d == index ? 14'h44 : _GEN_8780;
  wire [13:0] _GEN_8782 = 14'h224e == index ? 14'h44 : _GEN_8781;
  wire [13:0] _GEN_8783 = 14'h224f == index ? 14'h44 : _GEN_8782;
  wire [13:0] _GEN_8784 = 14'h2250 == index ? 14'h44 : _GEN_8783;
  wire [13:0] _GEN_8785 = 14'h2251 == index ? 14'h44 : _GEN_8784;
  wire [13:0] _GEN_8786 = 14'h2252 == index ? 14'h44 : _GEN_8785;
  wire [13:0] _GEN_8787 = 14'h2253 == index ? 14'h44 : _GEN_8786;
  wire [13:0] _GEN_8788 = 14'h2254 == index ? 14'h44 : _GEN_8787;
  wire [13:0] _GEN_8789 = 14'h2255 == index ? 14'h44 : _GEN_8788;
  wire [13:0] _GEN_8790 = 14'h2256 == index ? 14'h44 : _GEN_8789;
  wire [13:0] _GEN_8791 = 14'h2257 == index ? 14'h44 : _GEN_8790;
  wire [13:0] _GEN_8792 = 14'h2258 == index ? 14'h44 : _GEN_8791;
  wire [13:0] _GEN_8793 = 14'h2259 == index ? 14'h44 : _GEN_8792;
  wire [13:0] _GEN_8794 = 14'h225a == index ? 14'h44 : _GEN_8793;
  wire [13:0] _GEN_8795 = 14'h225b == index ? 14'h44 : _GEN_8794;
  wire [13:0] _GEN_8796 = 14'h225c == index ? 14'h44 : _GEN_8795;
  wire [13:0] _GEN_8797 = 14'h225d == index ? 14'h44 : _GEN_8796;
  wire [13:0] _GEN_8798 = 14'h225e == index ? 14'h44 : _GEN_8797;
  wire [13:0] _GEN_8799 = 14'h225f == index ? 14'h44 : _GEN_8798;
  wire [13:0] _GEN_8800 = 14'h2260 == index ? 14'h44 : _GEN_8799;
  wire [13:0] _GEN_8801 = 14'h2261 == index ? 14'h44 : _GEN_8800;
  wire [13:0] _GEN_8802 = 14'h2262 == index ? 14'h44 : _GEN_8801;
  wire [13:0] _GEN_8803 = 14'h2263 == index ? 14'h44 : _GEN_8802;
  wire [13:0] _GEN_8804 = 14'h2264 == index ? 14'h44 : _GEN_8803;
  wire [13:0] _GEN_8805 = 14'h2265 == index ? 14'h44 : _GEN_8804;
  wire [13:0] _GEN_8806 = 14'h2266 == index ? 14'h44 : _GEN_8805;
  wire [13:0] _GEN_8807 = 14'h2267 == index ? 14'h44 : _GEN_8806;
  wire [13:0] _GEN_8808 = 14'h2268 == index ? 14'h44 : _GEN_8807;
  wire [13:0] _GEN_8809 = 14'h2269 == index ? 14'h44 : _GEN_8808;
  wire [13:0] _GEN_8810 = 14'h226a == index ? 14'h44 : _GEN_8809;
  wire [13:0] _GEN_8811 = 14'h226b == index ? 14'h44 : _GEN_8810;
  wire [13:0] _GEN_8812 = 14'h226c == index ? 14'h44 : _GEN_8811;
  wire [13:0] _GEN_8813 = 14'h226d == index ? 14'h44 : _GEN_8812;
  wire [13:0] _GEN_8814 = 14'h226e == index ? 14'h44 : _GEN_8813;
  wire [13:0] _GEN_8815 = 14'h226f == index ? 14'h44 : _GEN_8814;
  wire [13:0] _GEN_8816 = 14'h2270 == index ? 14'h44 : _GEN_8815;
  wire [13:0] _GEN_8817 = 14'h2271 == index ? 14'h44 : _GEN_8816;
  wire [13:0] _GEN_8818 = 14'h2272 == index ? 14'h44 : _GEN_8817;
  wire [13:0] _GEN_8819 = 14'h2273 == index ? 14'h44 : _GEN_8818;
  wire [13:0] _GEN_8820 = 14'h2274 == index ? 14'h44 : _GEN_8819;
  wire [13:0] _GEN_8821 = 14'h2275 == index ? 14'h44 : _GEN_8820;
  wire [13:0] _GEN_8822 = 14'h2276 == index ? 14'h44 : _GEN_8821;
  wire [13:0] _GEN_8823 = 14'h2277 == index ? 14'h44 : _GEN_8822;
  wire [13:0] _GEN_8824 = 14'h2278 == index ? 14'h44 : _GEN_8823;
  wire [13:0] _GEN_8825 = 14'h2279 == index ? 14'h44 : _GEN_8824;
  wire [13:0] _GEN_8826 = 14'h227a == index ? 14'h44 : _GEN_8825;
  wire [13:0] _GEN_8827 = 14'h227b == index ? 14'h44 : _GEN_8826;
  wire [13:0] _GEN_8828 = 14'h227c == index ? 14'h44 : _GEN_8827;
  wire [13:0] _GEN_8829 = 14'h227d == index ? 14'h44 : _GEN_8828;
  wire [13:0] _GEN_8830 = 14'h227e == index ? 14'h44 : _GEN_8829;
  wire [13:0] _GEN_8831 = 14'h227f == index ? 14'h44 : _GEN_8830;
  wire [13:0] _GEN_8832 = 14'h2280 == index ? 14'h0 : _GEN_8831;
  wire [13:0] _GEN_8833 = 14'h2281 == index ? 14'h2280 : _GEN_8832;
  wire [13:0] _GEN_8834 = 14'h2282 == index ? 14'h1101 : _GEN_8833;
  wire [13:0] _GEN_8835 = 14'h2283 == index ? 14'hb80 : _GEN_8834;
  wire [13:0] _GEN_8836 = 14'h2284 == index ? 14'h881 : _GEN_8835;
  wire [13:0] _GEN_8837 = 14'h2285 == index ? 14'h684 : _GEN_8836;
  wire [13:0] _GEN_8838 = 14'h2286 == index ? 14'h583 : _GEN_8837;
  wire [13:0] _GEN_8839 = 14'h2287 == index ? 14'h486 : _GEN_8838;
  wire [13:0] _GEN_8840 = 14'h2288 == index ? 14'h405 : _GEN_8839;
  wire [13:0] _GEN_8841 = 14'h2289 == index ? 14'h386 : _GEN_8840;
  wire [13:0] _GEN_8842 = 14'h228a == index ? 14'h309 : _GEN_8841;
  wire [13:0] _GEN_8843 = 14'h228b == index ? 14'h303 : _GEN_8842;
  wire [13:0] _GEN_8844 = 14'h228c == index ? 14'h289 : _GEN_8843;
  wire [13:0] _GEN_8845 = 14'h228d == index ? 14'h284 : _GEN_8844;
  wire [13:0] _GEN_8846 = 14'h228e == index ? 14'h20d : _GEN_8845;
  wire [13:0] _GEN_8847 = 14'h228f == index ? 14'h209 : _GEN_8846;
  wire [13:0] _GEN_8848 = 14'h2290 == index ? 14'h205 : _GEN_8847;
  wire [13:0] _GEN_8849 = 14'h2291 == index ? 14'h201 : _GEN_8848;
  wire [13:0] _GEN_8850 = 14'h2292 == index ? 14'h18f : _GEN_8849;
  wire [13:0] _GEN_8851 = 14'h2293 == index ? 14'h18c : _GEN_8850;
  wire [13:0] _GEN_8852 = 14'h2294 == index ? 14'h189 : _GEN_8851;
  wire [13:0] _GEN_8853 = 14'h2295 == index ? 14'h186 : _GEN_8852;
  wire [13:0] _GEN_8854 = 14'h2296 == index ? 14'h183 : _GEN_8853;
  wire [13:0] _GEN_8855 = 14'h2297 == index ? 14'h180 : _GEN_8854;
  wire [13:0] _GEN_8856 = 14'h2298 == index ? 14'h115 : _GEN_8855;
  wire [13:0] _GEN_8857 = 14'h2299 == index ? 14'h113 : _GEN_8856;
  wire [13:0] _GEN_8858 = 14'h229a == index ? 14'h111 : _GEN_8857;
  wire [13:0] _GEN_8859 = 14'h229b == index ? 14'h10f : _GEN_8858;
  wire [13:0] _GEN_8860 = 14'h229c == index ? 14'h10d : _GEN_8859;
  wire [13:0] _GEN_8861 = 14'h229d == index ? 14'h10b : _GEN_8860;
  wire [13:0] _GEN_8862 = 14'h229e == index ? 14'h109 : _GEN_8861;
  wire [13:0] _GEN_8863 = 14'h229f == index ? 14'h107 : _GEN_8862;
  wire [13:0] _GEN_8864 = 14'h22a0 == index ? 14'h105 : _GEN_8863;
  wire [13:0] _GEN_8865 = 14'h22a1 == index ? 14'h103 : _GEN_8864;
  wire [13:0] _GEN_8866 = 14'h22a2 == index ? 14'h101 : _GEN_8865;
  wire [13:0] _GEN_8867 = 14'h22a3 == index ? 14'ha2 : _GEN_8866;
  wire [13:0] _GEN_8868 = 14'h22a4 == index ? 14'ha1 : _GEN_8867;
  wire [13:0] _GEN_8869 = 14'h22a5 == index ? 14'ha0 : _GEN_8868;
  wire [13:0] _GEN_8870 = 14'h22a6 == index ? 14'h9f : _GEN_8869;
  wire [13:0] _GEN_8871 = 14'h22a7 == index ? 14'h9e : _GEN_8870;
  wire [13:0] _GEN_8872 = 14'h22a8 == index ? 14'h9d : _GEN_8871;
  wire [13:0] _GEN_8873 = 14'h22a9 == index ? 14'h9c : _GEN_8872;
  wire [13:0] _GEN_8874 = 14'h22aa == index ? 14'h9b : _GEN_8873;
  wire [13:0] _GEN_8875 = 14'h22ab == index ? 14'h9a : _GEN_8874;
  wire [13:0] _GEN_8876 = 14'h22ac == index ? 14'h99 : _GEN_8875;
  wire [13:0] _GEN_8877 = 14'h22ad == index ? 14'h98 : _GEN_8876;
  wire [13:0] _GEN_8878 = 14'h22ae == index ? 14'h97 : _GEN_8877;
  wire [13:0] _GEN_8879 = 14'h22af == index ? 14'h96 : _GEN_8878;
  wire [13:0] _GEN_8880 = 14'h22b0 == index ? 14'h95 : _GEN_8879;
  wire [13:0] _GEN_8881 = 14'h22b1 == index ? 14'h94 : _GEN_8880;
  wire [13:0] _GEN_8882 = 14'h22b2 == index ? 14'h93 : _GEN_8881;
  wire [13:0] _GEN_8883 = 14'h22b3 == index ? 14'h92 : _GEN_8882;
  wire [13:0] _GEN_8884 = 14'h22b4 == index ? 14'h91 : _GEN_8883;
  wire [13:0] _GEN_8885 = 14'h22b5 == index ? 14'h90 : _GEN_8884;
  wire [13:0] _GEN_8886 = 14'h22b6 == index ? 14'h8f : _GEN_8885;
  wire [13:0] _GEN_8887 = 14'h22b7 == index ? 14'h8e : _GEN_8886;
  wire [13:0] _GEN_8888 = 14'h22b8 == index ? 14'h8d : _GEN_8887;
  wire [13:0] _GEN_8889 = 14'h22b9 == index ? 14'h8c : _GEN_8888;
  wire [13:0] _GEN_8890 = 14'h22ba == index ? 14'h8b : _GEN_8889;
  wire [13:0] _GEN_8891 = 14'h22bb == index ? 14'h8a : _GEN_8890;
  wire [13:0] _GEN_8892 = 14'h22bc == index ? 14'h89 : _GEN_8891;
  wire [13:0] _GEN_8893 = 14'h22bd == index ? 14'h88 : _GEN_8892;
  wire [13:0] _GEN_8894 = 14'h22be == index ? 14'h87 : _GEN_8893;
  wire [13:0] _GEN_8895 = 14'h22bf == index ? 14'h86 : _GEN_8894;
  wire [13:0] _GEN_8896 = 14'h22c0 == index ? 14'h85 : _GEN_8895;
  wire [13:0] _GEN_8897 = 14'h22c1 == index ? 14'h84 : _GEN_8896;
  wire [13:0] _GEN_8898 = 14'h22c2 == index ? 14'h83 : _GEN_8897;
  wire [13:0] _GEN_8899 = 14'h22c3 == index ? 14'h82 : _GEN_8898;
  wire [13:0] _GEN_8900 = 14'h22c4 == index ? 14'h81 : _GEN_8899;
  wire [13:0] _GEN_8901 = 14'h22c5 == index ? 14'h80 : _GEN_8900;
  wire [13:0] _GEN_8902 = 14'h22c6 == index ? 14'h45 : _GEN_8901;
  wire [13:0] _GEN_8903 = 14'h22c7 == index ? 14'h45 : _GEN_8902;
  wire [13:0] _GEN_8904 = 14'h22c8 == index ? 14'h45 : _GEN_8903;
  wire [13:0] _GEN_8905 = 14'h22c9 == index ? 14'h45 : _GEN_8904;
  wire [13:0] _GEN_8906 = 14'h22ca == index ? 14'h45 : _GEN_8905;
  wire [13:0] _GEN_8907 = 14'h22cb == index ? 14'h45 : _GEN_8906;
  wire [13:0] _GEN_8908 = 14'h22cc == index ? 14'h45 : _GEN_8907;
  wire [13:0] _GEN_8909 = 14'h22cd == index ? 14'h45 : _GEN_8908;
  wire [13:0] _GEN_8910 = 14'h22ce == index ? 14'h45 : _GEN_8909;
  wire [13:0] _GEN_8911 = 14'h22cf == index ? 14'h45 : _GEN_8910;
  wire [13:0] _GEN_8912 = 14'h22d0 == index ? 14'h45 : _GEN_8911;
  wire [13:0] _GEN_8913 = 14'h22d1 == index ? 14'h45 : _GEN_8912;
  wire [13:0] _GEN_8914 = 14'h22d2 == index ? 14'h45 : _GEN_8913;
  wire [13:0] _GEN_8915 = 14'h22d3 == index ? 14'h45 : _GEN_8914;
  wire [13:0] _GEN_8916 = 14'h22d4 == index ? 14'h45 : _GEN_8915;
  wire [13:0] _GEN_8917 = 14'h22d5 == index ? 14'h45 : _GEN_8916;
  wire [13:0] _GEN_8918 = 14'h22d6 == index ? 14'h45 : _GEN_8917;
  wire [13:0] _GEN_8919 = 14'h22d7 == index ? 14'h45 : _GEN_8918;
  wire [13:0] _GEN_8920 = 14'h22d8 == index ? 14'h45 : _GEN_8919;
  wire [13:0] _GEN_8921 = 14'h22d9 == index ? 14'h45 : _GEN_8920;
  wire [13:0] _GEN_8922 = 14'h22da == index ? 14'h45 : _GEN_8921;
  wire [13:0] _GEN_8923 = 14'h22db == index ? 14'h45 : _GEN_8922;
  wire [13:0] _GEN_8924 = 14'h22dc == index ? 14'h45 : _GEN_8923;
  wire [13:0] _GEN_8925 = 14'h22dd == index ? 14'h45 : _GEN_8924;
  wire [13:0] _GEN_8926 = 14'h22de == index ? 14'h45 : _GEN_8925;
  wire [13:0] _GEN_8927 = 14'h22df == index ? 14'h45 : _GEN_8926;
  wire [13:0] _GEN_8928 = 14'h22e0 == index ? 14'h45 : _GEN_8927;
  wire [13:0] _GEN_8929 = 14'h22e1 == index ? 14'h45 : _GEN_8928;
  wire [13:0] _GEN_8930 = 14'h22e2 == index ? 14'h45 : _GEN_8929;
  wire [13:0] _GEN_8931 = 14'h22e3 == index ? 14'h45 : _GEN_8930;
  wire [13:0] _GEN_8932 = 14'h22e4 == index ? 14'h45 : _GEN_8931;
  wire [13:0] _GEN_8933 = 14'h22e5 == index ? 14'h45 : _GEN_8932;
  wire [13:0] _GEN_8934 = 14'h22e6 == index ? 14'h45 : _GEN_8933;
  wire [13:0] _GEN_8935 = 14'h22e7 == index ? 14'h45 : _GEN_8934;
  wire [13:0] _GEN_8936 = 14'h22e8 == index ? 14'h45 : _GEN_8935;
  wire [13:0] _GEN_8937 = 14'h22e9 == index ? 14'h45 : _GEN_8936;
  wire [13:0] _GEN_8938 = 14'h22ea == index ? 14'h45 : _GEN_8937;
  wire [13:0] _GEN_8939 = 14'h22eb == index ? 14'h45 : _GEN_8938;
  wire [13:0] _GEN_8940 = 14'h22ec == index ? 14'h45 : _GEN_8939;
  wire [13:0] _GEN_8941 = 14'h22ed == index ? 14'h45 : _GEN_8940;
  wire [13:0] _GEN_8942 = 14'h22ee == index ? 14'h45 : _GEN_8941;
  wire [13:0] _GEN_8943 = 14'h22ef == index ? 14'h45 : _GEN_8942;
  wire [13:0] _GEN_8944 = 14'h22f0 == index ? 14'h45 : _GEN_8943;
  wire [13:0] _GEN_8945 = 14'h22f1 == index ? 14'h45 : _GEN_8944;
  wire [13:0] _GEN_8946 = 14'h22f2 == index ? 14'h45 : _GEN_8945;
  wire [13:0] _GEN_8947 = 14'h22f3 == index ? 14'h45 : _GEN_8946;
  wire [13:0] _GEN_8948 = 14'h22f4 == index ? 14'h45 : _GEN_8947;
  wire [13:0] _GEN_8949 = 14'h22f5 == index ? 14'h45 : _GEN_8948;
  wire [13:0] _GEN_8950 = 14'h22f6 == index ? 14'h45 : _GEN_8949;
  wire [13:0] _GEN_8951 = 14'h22f7 == index ? 14'h45 : _GEN_8950;
  wire [13:0] _GEN_8952 = 14'h22f8 == index ? 14'h45 : _GEN_8951;
  wire [13:0] _GEN_8953 = 14'h22f9 == index ? 14'h45 : _GEN_8952;
  wire [13:0] _GEN_8954 = 14'h22fa == index ? 14'h45 : _GEN_8953;
  wire [13:0] _GEN_8955 = 14'h22fb == index ? 14'h45 : _GEN_8954;
  wire [13:0] _GEN_8956 = 14'h22fc == index ? 14'h45 : _GEN_8955;
  wire [13:0] _GEN_8957 = 14'h22fd == index ? 14'h45 : _GEN_8956;
  wire [13:0] _GEN_8958 = 14'h22fe == index ? 14'h45 : _GEN_8957;
  wire [13:0] _GEN_8959 = 14'h22ff == index ? 14'h45 : _GEN_8958;
  wire [13:0] _GEN_8960 = 14'h2300 == index ? 14'h0 : _GEN_8959;
  wire [13:0] _GEN_8961 = 14'h2301 == index ? 14'h2300 : _GEN_8960;
  wire [13:0] _GEN_8962 = 14'h2302 == index ? 14'h1180 : _GEN_8961;
  wire [13:0] _GEN_8963 = 14'h2303 == index ? 14'hb81 : _GEN_8962;
  wire [13:0] _GEN_8964 = 14'h2304 == index ? 14'h882 : _GEN_8963;
  wire [13:0] _GEN_8965 = 14'h2305 == index ? 14'h700 : _GEN_8964;
  wire [13:0] _GEN_8966 = 14'h2306 == index ? 14'h584 : _GEN_8965;
  wire [13:0] _GEN_8967 = 14'h2307 == index ? 14'h500 : _GEN_8966;
  wire [13:0] _GEN_8968 = 14'h2308 == index ? 14'h406 : _GEN_8967;
  wire [13:0] _GEN_8969 = 14'h2309 == index ? 14'h387 : _GEN_8968;
  wire [13:0] _GEN_8970 = 14'h230a == index ? 14'h380 : _GEN_8969;
  wire [13:0] _GEN_8971 = 14'h230b == index ? 14'h304 : _GEN_8970;
  wire [13:0] _GEN_8972 = 14'h230c == index ? 14'h28a : _GEN_8971;
  wire [13:0] _GEN_8973 = 14'h230d == index ? 14'h285 : _GEN_8972;
  wire [13:0] _GEN_8974 = 14'h230e == index ? 14'h280 : _GEN_8973;
  wire [13:0] _GEN_8975 = 14'h230f == index ? 14'h20a : _GEN_8974;
  wire [13:0] _GEN_8976 = 14'h2310 == index ? 14'h206 : _GEN_8975;
  wire [13:0] _GEN_8977 = 14'h2311 == index ? 14'h202 : _GEN_8976;
  wire [13:0] _GEN_8978 = 14'h2312 == index ? 14'h190 : _GEN_8977;
  wire [13:0] _GEN_8979 = 14'h2313 == index ? 14'h18d : _GEN_8978;
  wire [13:0] _GEN_8980 = 14'h2314 == index ? 14'h18a : _GEN_8979;
  wire [13:0] _GEN_8981 = 14'h2315 == index ? 14'h187 : _GEN_8980;
  wire [13:0] _GEN_8982 = 14'h2316 == index ? 14'h184 : _GEN_8981;
  wire [13:0] _GEN_8983 = 14'h2317 == index ? 14'h181 : _GEN_8982;
  wire [13:0] _GEN_8984 = 14'h2318 == index ? 14'h116 : _GEN_8983;
  wire [13:0] _GEN_8985 = 14'h2319 == index ? 14'h114 : _GEN_8984;
  wire [13:0] _GEN_8986 = 14'h231a == index ? 14'h112 : _GEN_8985;
  wire [13:0] _GEN_8987 = 14'h231b == index ? 14'h110 : _GEN_8986;
  wire [13:0] _GEN_8988 = 14'h231c == index ? 14'h10e : _GEN_8987;
  wire [13:0] _GEN_8989 = 14'h231d == index ? 14'h10c : _GEN_8988;
  wire [13:0] _GEN_8990 = 14'h231e == index ? 14'h10a : _GEN_8989;
  wire [13:0] _GEN_8991 = 14'h231f == index ? 14'h108 : _GEN_8990;
  wire [13:0] _GEN_8992 = 14'h2320 == index ? 14'h106 : _GEN_8991;
  wire [13:0] _GEN_8993 = 14'h2321 == index ? 14'h104 : _GEN_8992;
  wire [13:0] _GEN_8994 = 14'h2322 == index ? 14'h102 : _GEN_8993;
  wire [13:0] _GEN_8995 = 14'h2323 == index ? 14'h100 : _GEN_8994;
  wire [13:0] _GEN_8996 = 14'h2324 == index ? 14'ha2 : _GEN_8995;
  wire [13:0] _GEN_8997 = 14'h2325 == index ? 14'ha1 : _GEN_8996;
  wire [13:0] _GEN_8998 = 14'h2326 == index ? 14'ha0 : _GEN_8997;
  wire [13:0] _GEN_8999 = 14'h2327 == index ? 14'h9f : _GEN_8998;
  wire [13:0] _GEN_9000 = 14'h2328 == index ? 14'h9e : _GEN_8999;
  wire [13:0] _GEN_9001 = 14'h2329 == index ? 14'h9d : _GEN_9000;
  wire [13:0] _GEN_9002 = 14'h232a == index ? 14'h9c : _GEN_9001;
  wire [13:0] _GEN_9003 = 14'h232b == index ? 14'h9b : _GEN_9002;
  wire [13:0] _GEN_9004 = 14'h232c == index ? 14'h9a : _GEN_9003;
  wire [13:0] _GEN_9005 = 14'h232d == index ? 14'h99 : _GEN_9004;
  wire [13:0] _GEN_9006 = 14'h232e == index ? 14'h98 : _GEN_9005;
  wire [13:0] _GEN_9007 = 14'h232f == index ? 14'h97 : _GEN_9006;
  wire [13:0] _GEN_9008 = 14'h2330 == index ? 14'h96 : _GEN_9007;
  wire [13:0] _GEN_9009 = 14'h2331 == index ? 14'h95 : _GEN_9008;
  wire [13:0] _GEN_9010 = 14'h2332 == index ? 14'h94 : _GEN_9009;
  wire [13:0] _GEN_9011 = 14'h2333 == index ? 14'h93 : _GEN_9010;
  wire [13:0] _GEN_9012 = 14'h2334 == index ? 14'h92 : _GEN_9011;
  wire [13:0] _GEN_9013 = 14'h2335 == index ? 14'h91 : _GEN_9012;
  wire [13:0] _GEN_9014 = 14'h2336 == index ? 14'h90 : _GEN_9013;
  wire [13:0] _GEN_9015 = 14'h2337 == index ? 14'h8f : _GEN_9014;
  wire [13:0] _GEN_9016 = 14'h2338 == index ? 14'h8e : _GEN_9015;
  wire [13:0] _GEN_9017 = 14'h2339 == index ? 14'h8d : _GEN_9016;
  wire [13:0] _GEN_9018 = 14'h233a == index ? 14'h8c : _GEN_9017;
  wire [13:0] _GEN_9019 = 14'h233b == index ? 14'h8b : _GEN_9018;
  wire [13:0] _GEN_9020 = 14'h233c == index ? 14'h8a : _GEN_9019;
  wire [13:0] _GEN_9021 = 14'h233d == index ? 14'h89 : _GEN_9020;
  wire [13:0] _GEN_9022 = 14'h233e == index ? 14'h88 : _GEN_9021;
  wire [13:0] _GEN_9023 = 14'h233f == index ? 14'h87 : _GEN_9022;
  wire [13:0] _GEN_9024 = 14'h2340 == index ? 14'h86 : _GEN_9023;
  wire [13:0] _GEN_9025 = 14'h2341 == index ? 14'h85 : _GEN_9024;
  wire [13:0] _GEN_9026 = 14'h2342 == index ? 14'h84 : _GEN_9025;
  wire [13:0] _GEN_9027 = 14'h2343 == index ? 14'h83 : _GEN_9026;
  wire [13:0] _GEN_9028 = 14'h2344 == index ? 14'h82 : _GEN_9027;
  wire [13:0] _GEN_9029 = 14'h2345 == index ? 14'h81 : _GEN_9028;
  wire [13:0] _GEN_9030 = 14'h2346 == index ? 14'h80 : _GEN_9029;
  wire [13:0] _GEN_9031 = 14'h2347 == index ? 14'h46 : _GEN_9030;
  wire [13:0] _GEN_9032 = 14'h2348 == index ? 14'h46 : _GEN_9031;
  wire [13:0] _GEN_9033 = 14'h2349 == index ? 14'h46 : _GEN_9032;
  wire [13:0] _GEN_9034 = 14'h234a == index ? 14'h46 : _GEN_9033;
  wire [13:0] _GEN_9035 = 14'h234b == index ? 14'h46 : _GEN_9034;
  wire [13:0] _GEN_9036 = 14'h234c == index ? 14'h46 : _GEN_9035;
  wire [13:0] _GEN_9037 = 14'h234d == index ? 14'h46 : _GEN_9036;
  wire [13:0] _GEN_9038 = 14'h234e == index ? 14'h46 : _GEN_9037;
  wire [13:0] _GEN_9039 = 14'h234f == index ? 14'h46 : _GEN_9038;
  wire [13:0] _GEN_9040 = 14'h2350 == index ? 14'h46 : _GEN_9039;
  wire [13:0] _GEN_9041 = 14'h2351 == index ? 14'h46 : _GEN_9040;
  wire [13:0] _GEN_9042 = 14'h2352 == index ? 14'h46 : _GEN_9041;
  wire [13:0] _GEN_9043 = 14'h2353 == index ? 14'h46 : _GEN_9042;
  wire [13:0] _GEN_9044 = 14'h2354 == index ? 14'h46 : _GEN_9043;
  wire [13:0] _GEN_9045 = 14'h2355 == index ? 14'h46 : _GEN_9044;
  wire [13:0] _GEN_9046 = 14'h2356 == index ? 14'h46 : _GEN_9045;
  wire [13:0] _GEN_9047 = 14'h2357 == index ? 14'h46 : _GEN_9046;
  wire [13:0] _GEN_9048 = 14'h2358 == index ? 14'h46 : _GEN_9047;
  wire [13:0] _GEN_9049 = 14'h2359 == index ? 14'h46 : _GEN_9048;
  wire [13:0] _GEN_9050 = 14'h235a == index ? 14'h46 : _GEN_9049;
  wire [13:0] _GEN_9051 = 14'h235b == index ? 14'h46 : _GEN_9050;
  wire [13:0] _GEN_9052 = 14'h235c == index ? 14'h46 : _GEN_9051;
  wire [13:0] _GEN_9053 = 14'h235d == index ? 14'h46 : _GEN_9052;
  wire [13:0] _GEN_9054 = 14'h235e == index ? 14'h46 : _GEN_9053;
  wire [13:0] _GEN_9055 = 14'h235f == index ? 14'h46 : _GEN_9054;
  wire [13:0] _GEN_9056 = 14'h2360 == index ? 14'h46 : _GEN_9055;
  wire [13:0] _GEN_9057 = 14'h2361 == index ? 14'h46 : _GEN_9056;
  wire [13:0] _GEN_9058 = 14'h2362 == index ? 14'h46 : _GEN_9057;
  wire [13:0] _GEN_9059 = 14'h2363 == index ? 14'h46 : _GEN_9058;
  wire [13:0] _GEN_9060 = 14'h2364 == index ? 14'h46 : _GEN_9059;
  wire [13:0] _GEN_9061 = 14'h2365 == index ? 14'h46 : _GEN_9060;
  wire [13:0] _GEN_9062 = 14'h2366 == index ? 14'h46 : _GEN_9061;
  wire [13:0] _GEN_9063 = 14'h2367 == index ? 14'h46 : _GEN_9062;
  wire [13:0] _GEN_9064 = 14'h2368 == index ? 14'h46 : _GEN_9063;
  wire [13:0] _GEN_9065 = 14'h2369 == index ? 14'h46 : _GEN_9064;
  wire [13:0] _GEN_9066 = 14'h236a == index ? 14'h46 : _GEN_9065;
  wire [13:0] _GEN_9067 = 14'h236b == index ? 14'h46 : _GEN_9066;
  wire [13:0] _GEN_9068 = 14'h236c == index ? 14'h46 : _GEN_9067;
  wire [13:0] _GEN_9069 = 14'h236d == index ? 14'h46 : _GEN_9068;
  wire [13:0] _GEN_9070 = 14'h236e == index ? 14'h46 : _GEN_9069;
  wire [13:0] _GEN_9071 = 14'h236f == index ? 14'h46 : _GEN_9070;
  wire [13:0] _GEN_9072 = 14'h2370 == index ? 14'h46 : _GEN_9071;
  wire [13:0] _GEN_9073 = 14'h2371 == index ? 14'h46 : _GEN_9072;
  wire [13:0] _GEN_9074 = 14'h2372 == index ? 14'h46 : _GEN_9073;
  wire [13:0] _GEN_9075 = 14'h2373 == index ? 14'h46 : _GEN_9074;
  wire [13:0] _GEN_9076 = 14'h2374 == index ? 14'h46 : _GEN_9075;
  wire [13:0] _GEN_9077 = 14'h2375 == index ? 14'h46 : _GEN_9076;
  wire [13:0] _GEN_9078 = 14'h2376 == index ? 14'h46 : _GEN_9077;
  wire [13:0] _GEN_9079 = 14'h2377 == index ? 14'h46 : _GEN_9078;
  wire [13:0] _GEN_9080 = 14'h2378 == index ? 14'h46 : _GEN_9079;
  wire [13:0] _GEN_9081 = 14'h2379 == index ? 14'h46 : _GEN_9080;
  wire [13:0] _GEN_9082 = 14'h237a == index ? 14'h46 : _GEN_9081;
  wire [13:0] _GEN_9083 = 14'h237b == index ? 14'h46 : _GEN_9082;
  wire [13:0] _GEN_9084 = 14'h237c == index ? 14'h46 : _GEN_9083;
  wire [13:0] _GEN_9085 = 14'h237d == index ? 14'h46 : _GEN_9084;
  wire [13:0] _GEN_9086 = 14'h237e == index ? 14'h46 : _GEN_9085;
  wire [13:0] _GEN_9087 = 14'h237f == index ? 14'h46 : _GEN_9086;
  wire [13:0] _GEN_9088 = 14'h2380 == index ? 14'h0 : _GEN_9087;
  wire [13:0] _GEN_9089 = 14'h2381 == index ? 14'h2380 : _GEN_9088;
  wire [13:0] _GEN_9090 = 14'h2382 == index ? 14'h1181 : _GEN_9089;
  wire [13:0] _GEN_9091 = 14'h2383 == index ? 14'hb82 : _GEN_9090;
  wire [13:0] _GEN_9092 = 14'h2384 == index ? 14'h883 : _GEN_9091;
  wire [13:0] _GEN_9093 = 14'h2385 == index ? 14'h701 : _GEN_9092;
  wire [13:0] _GEN_9094 = 14'h2386 == index ? 14'h585 : _GEN_9093;
  wire [13:0] _GEN_9095 = 14'h2387 == index ? 14'h501 : _GEN_9094;
  wire [13:0] _GEN_9096 = 14'h2388 == index ? 14'h407 : _GEN_9095;
  wire [13:0] _GEN_9097 = 14'h2389 == index ? 14'h388 : _GEN_9096;
  wire [13:0] _GEN_9098 = 14'h238a == index ? 14'h381 : _GEN_9097;
  wire [13:0] _GEN_9099 = 14'h238b == index ? 14'h305 : _GEN_9098;
  wire [13:0] _GEN_9100 = 14'h238c == index ? 14'h28b : _GEN_9099;
  wire [13:0] _GEN_9101 = 14'h238d == index ? 14'h286 : _GEN_9100;
  wire [13:0] _GEN_9102 = 14'h238e == index ? 14'h281 : _GEN_9101;
  wire [13:0] _GEN_9103 = 14'h238f == index ? 14'h20b : _GEN_9102;
  wire [13:0] _GEN_9104 = 14'h2390 == index ? 14'h207 : _GEN_9103;
  wire [13:0] _GEN_9105 = 14'h2391 == index ? 14'h203 : _GEN_9104;
  wire [13:0] _GEN_9106 = 14'h2392 == index ? 14'h191 : _GEN_9105;
  wire [13:0] _GEN_9107 = 14'h2393 == index ? 14'h18e : _GEN_9106;
  wire [13:0] _GEN_9108 = 14'h2394 == index ? 14'h18b : _GEN_9107;
  wire [13:0] _GEN_9109 = 14'h2395 == index ? 14'h188 : _GEN_9108;
  wire [13:0] _GEN_9110 = 14'h2396 == index ? 14'h185 : _GEN_9109;
  wire [13:0] _GEN_9111 = 14'h2397 == index ? 14'h182 : _GEN_9110;
  wire [13:0] _GEN_9112 = 14'h2398 == index ? 14'h117 : _GEN_9111;
  wire [13:0] _GEN_9113 = 14'h2399 == index ? 14'h115 : _GEN_9112;
  wire [13:0] _GEN_9114 = 14'h239a == index ? 14'h113 : _GEN_9113;
  wire [13:0] _GEN_9115 = 14'h239b == index ? 14'h111 : _GEN_9114;
  wire [13:0] _GEN_9116 = 14'h239c == index ? 14'h10f : _GEN_9115;
  wire [13:0] _GEN_9117 = 14'h239d == index ? 14'h10d : _GEN_9116;
  wire [13:0] _GEN_9118 = 14'h239e == index ? 14'h10b : _GEN_9117;
  wire [13:0] _GEN_9119 = 14'h239f == index ? 14'h109 : _GEN_9118;
  wire [13:0] _GEN_9120 = 14'h23a0 == index ? 14'h107 : _GEN_9119;
  wire [13:0] _GEN_9121 = 14'h23a1 == index ? 14'h105 : _GEN_9120;
  wire [13:0] _GEN_9122 = 14'h23a2 == index ? 14'h103 : _GEN_9121;
  wire [13:0] _GEN_9123 = 14'h23a3 == index ? 14'h101 : _GEN_9122;
  wire [13:0] _GEN_9124 = 14'h23a4 == index ? 14'ha3 : _GEN_9123;
  wire [13:0] _GEN_9125 = 14'h23a5 == index ? 14'ha2 : _GEN_9124;
  wire [13:0] _GEN_9126 = 14'h23a6 == index ? 14'ha1 : _GEN_9125;
  wire [13:0] _GEN_9127 = 14'h23a7 == index ? 14'ha0 : _GEN_9126;
  wire [13:0] _GEN_9128 = 14'h23a8 == index ? 14'h9f : _GEN_9127;
  wire [13:0] _GEN_9129 = 14'h23a9 == index ? 14'h9e : _GEN_9128;
  wire [13:0] _GEN_9130 = 14'h23aa == index ? 14'h9d : _GEN_9129;
  wire [13:0] _GEN_9131 = 14'h23ab == index ? 14'h9c : _GEN_9130;
  wire [13:0] _GEN_9132 = 14'h23ac == index ? 14'h9b : _GEN_9131;
  wire [13:0] _GEN_9133 = 14'h23ad == index ? 14'h9a : _GEN_9132;
  wire [13:0] _GEN_9134 = 14'h23ae == index ? 14'h99 : _GEN_9133;
  wire [13:0] _GEN_9135 = 14'h23af == index ? 14'h98 : _GEN_9134;
  wire [13:0] _GEN_9136 = 14'h23b0 == index ? 14'h97 : _GEN_9135;
  wire [13:0] _GEN_9137 = 14'h23b1 == index ? 14'h96 : _GEN_9136;
  wire [13:0] _GEN_9138 = 14'h23b2 == index ? 14'h95 : _GEN_9137;
  wire [13:0] _GEN_9139 = 14'h23b3 == index ? 14'h94 : _GEN_9138;
  wire [13:0] _GEN_9140 = 14'h23b4 == index ? 14'h93 : _GEN_9139;
  wire [13:0] _GEN_9141 = 14'h23b5 == index ? 14'h92 : _GEN_9140;
  wire [13:0] _GEN_9142 = 14'h23b6 == index ? 14'h91 : _GEN_9141;
  wire [13:0] _GEN_9143 = 14'h23b7 == index ? 14'h90 : _GEN_9142;
  wire [13:0] _GEN_9144 = 14'h23b8 == index ? 14'h8f : _GEN_9143;
  wire [13:0] _GEN_9145 = 14'h23b9 == index ? 14'h8e : _GEN_9144;
  wire [13:0] _GEN_9146 = 14'h23ba == index ? 14'h8d : _GEN_9145;
  wire [13:0] _GEN_9147 = 14'h23bb == index ? 14'h8c : _GEN_9146;
  wire [13:0] _GEN_9148 = 14'h23bc == index ? 14'h8b : _GEN_9147;
  wire [13:0] _GEN_9149 = 14'h23bd == index ? 14'h8a : _GEN_9148;
  wire [13:0] _GEN_9150 = 14'h23be == index ? 14'h89 : _GEN_9149;
  wire [13:0] _GEN_9151 = 14'h23bf == index ? 14'h88 : _GEN_9150;
  wire [13:0] _GEN_9152 = 14'h23c0 == index ? 14'h87 : _GEN_9151;
  wire [13:0] _GEN_9153 = 14'h23c1 == index ? 14'h86 : _GEN_9152;
  wire [13:0] _GEN_9154 = 14'h23c2 == index ? 14'h85 : _GEN_9153;
  wire [13:0] _GEN_9155 = 14'h23c3 == index ? 14'h84 : _GEN_9154;
  wire [13:0] _GEN_9156 = 14'h23c4 == index ? 14'h83 : _GEN_9155;
  wire [13:0] _GEN_9157 = 14'h23c5 == index ? 14'h82 : _GEN_9156;
  wire [13:0] _GEN_9158 = 14'h23c6 == index ? 14'h81 : _GEN_9157;
  wire [13:0] _GEN_9159 = 14'h23c7 == index ? 14'h80 : _GEN_9158;
  wire [13:0] _GEN_9160 = 14'h23c8 == index ? 14'h47 : _GEN_9159;
  wire [13:0] _GEN_9161 = 14'h23c9 == index ? 14'h47 : _GEN_9160;
  wire [13:0] _GEN_9162 = 14'h23ca == index ? 14'h47 : _GEN_9161;
  wire [13:0] _GEN_9163 = 14'h23cb == index ? 14'h47 : _GEN_9162;
  wire [13:0] _GEN_9164 = 14'h23cc == index ? 14'h47 : _GEN_9163;
  wire [13:0] _GEN_9165 = 14'h23cd == index ? 14'h47 : _GEN_9164;
  wire [13:0] _GEN_9166 = 14'h23ce == index ? 14'h47 : _GEN_9165;
  wire [13:0] _GEN_9167 = 14'h23cf == index ? 14'h47 : _GEN_9166;
  wire [13:0] _GEN_9168 = 14'h23d0 == index ? 14'h47 : _GEN_9167;
  wire [13:0] _GEN_9169 = 14'h23d1 == index ? 14'h47 : _GEN_9168;
  wire [13:0] _GEN_9170 = 14'h23d2 == index ? 14'h47 : _GEN_9169;
  wire [13:0] _GEN_9171 = 14'h23d3 == index ? 14'h47 : _GEN_9170;
  wire [13:0] _GEN_9172 = 14'h23d4 == index ? 14'h47 : _GEN_9171;
  wire [13:0] _GEN_9173 = 14'h23d5 == index ? 14'h47 : _GEN_9172;
  wire [13:0] _GEN_9174 = 14'h23d6 == index ? 14'h47 : _GEN_9173;
  wire [13:0] _GEN_9175 = 14'h23d7 == index ? 14'h47 : _GEN_9174;
  wire [13:0] _GEN_9176 = 14'h23d8 == index ? 14'h47 : _GEN_9175;
  wire [13:0] _GEN_9177 = 14'h23d9 == index ? 14'h47 : _GEN_9176;
  wire [13:0] _GEN_9178 = 14'h23da == index ? 14'h47 : _GEN_9177;
  wire [13:0] _GEN_9179 = 14'h23db == index ? 14'h47 : _GEN_9178;
  wire [13:0] _GEN_9180 = 14'h23dc == index ? 14'h47 : _GEN_9179;
  wire [13:0] _GEN_9181 = 14'h23dd == index ? 14'h47 : _GEN_9180;
  wire [13:0] _GEN_9182 = 14'h23de == index ? 14'h47 : _GEN_9181;
  wire [13:0] _GEN_9183 = 14'h23df == index ? 14'h47 : _GEN_9182;
  wire [13:0] _GEN_9184 = 14'h23e0 == index ? 14'h47 : _GEN_9183;
  wire [13:0] _GEN_9185 = 14'h23e1 == index ? 14'h47 : _GEN_9184;
  wire [13:0] _GEN_9186 = 14'h23e2 == index ? 14'h47 : _GEN_9185;
  wire [13:0] _GEN_9187 = 14'h23e3 == index ? 14'h47 : _GEN_9186;
  wire [13:0] _GEN_9188 = 14'h23e4 == index ? 14'h47 : _GEN_9187;
  wire [13:0] _GEN_9189 = 14'h23e5 == index ? 14'h47 : _GEN_9188;
  wire [13:0] _GEN_9190 = 14'h23e6 == index ? 14'h47 : _GEN_9189;
  wire [13:0] _GEN_9191 = 14'h23e7 == index ? 14'h47 : _GEN_9190;
  wire [13:0] _GEN_9192 = 14'h23e8 == index ? 14'h47 : _GEN_9191;
  wire [13:0] _GEN_9193 = 14'h23e9 == index ? 14'h47 : _GEN_9192;
  wire [13:0] _GEN_9194 = 14'h23ea == index ? 14'h47 : _GEN_9193;
  wire [13:0] _GEN_9195 = 14'h23eb == index ? 14'h47 : _GEN_9194;
  wire [13:0] _GEN_9196 = 14'h23ec == index ? 14'h47 : _GEN_9195;
  wire [13:0] _GEN_9197 = 14'h23ed == index ? 14'h47 : _GEN_9196;
  wire [13:0] _GEN_9198 = 14'h23ee == index ? 14'h47 : _GEN_9197;
  wire [13:0] _GEN_9199 = 14'h23ef == index ? 14'h47 : _GEN_9198;
  wire [13:0] _GEN_9200 = 14'h23f0 == index ? 14'h47 : _GEN_9199;
  wire [13:0] _GEN_9201 = 14'h23f1 == index ? 14'h47 : _GEN_9200;
  wire [13:0] _GEN_9202 = 14'h23f2 == index ? 14'h47 : _GEN_9201;
  wire [13:0] _GEN_9203 = 14'h23f3 == index ? 14'h47 : _GEN_9202;
  wire [13:0] _GEN_9204 = 14'h23f4 == index ? 14'h47 : _GEN_9203;
  wire [13:0] _GEN_9205 = 14'h23f5 == index ? 14'h47 : _GEN_9204;
  wire [13:0] _GEN_9206 = 14'h23f6 == index ? 14'h47 : _GEN_9205;
  wire [13:0] _GEN_9207 = 14'h23f7 == index ? 14'h47 : _GEN_9206;
  wire [13:0] _GEN_9208 = 14'h23f8 == index ? 14'h47 : _GEN_9207;
  wire [13:0] _GEN_9209 = 14'h23f9 == index ? 14'h47 : _GEN_9208;
  wire [13:0] _GEN_9210 = 14'h23fa == index ? 14'h47 : _GEN_9209;
  wire [13:0] _GEN_9211 = 14'h23fb == index ? 14'h47 : _GEN_9210;
  wire [13:0] _GEN_9212 = 14'h23fc == index ? 14'h47 : _GEN_9211;
  wire [13:0] _GEN_9213 = 14'h23fd == index ? 14'h47 : _GEN_9212;
  wire [13:0] _GEN_9214 = 14'h23fe == index ? 14'h47 : _GEN_9213;
  wire [13:0] _GEN_9215 = 14'h23ff == index ? 14'h47 : _GEN_9214;
  wire [13:0] _GEN_9216 = 14'h2400 == index ? 14'h0 : _GEN_9215;
  wire [13:0] _GEN_9217 = 14'h2401 == index ? 14'h2400 : _GEN_9216;
  wire [13:0] _GEN_9218 = 14'h2402 == index ? 14'h1200 : _GEN_9217;
  wire [13:0] _GEN_9219 = 14'h2403 == index ? 14'hc00 : _GEN_9218;
  wire [13:0] _GEN_9220 = 14'h2404 == index ? 14'h900 : _GEN_9219;
  wire [13:0] _GEN_9221 = 14'h2405 == index ? 14'h702 : _GEN_9220;
  wire [13:0] _GEN_9222 = 14'h2406 == index ? 14'h600 : _GEN_9221;
  wire [13:0] _GEN_9223 = 14'h2407 == index ? 14'h502 : _GEN_9222;
  wire [13:0] _GEN_9224 = 14'h2408 == index ? 14'h480 : _GEN_9223;
  wire [13:0] _GEN_9225 = 14'h2409 == index ? 14'h400 : _GEN_9224;
  wire [13:0] _GEN_9226 = 14'h240a == index ? 14'h382 : _GEN_9225;
  wire [13:0] _GEN_9227 = 14'h240b == index ? 14'h306 : _GEN_9226;
  wire [13:0] _GEN_9228 = 14'h240c == index ? 14'h300 : _GEN_9227;
  wire [13:0] _GEN_9229 = 14'h240d == index ? 14'h287 : _GEN_9228;
  wire [13:0] _GEN_9230 = 14'h240e == index ? 14'h282 : _GEN_9229;
  wire [13:0] _GEN_9231 = 14'h240f == index ? 14'h20c : _GEN_9230;
  wire [13:0] _GEN_9232 = 14'h2410 == index ? 14'h208 : _GEN_9231;
  wire [13:0] _GEN_9233 = 14'h2411 == index ? 14'h204 : _GEN_9232;
  wire [13:0] _GEN_9234 = 14'h2412 == index ? 14'h200 : _GEN_9233;
  wire [13:0] _GEN_9235 = 14'h2413 == index ? 14'h18f : _GEN_9234;
  wire [13:0] _GEN_9236 = 14'h2414 == index ? 14'h18c : _GEN_9235;
  wire [13:0] _GEN_9237 = 14'h2415 == index ? 14'h189 : _GEN_9236;
  wire [13:0] _GEN_9238 = 14'h2416 == index ? 14'h186 : _GEN_9237;
  wire [13:0] _GEN_9239 = 14'h2417 == index ? 14'h183 : _GEN_9238;
  wire [13:0] _GEN_9240 = 14'h2418 == index ? 14'h180 : _GEN_9239;
  wire [13:0] _GEN_9241 = 14'h2419 == index ? 14'h116 : _GEN_9240;
  wire [13:0] _GEN_9242 = 14'h241a == index ? 14'h114 : _GEN_9241;
  wire [13:0] _GEN_9243 = 14'h241b == index ? 14'h112 : _GEN_9242;
  wire [13:0] _GEN_9244 = 14'h241c == index ? 14'h110 : _GEN_9243;
  wire [13:0] _GEN_9245 = 14'h241d == index ? 14'h10e : _GEN_9244;
  wire [13:0] _GEN_9246 = 14'h241e == index ? 14'h10c : _GEN_9245;
  wire [13:0] _GEN_9247 = 14'h241f == index ? 14'h10a : _GEN_9246;
  wire [13:0] _GEN_9248 = 14'h2420 == index ? 14'h108 : _GEN_9247;
  wire [13:0] _GEN_9249 = 14'h2421 == index ? 14'h106 : _GEN_9248;
  wire [13:0] _GEN_9250 = 14'h2422 == index ? 14'h104 : _GEN_9249;
  wire [13:0] _GEN_9251 = 14'h2423 == index ? 14'h102 : _GEN_9250;
  wire [13:0] _GEN_9252 = 14'h2424 == index ? 14'h100 : _GEN_9251;
  wire [13:0] _GEN_9253 = 14'h2425 == index ? 14'ha3 : _GEN_9252;
  wire [13:0] _GEN_9254 = 14'h2426 == index ? 14'ha2 : _GEN_9253;
  wire [13:0] _GEN_9255 = 14'h2427 == index ? 14'ha1 : _GEN_9254;
  wire [13:0] _GEN_9256 = 14'h2428 == index ? 14'ha0 : _GEN_9255;
  wire [13:0] _GEN_9257 = 14'h2429 == index ? 14'h9f : _GEN_9256;
  wire [13:0] _GEN_9258 = 14'h242a == index ? 14'h9e : _GEN_9257;
  wire [13:0] _GEN_9259 = 14'h242b == index ? 14'h9d : _GEN_9258;
  wire [13:0] _GEN_9260 = 14'h242c == index ? 14'h9c : _GEN_9259;
  wire [13:0] _GEN_9261 = 14'h242d == index ? 14'h9b : _GEN_9260;
  wire [13:0] _GEN_9262 = 14'h242e == index ? 14'h9a : _GEN_9261;
  wire [13:0] _GEN_9263 = 14'h242f == index ? 14'h99 : _GEN_9262;
  wire [13:0] _GEN_9264 = 14'h2430 == index ? 14'h98 : _GEN_9263;
  wire [13:0] _GEN_9265 = 14'h2431 == index ? 14'h97 : _GEN_9264;
  wire [13:0] _GEN_9266 = 14'h2432 == index ? 14'h96 : _GEN_9265;
  wire [13:0] _GEN_9267 = 14'h2433 == index ? 14'h95 : _GEN_9266;
  wire [13:0] _GEN_9268 = 14'h2434 == index ? 14'h94 : _GEN_9267;
  wire [13:0] _GEN_9269 = 14'h2435 == index ? 14'h93 : _GEN_9268;
  wire [13:0] _GEN_9270 = 14'h2436 == index ? 14'h92 : _GEN_9269;
  wire [13:0] _GEN_9271 = 14'h2437 == index ? 14'h91 : _GEN_9270;
  wire [13:0] _GEN_9272 = 14'h2438 == index ? 14'h90 : _GEN_9271;
  wire [13:0] _GEN_9273 = 14'h2439 == index ? 14'h8f : _GEN_9272;
  wire [13:0] _GEN_9274 = 14'h243a == index ? 14'h8e : _GEN_9273;
  wire [13:0] _GEN_9275 = 14'h243b == index ? 14'h8d : _GEN_9274;
  wire [13:0] _GEN_9276 = 14'h243c == index ? 14'h8c : _GEN_9275;
  wire [13:0] _GEN_9277 = 14'h243d == index ? 14'h8b : _GEN_9276;
  wire [13:0] _GEN_9278 = 14'h243e == index ? 14'h8a : _GEN_9277;
  wire [13:0] _GEN_9279 = 14'h243f == index ? 14'h89 : _GEN_9278;
  wire [13:0] _GEN_9280 = 14'h2440 == index ? 14'h88 : _GEN_9279;
  wire [13:0] _GEN_9281 = 14'h2441 == index ? 14'h87 : _GEN_9280;
  wire [13:0] _GEN_9282 = 14'h2442 == index ? 14'h86 : _GEN_9281;
  wire [13:0] _GEN_9283 = 14'h2443 == index ? 14'h85 : _GEN_9282;
  wire [13:0] _GEN_9284 = 14'h2444 == index ? 14'h84 : _GEN_9283;
  wire [13:0] _GEN_9285 = 14'h2445 == index ? 14'h83 : _GEN_9284;
  wire [13:0] _GEN_9286 = 14'h2446 == index ? 14'h82 : _GEN_9285;
  wire [13:0] _GEN_9287 = 14'h2447 == index ? 14'h81 : _GEN_9286;
  wire [13:0] _GEN_9288 = 14'h2448 == index ? 14'h80 : _GEN_9287;
  wire [13:0] _GEN_9289 = 14'h2449 == index ? 14'h48 : _GEN_9288;
  wire [13:0] _GEN_9290 = 14'h244a == index ? 14'h48 : _GEN_9289;
  wire [13:0] _GEN_9291 = 14'h244b == index ? 14'h48 : _GEN_9290;
  wire [13:0] _GEN_9292 = 14'h244c == index ? 14'h48 : _GEN_9291;
  wire [13:0] _GEN_9293 = 14'h244d == index ? 14'h48 : _GEN_9292;
  wire [13:0] _GEN_9294 = 14'h244e == index ? 14'h48 : _GEN_9293;
  wire [13:0] _GEN_9295 = 14'h244f == index ? 14'h48 : _GEN_9294;
  wire [13:0] _GEN_9296 = 14'h2450 == index ? 14'h48 : _GEN_9295;
  wire [13:0] _GEN_9297 = 14'h2451 == index ? 14'h48 : _GEN_9296;
  wire [13:0] _GEN_9298 = 14'h2452 == index ? 14'h48 : _GEN_9297;
  wire [13:0] _GEN_9299 = 14'h2453 == index ? 14'h48 : _GEN_9298;
  wire [13:0] _GEN_9300 = 14'h2454 == index ? 14'h48 : _GEN_9299;
  wire [13:0] _GEN_9301 = 14'h2455 == index ? 14'h48 : _GEN_9300;
  wire [13:0] _GEN_9302 = 14'h2456 == index ? 14'h48 : _GEN_9301;
  wire [13:0] _GEN_9303 = 14'h2457 == index ? 14'h48 : _GEN_9302;
  wire [13:0] _GEN_9304 = 14'h2458 == index ? 14'h48 : _GEN_9303;
  wire [13:0] _GEN_9305 = 14'h2459 == index ? 14'h48 : _GEN_9304;
  wire [13:0] _GEN_9306 = 14'h245a == index ? 14'h48 : _GEN_9305;
  wire [13:0] _GEN_9307 = 14'h245b == index ? 14'h48 : _GEN_9306;
  wire [13:0] _GEN_9308 = 14'h245c == index ? 14'h48 : _GEN_9307;
  wire [13:0] _GEN_9309 = 14'h245d == index ? 14'h48 : _GEN_9308;
  wire [13:0] _GEN_9310 = 14'h245e == index ? 14'h48 : _GEN_9309;
  wire [13:0] _GEN_9311 = 14'h245f == index ? 14'h48 : _GEN_9310;
  wire [13:0] _GEN_9312 = 14'h2460 == index ? 14'h48 : _GEN_9311;
  wire [13:0] _GEN_9313 = 14'h2461 == index ? 14'h48 : _GEN_9312;
  wire [13:0] _GEN_9314 = 14'h2462 == index ? 14'h48 : _GEN_9313;
  wire [13:0] _GEN_9315 = 14'h2463 == index ? 14'h48 : _GEN_9314;
  wire [13:0] _GEN_9316 = 14'h2464 == index ? 14'h48 : _GEN_9315;
  wire [13:0] _GEN_9317 = 14'h2465 == index ? 14'h48 : _GEN_9316;
  wire [13:0] _GEN_9318 = 14'h2466 == index ? 14'h48 : _GEN_9317;
  wire [13:0] _GEN_9319 = 14'h2467 == index ? 14'h48 : _GEN_9318;
  wire [13:0] _GEN_9320 = 14'h2468 == index ? 14'h48 : _GEN_9319;
  wire [13:0] _GEN_9321 = 14'h2469 == index ? 14'h48 : _GEN_9320;
  wire [13:0] _GEN_9322 = 14'h246a == index ? 14'h48 : _GEN_9321;
  wire [13:0] _GEN_9323 = 14'h246b == index ? 14'h48 : _GEN_9322;
  wire [13:0] _GEN_9324 = 14'h246c == index ? 14'h48 : _GEN_9323;
  wire [13:0] _GEN_9325 = 14'h246d == index ? 14'h48 : _GEN_9324;
  wire [13:0] _GEN_9326 = 14'h246e == index ? 14'h48 : _GEN_9325;
  wire [13:0] _GEN_9327 = 14'h246f == index ? 14'h48 : _GEN_9326;
  wire [13:0] _GEN_9328 = 14'h2470 == index ? 14'h48 : _GEN_9327;
  wire [13:0] _GEN_9329 = 14'h2471 == index ? 14'h48 : _GEN_9328;
  wire [13:0] _GEN_9330 = 14'h2472 == index ? 14'h48 : _GEN_9329;
  wire [13:0] _GEN_9331 = 14'h2473 == index ? 14'h48 : _GEN_9330;
  wire [13:0] _GEN_9332 = 14'h2474 == index ? 14'h48 : _GEN_9331;
  wire [13:0] _GEN_9333 = 14'h2475 == index ? 14'h48 : _GEN_9332;
  wire [13:0] _GEN_9334 = 14'h2476 == index ? 14'h48 : _GEN_9333;
  wire [13:0] _GEN_9335 = 14'h2477 == index ? 14'h48 : _GEN_9334;
  wire [13:0] _GEN_9336 = 14'h2478 == index ? 14'h48 : _GEN_9335;
  wire [13:0] _GEN_9337 = 14'h2479 == index ? 14'h48 : _GEN_9336;
  wire [13:0] _GEN_9338 = 14'h247a == index ? 14'h48 : _GEN_9337;
  wire [13:0] _GEN_9339 = 14'h247b == index ? 14'h48 : _GEN_9338;
  wire [13:0] _GEN_9340 = 14'h247c == index ? 14'h48 : _GEN_9339;
  wire [13:0] _GEN_9341 = 14'h247d == index ? 14'h48 : _GEN_9340;
  wire [13:0] _GEN_9342 = 14'h247e == index ? 14'h48 : _GEN_9341;
  wire [13:0] _GEN_9343 = 14'h247f == index ? 14'h48 : _GEN_9342;
  wire [13:0] _GEN_9344 = 14'h2480 == index ? 14'h0 : _GEN_9343;
  wire [13:0] _GEN_9345 = 14'h2481 == index ? 14'h2480 : _GEN_9344;
  wire [13:0] _GEN_9346 = 14'h2482 == index ? 14'h1201 : _GEN_9345;
  wire [13:0] _GEN_9347 = 14'h2483 == index ? 14'hc01 : _GEN_9346;
  wire [13:0] _GEN_9348 = 14'h2484 == index ? 14'h901 : _GEN_9347;
  wire [13:0] _GEN_9349 = 14'h2485 == index ? 14'h703 : _GEN_9348;
  wire [13:0] _GEN_9350 = 14'h2486 == index ? 14'h601 : _GEN_9349;
  wire [13:0] _GEN_9351 = 14'h2487 == index ? 14'h503 : _GEN_9350;
  wire [13:0] _GEN_9352 = 14'h2488 == index ? 14'h481 : _GEN_9351;
  wire [13:0] _GEN_9353 = 14'h2489 == index ? 14'h401 : _GEN_9352;
  wire [13:0] _GEN_9354 = 14'h248a == index ? 14'h383 : _GEN_9353;
  wire [13:0] _GEN_9355 = 14'h248b == index ? 14'h307 : _GEN_9354;
  wire [13:0] _GEN_9356 = 14'h248c == index ? 14'h301 : _GEN_9355;
  wire [13:0] _GEN_9357 = 14'h248d == index ? 14'h288 : _GEN_9356;
  wire [13:0] _GEN_9358 = 14'h248e == index ? 14'h283 : _GEN_9357;
  wire [13:0] _GEN_9359 = 14'h248f == index ? 14'h20d : _GEN_9358;
  wire [13:0] _GEN_9360 = 14'h2490 == index ? 14'h209 : _GEN_9359;
  wire [13:0] _GEN_9361 = 14'h2491 == index ? 14'h205 : _GEN_9360;
  wire [13:0] _GEN_9362 = 14'h2492 == index ? 14'h201 : _GEN_9361;
  wire [13:0] _GEN_9363 = 14'h2493 == index ? 14'h190 : _GEN_9362;
  wire [13:0] _GEN_9364 = 14'h2494 == index ? 14'h18d : _GEN_9363;
  wire [13:0] _GEN_9365 = 14'h2495 == index ? 14'h18a : _GEN_9364;
  wire [13:0] _GEN_9366 = 14'h2496 == index ? 14'h187 : _GEN_9365;
  wire [13:0] _GEN_9367 = 14'h2497 == index ? 14'h184 : _GEN_9366;
  wire [13:0] _GEN_9368 = 14'h2498 == index ? 14'h181 : _GEN_9367;
  wire [13:0] _GEN_9369 = 14'h2499 == index ? 14'h117 : _GEN_9368;
  wire [13:0] _GEN_9370 = 14'h249a == index ? 14'h115 : _GEN_9369;
  wire [13:0] _GEN_9371 = 14'h249b == index ? 14'h113 : _GEN_9370;
  wire [13:0] _GEN_9372 = 14'h249c == index ? 14'h111 : _GEN_9371;
  wire [13:0] _GEN_9373 = 14'h249d == index ? 14'h10f : _GEN_9372;
  wire [13:0] _GEN_9374 = 14'h249e == index ? 14'h10d : _GEN_9373;
  wire [13:0] _GEN_9375 = 14'h249f == index ? 14'h10b : _GEN_9374;
  wire [13:0] _GEN_9376 = 14'h24a0 == index ? 14'h109 : _GEN_9375;
  wire [13:0] _GEN_9377 = 14'h24a1 == index ? 14'h107 : _GEN_9376;
  wire [13:0] _GEN_9378 = 14'h24a2 == index ? 14'h105 : _GEN_9377;
  wire [13:0] _GEN_9379 = 14'h24a3 == index ? 14'h103 : _GEN_9378;
  wire [13:0] _GEN_9380 = 14'h24a4 == index ? 14'h101 : _GEN_9379;
  wire [13:0] _GEN_9381 = 14'h24a5 == index ? 14'ha4 : _GEN_9380;
  wire [13:0] _GEN_9382 = 14'h24a6 == index ? 14'ha3 : _GEN_9381;
  wire [13:0] _GEN_9383 = 14'h24a7 == index ? 14'ha2 : _GEN_9382;
  wire [13:0] _GEN_9384 = 14'h24a8 == index ? 14'ha1 : _GEN_9383;
  wire [13:0] _GEN_9385 = 14'h24a9 == index ? 14'ha0 : _GEN_9384;
  wire [13:0] _GEN_9386 = 14'h24aa == index ? 14'h9f : _GEN_9385;
  wire [13:0] _GEN_9387 = 14'h24ab == index ? 14'h9e : _GEN_9386;
  wire [13:0] _GEN_9388 = 14'h24ac == index ? 14'h9d : _GEN_9387;
  wire [13:0] _GEN_9389 = 14'h24ad == index ? 14'h9c : _GEN_9388;
  wire [13:0] _GEN_9390 = 14'h24ae == index ? 14'h9b : _GEN_9389;
  wire [13:0] _GEN_9391 = 14'h24af == index ? 14'h9a : _GEN_9390;
  wire [13:0] _GEN_9392 = 14'h24b0 == index ? 14'h99 : _GEN_9391;
  wire [13:0] _GEN_9393 = 14'h24b1 == index ? 14'h98 : _GEN_9392;
  wire [13:0] _GEN_9394 = 14'h24b2 == index ? 14'h97 : _GEN_9393;
  wire [13:0] _GEN_9395 = 14'h24b3 == index ? 14'h96 : _GEN_9394;
  wire [13:0] _GEN_9396 = 14'h24b4 == index ? 14'h95 : _GEN_9395;
  wire [13:0] _GEN_9397 = 14'h24b5 == index ? 14'h94 : _GEN_9396;
  wire [13:0] _GEN_9398 = 14'h24b6 == index ? 14'h93 : _GEN_9397;
  wire [13:0] _GEN_9399 = 14'h24b7 == index ? 14'h92 : _GEN_9398;
  wire [13:0] _GEN_9400 = 14'h24b8 == index ? 14'h91 : _GEN_9399;
  wire [13:0] _GEN_9401 = 14'h24b9 == index ? 14'h90 : _GEN_9400;
  wire [13:0] _GEN_9402 = 14'h24ba == index ? 14'h8f : _GEN_9401;
  wire [13:0] _GEN_9403 = 14'h24bb == index ? 14'h8e : _GEN_9402;
  wire [13:0] _GEN_9404 = 14'h24bc == index ? 14'h8d : _GEN_9403;
  wire [13:0] _GEN_9405 = 14'h24bd == index ? 14'h8c : _GEN_9404;
  wire [13:0] _GEN_9406 = 14'h24be == index ? 14'h8b : _GEN_9405;
  wire [13:0] _GEN_9407 = 14'h24bf == index ? 14'h8a : _GEN_9406;
  wire [13:0] _GEN_9408 = 14'h24c0 == index ? 14'h89 : _GEN_9407;
  wire [13:0] _GEN_9409 = 14'h24c1 == index ? 14'h88 : _GEN_9408;
  wire [13:0] _GEN_9410 = 14'h24c2 == index ? 14'h87 : _GEN_9409;
  wire [13:0] _GEN_9411 = 14'h24c3 == index ? 14'h86 : _GEN_9410;
  wire [13:0] _GEN_9412 = 14'h24c4 == index ? 14'h85 : _GEN_9411;
  wire [13:0] _GEN_9413 = 14'h24c5 == index ? 14'h84 : _GEN_9412;
  wire [13:0] _GEN_9414 = 14'h24c6 == index ? 14'h83 : _GEN_9413;
  wire [13:0] _GEN_9415 = 14'h24c7 == index ? 14'h82 : _GEN_9414;
  wire [13:0] _GEN_9416 = 14'h24c8 == index ? 14'h81 : _GEN_9415;
  wire [13:0] _GEN_9417 = 14'h24c9 == index ? 14'h80 : _GEN_9416;
  wire [13:0] _GEN_9418 = 14'h24ca == index ? 14'h49 : _GEN_9417;
  wire [13:0] _GEN_9419 = 14'h24cb == index ? 14'h49 : _GEN_9418;
  wire [13:0] _GEN_9420 = 14'h24cc == index ? 14'h49 : _GEN_9419;
  wire [13:0] _GEN_9421 = 14'h24cd == index ? 14'h49 : _GEN_9420;
  wire [13:0] _GEN_9422 = 14'h24ce == index ? 14'h49 : _GEN_9421;
  wire [13:0] _GEN_9423 = 14'h24cf == index ? 14'h49 : _GEN_9422;
  wire [13:0] _GEN_9424 = 14'h24d0 == index ? 14'h49 : _GEN_9423;
  wire [13:0] _GEN_9425 = 14'h24d1 == index ? 14'h49 : _GEN_9424;
  wire [13:0] _GEN_9426 = 14'h24d2 == index ? 14'h49 : _GEN_9425;
  wire [13:0] _GEN_9427 = 14'h24d3 == index ? 14'h49 : _GEN_9426;
  wire [13:0] _GEN_9428 = 14'h24d4 == index ? 14'h49 : _GEN_9427;
  wire [13:0] _GEN_9429 = 14'h24d5 == index ? 14'h49 : _GEN_9428;
  wire [13:0] _GEN_9430 = 14'h24d6 == index ? 14'h49 : _GEN_9429;
  wire [13:0] _GEN_9431 = 14'h24d7 == index ? 14'h49 : _GEN_9430;
  wire [13:0] _GEN_9432 = 14'h24d8 == index ? 14'h49 : _GEN_9431;
  wire [13:0] _GEN_9433 = 14'h24d9 == index ? 14'h49 : _GEN_9432;
  wire [13:0] _GEN_9434 = 14'h24da == index ? 14'h49 : _GEN_9433;
  wire [13:0] _GEN_9435 = 14'h24db == index ? 14'h49 : _GEN_9434;
  wire [13:0] _GEN_9436 = 14'h24dc == index ? 14'h49 : _GEN_9435;
  wire [13:0] _GEN_9437 = 14'h24dd == index ? 14'h49 : _GEN_9436;
  wire [13:0] _GEN_9438 = 14'h24de == index ? 14'h49 : _GEN_9437;
  wire [13:0] _GEN_9439 = 14'h24df == index ? 14'h49 : _GEN_9438;
  wire [13:0] _GEN_9440 = 14'h24e0 == index ? 14'h49 : _GEN_9439;
  wire [13:0] _GEN_9441 = 14'h24e1 == index ? 14'h49 : _GEN_9440;
  wire [13:0] _GEN_9442 = 14'h24e2 == index ? 14'h49 : _GEN_9441;
  wire [13:0] _GEN_9443 = 14'h24e3 == index ? 14'h49 : _GEN_9442;
  wire [13:0] _GEN_9444 = 14'h24e4 == index ? 14'h49 : _GEN_9443;
  wire [13:0] _GEN_9445 = 14'h24e5 == index ? 14'h49 : _GEN_9444;
  wire [13:0] _GEN_9446 = 14'h24e6 == index ? 14'h49 : _GEN_9445;
  wire [13:0] _GEN_9447 = 14'h24e7 == index ? 14'h49 : _GEN_9446;
  wire [13:0] _GEN_9448 = 14'h24e8 == index ? 14'h49 : _GEN_9447;
  wire [13:0] _GEN_9449 = 14'h24e9 == index ? 14'h49 : _GEN_9448;
  wire [13:0] _GEN_9450 = 14'h24ea == index ? 14'h49 : _GEN_9449;
  wire [13:0] _GEN_9451 = 14'h24eb == index ? 14'h49 : _GEN_9450;
  wire [13:0] _GEN_9452 = 14'h24ec == index ? 14'h49 : _GEN_9451;
  wire [13:0] _GEN_9453 = 14'h24ed == index ? 14'h49 : _GEN_9452;
  wire [13:0] _GEN_9454 = 14'h24ee == index ? 14'h49 : _GEN_9453;
  wire [13:0] _GEN_9455 = 14'h24ef == index ? 14'h49 : _GEN_9454;
  wire [13:0] _GEN_9456 = 14'h24f0 == index ? 14'h49 : _GEN_9455;
  wire [13:0] _GEN_9457 = 14'h24f1 == index ? 14'h49 : _GEN_9456;
  wire [13:0] _GEN_9458 = 14'h24f2 == index ? 14'h49 : _GEN_9457;
  wire [13:0] _GEN_9459 = 14'h24f3 == index ? 14'h49 : _GEN_9458;
  wire [13:0] _GEN_9460 = 14'h24f4 == index ? 14'h49 : _GEN_9459;
  wire [13:0] _GEN_9461 = 14'h24f5 == index ? 14'h49 : _GEN_9460;
  wire [13:0] _GEN_9462 = 14'h24f6 == index ? 14'h49 : _GEN_9461;
  wire [13:0] _GEN_9463 = 14'h24f7 == index ? 14'h49 : _GEN_9462;
  wire [13:0] _GEN_9464 = 14'h24f8 == index ? 14'h49 : _GEN_9463;
  wire [13:0] _GEN_9465 = 14'h24f9 == index ? 14'h49 : _GEN_9464;
  wire [13:0] _GEN_9466 = 14'h24fa == index ? 14'h49 : _GEN_9465;
  wire [13:0] _GEN_9467 = 14'h24fb == index ? 14'h49 : _GEN_9466;
  wire [13:0] _GEN_9468 = 14'h24fc == index ? 14'h49 : _GEN_9467;
  wire [13:0] _GEN_9469 = 14'h24fd == index ? 14'h49 : _GEN_9468;
  wire [13:0] _GEN_9470 = 14'h24fe == index ? 14'h49 : _GEN_9469;
  wire [13:0] _GEN_9471 = 14'h24ff == index ? 14'h49 : _GEN_9470;
  wire [13:0] _GEN_9472 = 14'h2500 == index ? 14'h0 : _GEN_9471;
  wire [13:0] _GEN_9473 = 14'h2501 == index ? 14'h2500 : _GEN_9472;
  wire [13:0] _GEN_9474 = 14'h2502 == index ? 14'h1280 : _GEN_9473;
  wire [13:0] _GEN_9475 = 14'h2503 == index ? 14'hc02 : _GEN_9474;
  wire [13:0] _GEN_9476 = 14'h2504 == index ? 14'h902 : _GEN_9475;
  wire [13:0] _GEN_9477 = 14'h2505 == index ? 14'h704 : _GEN_9476;
  wire [13:0] _GEN_9478 = 14'h2506 == index ? 14'h602 : _GEN_9477;
  wire [13:0] _GEN_9479 = 14'h2507 == index ? 14'h504 : _GEN_9478;
  wire [13:0] _GEN_9480 = 14'h2508 == index ? 14'h482 : _GEN_9479;
  wire [13:0] _GEN_9481 = 14'h2509 == index ? 14'h402 : _GEN_9480;
  wire [13:0] _GEN_9482 = 14'h250a == index ? 14'h384 : _GEN_9481;
  wire [13:0] _GEN_9483 = 14'h250b == index ? 14'h308 : _GEN_9482;
  wire [13:0] _GEN_9484 = 14'h250c == index ? 14'h302 : _GEN_9483;
  wire [13:0] _GEN_9485 = 14'h250d == index ? 14'h289 : _GEN_9484;
  wire [13:0] _GEN_9486 = 14'h250e == index ? 14'h284 : _GEN_9485;
  wire [13:0] _GEN_9487 = 14'h250f == index ? 14'h20e : _GEN_9486;
  wire [13:0] _GEN_9488 = 14'h2510 == index ? 14'h20a : _GEN_9487;
  wire [13:0] _GEN_9489 = 14'h2511 == index ? 14'h206 : _GEN_9488;
  wire [13:0] _GEN_9490 = 14'h2512 == index ? 14'h202 : _GEN_9489;
  wire [13:0] _GEN_9491 = 14'h2513 == index ? 14'h191 : _GEN_9490;
  wire [13:0] _GEN_9492 = 14'h2514 == index ? 14'h18e : _GEN_9491;
  wire [13:0] _GEN_9493 = 14'h2515 == index ? 14'h18b : _GEN_9492;
  wire [13:0] _GEN_9494 = 14'h2516 == index ? 14'h188 : _GEN_9493;
  wire [13:0] _GEN_9495 = 14'h2517 == index ? 14'h185 : _GEN_9494;
  wire [13:0] _GEN_9496 = 14'h2518 == index ? 14'h182 : _GEN_9495;
  wire [13:0] _GEN_9497 = 14'h2519 == index ? 14'h118 : _GEN_9496;
  wire [13:0] _GEN_9498 = 14'h251a == index ? 14'h116 : _GEN_9497;
  wire [13:0] _GEN_9499 = 14'h251b == index ? 14'h114 : _GEN_9498;
  wire [13:0] _GEN_9500 = 14'h251c == index ? 14'h112 : _GEN_9499;
  wire [13:0] _GEN_9501 = 14'h251d == index ? 14'h110 : _GEN_9500;
  wire [13:0] _GEN_9502 = 14'h251e == index ? 14'h10e : _GEN_9501;
  wire [13:0] _GEN_9503 = 14'h251f == index ? 14'h10c : _GEN_9502;
  wire [13:0] _GEN_9504 = 14'h2520 == index ? 14'h10a : _GEN_9503;
  wire [13:0] _GEN_9505 = 14'h2521 == index ? 14'h108 : _GEN_9504;
  wire [13:0] _GEN_9506 = 14'h2522 == index ? 14'h106 : _GEN_9505;
  wire [13:0] _GEN_9507 = 14'h2523 == index ? 14'h104 : _GEN_9506;
  wire [13:0] _GEN_9508 = 14'h2524 == index ? 14'h102 : _GEN_9507;
  wire [13:0] _GEN_9509 = 14'h2525 == index ? 14'h100 : _GEN_9508;
  wire [13:0] _GEN_9510 = 14'h2526 == index ? 14'ha4 : _GEN_9509;
  wire [13:0] _GEN_9511 = 14'h2527 == index ? 14'ha3 : _GEN_9510;
  wire [13:0] _GEN_9512 = 14'h2528 == index ? 14'ha2 : _GEN_9511;
  wire [13:0] _GEN_9513 = 14'h2529 == index ? 14'ha1 : _GEN_9512;
  wire [13:0] _GEN_9514 = 14'h252a == index ? 14'ha0 : _GEN_9513;
  wire [13:0] _GEN_9515 = 14'h252b == index ? 14'h9f : _GEN_9514;
  wire [13:0] _GEN_9516 = 14'h252c == index ? 14'h9e : _GEN_9515;
  wire [13:0] _GEN_9517 = 14'h252d == index ? 14'h9d : _GEN_9516;
  wire [13:0] _GEN_9518 = 14'h252e == index ? 14'h9c : _GEN_9517;
  wire [13:0] _GEN_9519 = 14'h252f == index ? 14'h9b : _GEN_9518;
  wire [13:0] _GEN_9520 = 14'h2530 == index ? 14'h9a : _GEN_9519;
  wire [13:0] _GEN_9521 = 14'h2531 == index ? 14'h99 : _GEN_9520;
  wire [13:0] _GEN_9522 = 14'h2532 == index ? 14'h98 : _GEN_9521;
  wire [13:0] _GEN_9523 = 14'h2533 == index ? 14'h97 : _GEN_9522;
  wire [13:0] _GEN_9524 = 14'h2534 == index ? 14'h96 : _GEN_9523;
  wire [13:0] _GEN_9525 = 14'h2535 == index ? 14'h95 : _GEN_9524;
  wire [13:0] _GEN_9526 = 14'h2536 == index ? 14'h94 : _GEN_9525;
  wire [13:0] _GEN_9527 = 14'h2537 == index ? 14'h93 : _GEN_9526;
  wire [13:0] _GEN_9528 = 14'h2538 == index ? 14'h92 : _GEN_9527;
  wire [13:0] _GEN_9529 = 14'h2539 == index ? 14'h91 : _GEN_9528;
  wire [13:0] _GEN_9530 = 14'h253a == index ? 14'h90 : _GEN_9529;
  wire [13:0] _GEN_9531 = 14'h253b == index ? 14'h8f : _GEN_9530;
  wire [13:0] _GEN_9532 = 14'h253c == index ? 14'h8e : _GEN_9531;
  wire [13:0] _GEN_9533 = 14'h253d == index ? 14'h8d : _GEN_9532;
  wire [13:0] _GEN_9534 = 14'h253e == index ? 14'h8c : _GEN_9533;
  wire [13:0] _GEN_9535 = 14'h253f == index ? 14'h8b : _GEN_9534;
  wire [13:0] _GEN_9536 = 14'h2540 == index ? 14'h8a : _GEN_9535;
  wire [13:0] _GEN_9537 = 14'h2541 == index ? 14'h89 : _GEN_9536;
  wire [13:0] _GEN_9538 = 14'h2542 == index ? 14'h88 : _GEN_9537;
  wire [13:0] _GEN_9539 = 14'h2543 == index ? 14'h87 : _GEN_9538;
  wire [13:0] _GEN_9540 = 14'h2544 == index ? 14'h86 : _GEN_9539;
  wire [13:0] _GEN_9541 = 14'h2545 == index ? 14'h85 : _GEN_9540;
  wire [13:0] _GEN_9542 = 14'h2546 == index ? 14'h84 : _GEN_9541;
  wire [13:0] _GEN_9543 = 14'h2547 == index ? 14'h83 : _GEN_9542;
  wire [13:0] _GEN_9544 = 14'h2548 == index ? 14'h82 : _GEN_9543;
  wire [13:0] _GEN_9545 = 14'h2549 == index ? 14'h81 : _GEN_9544;
  wire [13:0] _GEN_9546 = 14'h254a == index ? 14'h80 : _GEN_9545;
  wire [13:0] _GEN_9547 = 14'h254b == index ? 14'h4a : _GEN_9546;
  wire [13:0] _GEN_9548 = 14'h254c == index ? 14'h4a : _GEN_9547;
  wire [13:0] _GEN_9549 = 14'h254d == index ? 14'h4a : _GEN_9548;
  wire [13:0] _GEN_9550 = 14'h254e == index ? 14'h4a : _GEN_9549;
  wire [13:0] _GEN_9551 = 14'h254f == index ? 14'h4a : _GEN_9550;
  wire [13:0] _GEN_9552 = 14'h2550 == index ? 14'h4a : _GEN_9551;
  wire [13:0] _GEN_9553 = 14'h2551 == index ? 14'h4a : _GEN_9552;
  wire [13:0] _GEN_9554 = 14'h2552 == index ? 14'h4a : _GEN_9553;
  wire [13:0] _GEN_9555 = 14'h2553 == index ? 14'h4a : _GEN_9554;
  wire [13:0] _GEN_9556 = 14'h2554 == index ? 14'h4a : _GEN_9555;
  wire [13:0] _GEN_9557 = 14'h2555 == index ? 14'h4a : _GEN_9556;
  wire [13:0] _GEN_9558 = 14'h2556 == index ? 14'h4a : _GEN_9557;
  wire [13:0] _GEN_9559 = 14'h2557 == index ? 14'h4a : _GEN_9558;
  wire [13:0] _GEN_9560 = 14'h2558 == index ? 14'h4a : _GEN_9559;
  wire [13:0] _GEN_9561 = 14'h2559 == index ? 14'h4a : _GEN_9560;
  wire [13:0] _GEN_9562 = 14'h255a == index ? 14'h4a : _GEN_9561;
  wire [13:0] _GEN_9563 = 14'h255b == index ? 14'h4a : _GEN_9562;
  wire [13:0] _GEN_9564 = 14'h255c == index ? 14'h4a : _GEN_9563;
  wire [13:0] _GEN_9565 = 14'h255d == index ? 14'h4a : _GEN_9564;
  wire [13:0] _GEN_9566 = 14'h255e == index ? 14'h4a : _GEN_9565;
  wire [13:0] _GEN_9567 = 14'h255f == index ? 14'h4a : _GEN_9566;
  wire [13:0] _GEN_9568 = 14'h2560 == index ? 14'h4a : _GEN_9567;
  wire [13:0] _GEN_9569 = 14'h2561 == index ? 14'h4a : _GEN_9568;
  wire [13:0] _GEN_9570 = 14'h2562 == index ? 14'h4a : _GEN_9569;
  wire [13:0] _GEN_9571 = 14'h2563 == index ? 14'h4a : _GEN_9570;
  wire [13:0] _GEN_9572 = 14'h2564 == index ? 14'h4a : _GEN_9571;
  wire [13:0] _GEN_9573 = 14'h2565 == index ? 14'h4a : _GEN_9572;
  wire [13:0] _GEN_9574 = 14'h2566 == index ? 14'h4a : _GEN_9573;
  wire [13:0] _GEN_9575 = 14'h2567 == index ? 14'h4a : _GEN_9574;
  wire [13:0] _GEN_9576 = 14'h2568 == index ? 14'h4a : _GEN_9575;
  wire [13:0] _GEN_9577 = 14'h2569 == index ? 14'h4a : _GEN_9576;
  wire [13:0] _GEN_9578 = 14'h256a == index ? 14'h4a : _GEN_9577;
  wire [13:0] _GEN_9579 = 14'h256b == index ? 14'h4a : _GEN_9578;
  wire [13:0] _GEN_9580 = 14'h256c == index ? 14'h4a : _GEN_9579;
  wire [13:0] _GEN_9581 = 14'h256d == index ? 14'h4a : _GEN_9580;
  wire [13:0] _GEN_9582 = 14'h256e == index ? 14'h4a : _GEN_9581;
  wire [13:0] _GEN_9583 = 14'h256f == index ? 14'h4a : _GEN_9582;
  wire [13:0] _GEN_9584 = 14'h2570 == index ? 14'h4a : _GEN_9583;
  wire [13:0] _GEN_9585 = 14'h2571 == index ? 14'h4a : _GEN_9584;
  wire [13:0] _GEN_9586 = 14'h2572 == index ? 14'h4a : _GEN_9585;
  wire [13:0] _GEN_9587 = 14'h2573 == index ? 14'h4a : _GEN_9586;
  wire [13:0] _GEN_9588 = 14'h2574 == index ? 14'h4a : _GEN_9587;
  wire [13:0] _GEN_9589 = 14'h2575 == index ? 14'h4a : _GEN_9588;
  wire [13:0] _GEN_9590 = 14'h2576 == index ? 14'h4a : _GEN_9589;
  wire [13:0] _GEN_9591 = 14'h2577 == index ? 14'h4a : _GEN_9590;
  wire [13:0] _GEN_9592 = 14'h2578 == index ? 14'h4a : _GEN_9591;
  wire [13:0] _GEN_9593 = 14'h2579 == index ? 14'h4a : _GEN_9592;
  wire [13:0] _GEN_9594 = 14'h257a == index ? 14'h4a : _GEN_9593;
  wire [13:0] _GEN_9595 = 14'h257b == index ? 14'h4a : _GEN_9594;
  wire [13:0] _GEN_9596 = 14'h257c == index ? 14'h4a : _GEN_9595;
  wire [13:0] _GEN_9597 = 14'h257d == index ? 14'h4a : _GEN_9596;
  wire [13:0] _GEN_9598 = 14'h257e == index ? 14'h4a : _GEN_9597;
  wire [13:0] _GEN_9599 = 14'h257f == index ? 14'h4a : _GEN_9598;
  wire [13:0] _GEN_9600 = 14'h2580 == index ? 14'h0 : _GEN_9599;
  wire [13:0] _GEN_9601 = 14'h2581 == index ? 14'h2580 : _GEN_9600;
  wire [13:0] _GEN_9602 = 14'h2582 == index ? 14'h1281 : _GEN_9601;
  wire [13:0] _GEN_9603 = 14'h2583 == index ? 14'hc80 : _GEN_9602;
  wire [13:0] _GEN_9604 = 14'h2584 == index ? 14'h903 : _GEN_9603;
  wire [13:0] _GEN_9605 = 14'h2585 == index ? 14'h780 : _GEN_9604;
  wire [13:0] _GEN_9606 = 14'h2586 == index ? 14'h603 : _GEN_9605;
  wire [13:0] _GEN_9607 = 14'h2587 == index ? 14'h505 : _GEN_9606;
  wire [13:0] _GEN_9608 = 14'h2588 == index ? 14'h483 : _GEN_9607;
  wire [13:0] _GEN_9609 = 14'h2589 == index ? 14'h403 : _GEN_9608;
  wire [13:0] _GEN_9610 = 14'h258a == index ? 14'h385 : _GEN_9609;
  wire [13:0] _GEN_9611 = 14'h258b == index ? 14'h309 : _GEN_9610;
  wire [13:0] _GEN_9612 = 14'h258c == index ? 14'h303 : _GEN_9611;
  wire [13:0] _GEN_9613 = 14'h258d == index ? 14'h28a : _GEN_9612;
  wire [13:0] _GEN_9614 = 14'h258e == index ? 14'h285 : _GEN_9613;
  wire [13:0] _GEN_9615 = 14'h258f == index ? 14'h280 : _GEN_9614;
  wire [13:0] _GEN_9616 = 14'h2590 == index ? 14'h20b : _GEN_9615;
  wire [13:0] _GEN_9617 = 14'h2591 == index ? 14'h207 : _GEN_9616;
  wire [13:0] _GEN_9618 = 14'h2592 == index ? 14'h203 : _GEN_9617;
  wire [13:0] _GEN_9619 = 14'h2593 == index ? 14'h192 : _GEN_9618;
  wire [13:0] _GEN_9620 = 14'h2594 == index ? 14'h18f : _GEN_9619;
  wire [13:0] _GEN_9621 = 14'h2595 == index ? 14'h18c : _GEN_9620;
  wire [13:0] _GEN_9622 = 14'h2596 == index ? 14'h189 : _GEN_9621;
  wire [13:0] _GEN_9623 = 14'h2597 == index ? 14'h186 : _GEN_9622;
  wire [13:0] _GEN_9624 = 14'h2598 == index ? 14'h183 : _GEN_9623;
  wire [13:0] _GEN_9625 = 14'h2599 == index ? 14'h180 : _GEN_9624;
  wire [13:0] _GEN_9626 = 14'h259a == index ? 14'h117 : _GEN_9625;
  wire [13:0] _GEN_9627 = 14'h259b == index ? 14'h115 : _GEN_9626;
  wire [13:0] _GEN_9628 = 14'h259c == index ? 14'h113 : _GEN_9627;
  wire [13:0] _GEN_9629 = 14'h259d == index ? 14'h111 : _GEN_9628;
  wire [13:0] _GEN_9630 = 14'h259e == index ? 14'h10f : _GEN_9629;
  wire [13:0] _GEN_9631 = 14'h259f == index ? 14'h10d : _GEN_9630;
  wire [13:0] _GEN_9632 = 14'h25a0 == index ? 14'h10b : _GEN_9631;
  wire [13:0] _GEN_9633 = 14'h25a1 == index ? 14'h109 : _GEN_9632;
  wire [13:0] _GEN_9634 = 14'h25a2 == index ? 14'h107 : _GEN_9633;
  wire [13:0] _GEN_9635 = 14'h25a3 == index ? 14'h105 : _GEN_9634;
  wire [13:0] _GEN_9636 = 14'h25a4 == index ? 14'h103 : _GEN_9635;
  wire [13:0] _GEN_9637 = 14'h25a5 == index ? 14'h101 : _GEN_9636;
  wire [13:0] _GEN_9638 = 14'h25a6 == index ? 14'ha5 : _GEN_9637;
  wire [13:0] _GEN_9639 = 14'h25a7 == index ? 14'ha4 : _GEN_9638;
  wire [13:0] _GEN_9640 = 14'h25a8 == index ? 14'ha3 : _GEN_9639;
  wire [13:0] _GEN_9641 = 14'h25a9 == index ? 14'ha2 : _GEN_9640;
  wire [13:0] _GEN_9642 = 14'h25aa == index ? 14'ha1 : _GEN_9641;
  wire [13:0] _GEN_9643 = 14'h25ab == index ? 14'ha0 : _GEN_9642;
  wire [13:0] _GEN_9644 = 14'h25ac == index ? 14'h9f : _GEN_9643;
  wire [13:0] _GEN_9645 = 14'h25ad == index ? 14'h9e : _GEN_9644;
  wire [13:0] _GEN_9646 = 14'h25ae == index ? 14'h9d : _GEN_9645;
  wire [13:0] _GEN_9647 = 14'h25af == index ? 14'h9c : _GEN_9646;
  wire [13:0] _GEN_9648 = 14'h25b0 == index ? 14'h9b : _GEN_9647;
  wire [13:0] _GEN_9649 = 14'h25b1 == index ? 14'h9a : _GEN_9648;
  wire [13:0] _GEN_9650 = 14'h25b2 == index ? 14'h99 : _GEN_9649;
  wire [13:0] _GEN_9651 = 14'h25b3 == index ? 14'h98 : _GEN_9650;
  wire [13:0] _GEN_9652 = 14'h25b4 == index ? 14'h97 : _GEN_9651;
  wire [13:0] _GEN_9653 = 14'h25b5 == index ? 14'h96 : _GEN_9652;
  wire [13:0] _GEN_9654 = 14'h25b6 == index ? 14'h95 : _GEN_9653;
  wire [13:0] _GEN_9655 = 14'h25b7 == index ? 14'h94 : _GEN_9654;
  wire [13:0] _GEN_9656 = 14'h25b8 == index ? 14'h93 : _GEN_9655;
  wire [13:0] _GEN_9657 = 14'h25b9 == index ? 14'h92 : _GEN_9656;
  wire [13:0] _GEN_9658 = 14'h25ba == index ? 14'h91 : _GEN_9657;
  wire [13:0] _GEN_9659 = 14'h25bb == index ? 14'h90 : _GEN_9658;
  wire [13:0] _GEN_9660 = 14'h25bc == index ? 14'h8f : _GEN_9659;
  wire [13:0] _GEN_9661 = 14'h25bd == index ? 14'h8e : _GEN_9660;
  wire [13:0] _GEN_9662 = 14'h25be == index ? 14'h8d : _GEN_9661;
  wire [13:0] _GEN_9663 = 14'h25bf == index ? 14'h8c : _GEN_9662;
  wire [13:0] _GEN_9664 = 14'h25c0 == index ? 14'h8b : _GEN_9663;
  wire [13:0] _GEN_9665 = 14'h25c1 == index ? 14'h8a : _GEN_9664;
  wire [13:0] _GEN_9666 = 14'h25c2 == index ? 14'h89 : _GEN_9665;
  wire [13:0] _GEN_9667 = 14'h25c3 == index ? 14'h88 : _GEN_9666;
  wire [13:0] _GEN_9668 = 14'h25c4 == index ? 14'h87 : _GEN_9667;
  wire [13:0] _GEN_9669 = 14'h25c5 == index ? 14'h86 : _GEN_9668;
  wire [13:0] _GEN_9670 = 14'h25c6 == index ? 14'h85 : _GEN_9669;
  wire [13:0] _GEN_9671 = 14'h25c7 == index ? 14'h84 : _GEN_9670;
  wire [13:0] _GEN_9672 = 14'h25c8 == index ? 14'h83 : _GEN_9671;
  wire [13:0] _GEN_9673 = 14'h25c9 == index ? 14'h82 : _GEN_9672;
  wire [13:0] _GEN_9674 = 14'h25ca == index ? 14'h81 : _GEN_9673;
  wire [13:0] _GEN_9675 = 14'h25cb == index ? 14'h80 : _GEN_9674;
  wire [13:0] _GEN_9676 = 14'h25cc == index ? 14'h4b : _GEN_9675;
  wire [13:0] _GEN_9677 = 14'h25cd == index ? 14'h4b : _GEN_9676;
  wire [13:0] _GEN_9678 = 14'h25ce == index ? 14'h4b : _GEN_9677;
  wire [13:0] _GEN_9679 = 14'h25cf == index ? 14'h4b : _GEN_9678;
  wire [13:0] _GEN_9680 = 14'h25d0 == index ? 14'h4b : _GEN_9679;
  wire [13:0] _GEN_9681 = 14'h25d1 == index ? 14'h4b : _GEN_9680;
  wire [13:0] _GEN_9682 = 14'h25d2 == index ? 14'h4b : _GEN_9681;
  wire [13:0] _GEN_9683 = 14'h25d3 == index ? 14'h4b : _GEN_9682;
  wire [13:0] _GEN_9684 = 14'h25d4 == index ? 14'h4b : _GEN_9683;
  wire [13:0] _GEN_9685 = 14'h25d5 == index ? 14'h4b : _GEN_9684;
  wire [13:0] _GEN_9686 = 14'h25d6 == index ? 14'h4b : _GEN_9685;
  wire [13:0] _GEN_9687 = 14'h25d7 == index ? 14'h4b : _GEN_9686;
  wire [13:0] _GEN_9688 = 14'h25d8 == index ? 14'h4b : _GEN_9687;
  wire [13:0] _GEN_9689 = 14'h25d9 == index ? 14'h4b : _GEN_9688;
  wire [13:0] _GEN_9690 = 14'h25da == index ? 14'h4b : _GEN_9689;
  wire [13:0] _GEN_9691 = 14'h25db == index ? 14'h4b : _GEN_9690;
  wire [13:0] _GEN_9692 = 14'h25dc == index ? 14'h4b : _GEN_9691;
  wire [13:0] _GEN_9693 = 14'h25dd == index ? 14'h4b : _GEN_9692;
  wire [13:0] _GEN_9694 = 14'h25de == index ? 14'h4b : _GEN_9693;
  wire [13:0] _GEN_9695 = 14'h25df == index ? 14'h4b : _GEN_9694;
  wire [13:0] _GEN_9696 = 14'h25e0 == index ? 14'h4b : _GEN_9695;
  wire [13:0] _GEN_9697 = 14'h25e1 == index ? 14'h4b : _GEN_9696;
  wire [13:0] _GEN_9698 = 14'h25e2 == index ? 14'h4b : _GEN_9697;
  wire [13:0] _GEN_9699 = 14'h25e3 == index ? 14'h4b : _GEN_9698;
  wire [13:0] _GEN_9700 = 14'h25e4 == index ? 14'h4b : _GEN_9699;
  wire [13:0] _GEN_9701 = 14'h25e5 == index ? 14'h4b : _GEN_9700;
  wire [13:0] _GEN_9702 = 14'h25e6 == index ? 14'h4b : _GEN_9701;
  wire [13:0] _GEN_9703 = 14'h25e7 == index ? 14'h4b : _GEN_9702;
  wire [13:0] _GEN_9704 = 14'h25e8 == index ? 14'h4b : _GEN_9703;
  wire [13:0] _GEN_9705 = 14'h25e9 == index ? 14'h4b : _GEN_9704;
  wire [13:0] _GEN_9706 = 14'h25ea == index ? 14'h4b : _GEN_9705;
  wire [13:0] _GEN_9707 = 14'h25eb == index ? 14'h4b : _GEN_9706;
  wire [13:0] _GEN_9708 = 14'h25ec == index ? 14'h4b : _GEN_9707;
  wire [13:0] _GEN_9709 = 14'h25ed == index ? 14'h4b : _GEN_9708;
  wire [13:0] _GEN_9710 = 14'h25ee == index ? 14'h4b : _GEN_9709;
  wire [13:0] _GEN_9711 = 14'h25ef == index ? 14'h4b : _GEN_9710;
  wire [13:0] _GEN_9712 = 14'h25f0 == index ? 14'h4b : _GEN_9711;
  wire [13:0] _GEN_9713 = 14'h25f1 == index ? 14'h4b : _GEN_9712;
  wire [13:0] _GEN_9714 = 14'h25f2 == index ? 14'h4b : _GEN_9713;
  wire [13:0] _GEN_9715 = 14'h25f3 == index ? 14'h4b : _GEN_9714;
  wire [13:0] _GEN_9716 = 14'h25f4 == index ? 14'h4b : _GEN_9715;
  wire [13:0] _GEN_9717 = 14'h25f5 == index ? 14'h4b : _GEN_9716;
  wire [13:0] _GEN_9718 = 14'h25f6 == index ? 14'h4b : _GEN_9717;
  wire [13:0] _GEN_9719 = 14'h25f7 == index ? 14'h4b : _GEN_9718;
  wire [13:0] _GEN_9720 = 14'h25f8 == index ? 14'h4b : _GEN_9719;
  wire [13:0] _GEN_9721 = 14'h25f9 == index ? 14'h4b : _GEN_9720;
  wire [13:0] _GEN_9722 = 14'h25fa == index ? 14'h4b : _GEN_9721;
  wire [13:0] _GEN_9723 = 14'h25fb == index ? 14'h4b : _GEN_9722;
  wire [13:0] _GEN_9724 = 14'h25fc == index ? 14'h4b : _GEN_9723;
  wire [13:0] _GEN_9725 = 14'h25fd == index ? 14'h4b : _GEN_9724;
  wire [13:0] _GEN_9726 = 14'h25fe == index ? 14'h4b : _GEN_9725;
  wire [13:0] _GEN_9727 = 14'h25ff == index ? 14'h4b : _GEN_9726;
  wire [13:0] _GEN_9728 = 14'h2600 == index ? 14'h0 : _GEN_9727;
  wire [13:0] _GEN_9729 = 14'h2601 == index ? 14'h2600 : _GEN_9728;
  wire [13:0] _GEN_9730 = 14'h2602 == index ? 14'h1300 : _GEN_9729;
  wire [13:0] _GEN_9731 = 14'h2603 == index ? 14'hc81 : _GEN_9730;
  wire [13:0] _GEN_9732 = 14'h2604 == index ? 14'h980 : _GEN_9731;
  wire [13:0] _GEN_9733 = 14'h2605 == index ? 14'h781 : _GEN_9732;
  wire [13:0] _GEN_9734 = 14'h2606 == index ? 14'h604 : _GEN_9733;
  wire [13:0] _GEN_9735 = 14'h2607 == index ? 14'h506 : _GEN_9734;
  wire [13:0] _GEN_9736 = 14'h2608 == index ? 14'h484 : _GEN_9735;
  wire [13:0] _GEN_9737 = 14'h2609 == index ? 14'h404 : _GEN_9736;
  wire [13:0] _GEN_9738 = 14'h260a == index ? 14'h386 : _GEN_9737;
  wire [13:0] _GEN_9739 = 14'h260b == index ? 14'h30a : _GEN_9738;
  wire [13:0] _GEN_9740 = 14'h260c == index ? 14'h304 : _GEN_9739;
  wire [13:0] _GEN_9741 = 14'h260d == index ? 14'h28b : _GEN_9740;
  wire [13:0] _GEN_9742 = 14'h260e == index ? 14'h286 : _GEN_9741;
  wire [13:0] _GEN_9743 = 14'h260f == index ? 14'h281 : _GEN_9742;
  wire [13:0] _GEN_9744 = 14'h2610 == index ? 14'h20c : _GEN_9743;
  wire [13:0] _GEN_9745 = 14'h2611 == index ? 14'h208 : _GEN_9744;
  wire [13:0] _GEN_9746 = 14'h2612 == index ? 14'h204 : _GEN_9745;
  wire [13:0] _GEN_9747 = 14'h2613 == index ? 14'h200 : _GEN_9746;
  wire [13:0] _GEN_9748 = 14'h2614 == index ? 14'h190 : _GEN_9747;
  wire [13:0] _GEN_9749 = 14'h2615 == index ? 14'h18d : _GEN_9748;
  wire [13:0] _GEN_9750 = 14'h2616 == index ? 14'h18a : _GEN_9749;
  wire [13:0] _GEN_9751 = 14'h2617 == index ? 14'h187 : _GEN_9750;
  wire [13:0] _GEN_9752 = 14'h2618 == index ? 14'h184 : _GEN_9751;
  wire [13:0] _GEN_9753 = 14'h2619 == index ? 14'h181 : _GEN_9752;
  wire [13:0] _GEN_9754 = 14'h261a == index ? 14'h118 : _GEN_9753;
  wire [13:0] _GEN_9755 = 14'h261b == index ? 14'h116 : _GEN_9754;
  wire [13:0] _GEN_9756 = 14'h261c == index ? 14'h114 : _GEN_9755;
  wire [13:0] _GEN_9757 = 14'h261d == index ? 14'h112 : _GEN_9756;
  wire [13:0] _GEN_9758 = 14'h261e == index ? 14'h110 : _GEN_9757;
  wire [13:0] _GEN_9759 = 14'h261f == index ? 14'h10e : _GEN_9758;
  wire [13:0] _GEN_9760 = 14'h2620 == index ? 14'h10c : _GEN_9759;
  wire [13:0] _GEN_9761 = 14'h2621 == index ? 14'h10a : _GEN_9760;
  wire [13:0] _GEN_9762 = 14'h2622 == index ? 14'h108 : _GEN_9761;
  wire [13:0] _GEN_9763 = 14'h2623 == index ? 14'h106 : _GEN_9762;
  wire [13:0] _GEN_9764 = 14'h2624 == index ? 14'h104 : _GEN_9763;
  wire [13:0] _GEN_9765 = 14'h2625 == index ? 14'h102 : _GEN_9764;
  wire [13:0] _GEN_9766 = 14'h2626 == index ? 14'h100 : _GEN_9765;
  wire [13:0] _GEN_9767 = 14'h2627 == index ? 14'ha5 : _GEN_9766;
  wire [13:0] _GEN_9768 = 14'h2628 == index ? 14'ha4 : _GEN_9767;
  wire [13:0] _GEN_9769 = 14'h2629 == index ? 14'ha3 : _GEN_9768;
  wire [13:0] _GEN_9770 = 14'h262a == index ? 14'ha2 : _GEN_9769;
  wire [13:0] _GEN_9771 = 14'h262b == index ? 14'ha1 : _GEN_9770;
  wire [13:0] _GEN_9772 = 14'h262c == index ? 14'ha0 : _GEN_9771;
  wire [13:0] _GEN_9773 = 14'h262d == index ? 14'h9f : _GEN_9772;
  wire [13:0] _GEN_9774 = 14'h262e == index ? 14'h9e : _GEN_9773;
  wire [13:0] _GEN_9775 = 14'h262f == index ? 14'h9d : _GEN_9774;
  wire [13:0] _GEN_9776 = 14'h2630 == index ? 14'h9c : _GEN_9775;
  wire [13:0] _GEN_9777 = 14'h2631 == index ? 14'h9b : _GEN_9776;
  wire [13:0] _GEN_9778 = 14'h2632 == index ? 14'h9a : _GEN_9777;
  wire [13:0] _GEN_9779 = 14'h2633 == index ? 14'h99 : _GEN_9778;
  wire [13:0] _GEN_9780 = 14'h2634 == index ? 14'h98 : _GEN_9779;
  wire [13:0] _GEN_9781 = 14'h2635 == index ? 14'h97 : _GEN_9780;
  wire [13:0] _GEN_9782 = 14'h2636 == index ? 14'h96 : _GEN_9781;
  wire [13:0] _GEN_9783 = 14'h2637 == index ? 14'h95 : _GEN_9782;
  wire [13:0] _GEN_9784 = 14'h2638 == index ? 14'h94 : _GEN_9783;
  wire [13:0] _GEN_9785 = 14'h2639 == index ? 14'h93 : _GEN_9784;
  wire [13:0] _GEN_9786 = 14'h263a == index ? 14'h92 : _GEN_9785;
  wire [13:0] _GEN_9787 = 14'h263b == index ? 14'h91 : _GEN_9786;
  wire [13:0] _GEN_9788 = 14'h263c == index ? 14'h90 : _GEN_9787;
  wire [13:0] _GEN_9789 = 14'h263d == index ? 14'h8f : _GEN_9788;
  wire [13:0] _GEN_9790 = 14'h263e == index ? 14'h8e : _GEN_9789;
  wire [13:0] _GEN_9791 = 14'h263f == index ? 14'h8d : _GEN_9790;
  wire [13:0] _GEN_9792 = 14'h2640 == index ? 14'h8c : _GEN_9791;
  wire [13:0] _GEN_9793 = 14'h2641 == index ? 14'h8b : _GEN_9792;
  wire [13:0] _GEN_9794 = 14'h2642 == index ? 14'h8a : _GEN_9793;
  wire [13:0] _GEN_9795 = 14'h2643 == index ? 14'h89 : _GEN_9794;
  wire [13:0] _GEN_9796 = 14'h2644 == index ? 14'h88 : _GEN_9795;
  wire [13:0] _GEN_9797 = 14'h2645 == index ? 14'h87 : _GEN_9796;
  wire [13:0] _GEN_9798 = 14'h2646 == index ? 14'h86 : _GEN_9797;
  wire [13:0] _GEN_9799 = 14'h2647 == index ? 14'h85 : _GEN_9798;
  wire [13:0] _GEN_9800 = 14'h2648 == index ? 14'h84 : _GEN_9799;
  wire [13:0] _GEN_9801 = 14'h2649 == index ? 14'h83 : _GEN_9800;
  wire [13:0] _GEN_9802 = 14'h264a == index ? 14'h82 : _GEN_9801;
  wire [13:0] _GEN_9803 = 14'h264b == index ? 14'h81 : _GEN_9802;
  wire [13:0] _GEN_9804 = 14'h264c == index ? 14'h80 : _GEN_9803;
  wire [13:0] _GEN_9805 = 14'h264d == index ? 14'h4c : _GEN_9804;
  wire [13:0] _GEN_9806 = 14'h264e == index ? 14'h4c : _GEN_9805;
  wire [13:0] _GEN_9807 = 14'h264f == index ? 14'h4c : _GEN_9806;
  wire [13:0] _GEN_9808 = 14'h2650 == index ? 14'h4c : _GEN_9807;
  wire [13:0] _GEN_9809 = 14'h2651 == index ? 14'h4c : _GEN_9808;
  wire [13:0] _GEN_9810 = 14'h2652 == index ? 14'h4c : _GEN_9809;
  wire [13:0] _GEN_9811 = 14'h2653 == index ? 14'h4c : _GEN_9810;
  wire [13:0] _GEN_9812 = 14'h2654 == index ? 14'h4c : _GEN_9811;
  wire [13:0] _GEN_9813 = 14'h2655 == index ? 14'h4c : _GEN_9812;
  wire [13:0] _GEN_9814 = 14'h2656 == index ? 14'h4c : _GEN_9813;
  wire [13:0] _GEN_9815 = 14'h2657 == index ? 14'h4c : _GEN_9814;
  wire [13:0] _GEN_9816 = 14'h2658 == index ? 14'h4c : _GEN_9815;
  wire [13:0] _GEN_9817 = 14'h2659 == index ? 14'h4c : _GEN_9816;
  wire [13:0] _GEN_9818 = 14'h265a == index ? 14'h4c : _GEN_9817;
  wire [13:0] _GEN_9819 = 14'h265b == index ? 14'h4c : _GEN_9818;
  wire [13:0] _GEN_9820 = 14'h265c == index ? 14'h4c : _GEN_9819;
  wire [13:0] _GEN_9821 = 14'h265d == index ? 14'h4c : _GEN_9820;
  wire [13:0] _GEN_9822 = 14'h265e == index ? 14'h4c : _GEN_9821;
  wire [13:0] _GEN_9823 = 14'h265f == index ? 14'h4c : _GEN_9822;
  wire [13:0] _GEN_9824 = 14'h2660 == index ? 14'h4c : _GEN_9823;
  wire [13:0] _GEN_9825 = 14'h2661 == index ? 14'h4c : _GEN_9824;
  wire [13:0] _GEN_9826 = 14'h2662 == index ? 14'h4c : _GEN_9825;
  wire [13:0] _GEN_9827 = 14'h2663 == index ? 14'h4c : _GEN_9826;
  wire [13:0] _GEN_9828 = 14'h2664 == index ? 14'h4c : _GEN_9827;
  wire [13:0] _GEN_9829 = 14'h2665 == index ? 14'h4c : _GEN_9828;
  wire [13:0] _GEN_9830 = 14'h2666 == index ? 14'h4c : _GEN_9829;
  wire [13:0] _GEN_9831 = 14'h2667 == index ? 14'h4c : _GEN_9830;
  wire [13:0] _GEN_9832 = 14'h2668 == index ? 14'h4c : _GEN_9831;
  wire [13:0] _GEN_9833 = 14'h2669 == index ? 14'h4c : _GEN_9832;
  wire [13:0] _GEN_9834 = 14'h266a == index ? 14'h4c : _GEN_9833;
  wire [13:0] _GEN_9835 = 14'h266b == index ? 14'h4c : _GEN_9834;
  wire [13:0] _GEN_9836 = 14'h266c == index ? 14'h4c : _GEN_9835;
  wire [13:0] _GEN_9837 = 14'h266d == index ? 14'h4c : _GEN_9836;
  wire [13:0] _GEN_9838 = 14'h266e == index ? 14'h4c : _GEN_9837;
  wire [13:0] _GEN_9839 = 14'h266f == index ? 14'h4c : _GEN_9838;
  wire [13:0] _GEN_9840 = 14'h2670 == index ? 14'h4c : _GEN_9839;
  wire [13:0] _GEN_9841 = 14'h2671 == index ? 14'h4c : _GEN_9840;
  wire [13:0] _GEN_9842 = 14'h2672 == index ? 14'h4c : _GEN_9841;
  wire [13:0] _GEN_9843 = 14'h2673 == index ? 14'h4c : _GEN_9842;
  wire [13:0] _GEN_9844 = 14'h2674 == index ? 14'h4c : _GEN_9843;
  wire [13:0] _GEN_9845 = 14'h2675 == index ? 14'h4c : _GEN_9844;
  wire [13:0] _GEN_9846 = 14'h2676 == index ? 14'h4c : _GEN_9845;
  wire [13:0] _GEN_9847 = 14'h2677 == index ? 14'h4c : _GEN_9846;
  wire [13:0] _GEN_9848 = 14'h2678 == index ? 14'h4c : _GEN_9847;
  wire [13:0] _GEN_9849 = 14'h2679 == index ? 14'h4c : _GEN_9848;
  wire [13:0] _GEN_9850 = 14'h267a == index ? 14'h4c : _GEN_9849;
  wire [13:0] _GEN_9851 = 14'h267b == index ? 14'h4c : _GEN_9850;
  wire [13:0] _GEN_9852 = 14'h267c == index ? 14'h4c : _GEN_9851;
  wire [13:0] _GEN_9853 = 14'h267d == index ? 14'h4c : _GEN_9852;
  wire [13:0] _GEN_9854 = 14'h267e == index ? 14'h4c : _GEN_9853;
  wire [13:0] _GEN_9855 = 14'h267f == index ? 14'h4c : _GEN_9854;
  wire [13:0] _GEN_9856 = 14'h2680 == index ? 14'h0 : _GEN_9855;
  wire [13:0] _GEN_9857 = 14'h2681 == index ? 14'h2680 : _GEN_9856;
  wire [13:0] _GEN_9858 = 14'h2682 == index ? 14'h1301 : _GEN_9857;
  wire [13:0] _GEN_9859 = 14'h2683 == index ? 14'hc82 : _GEN_9858;
  wire [13:0] _GEN_9860 = 14'h2684 == index ? 14'h981 : _GEN_9859;
  wire [13:0] _GEN_9861 = 14'h2685 == index ? 14'h782 : _GEN_9860;
  wire [13:0] _GEN_9862 = 14'h2686 == index ? 14'h605 : _GEN_9861;
  wire [13:0] _GEN_9863 = 14'h2687 == index ? 14'h580 : _GEN_9862;
  wire [13:0] _GEN_9864 = 14'h2688 == index ? 14'h485 : _GEN_9863;
  wire [13:0] _GEN_9865 = 14'h2689 == index ? 14'h405 : _GEN_9864;
  wire [13:0] _GEN_9866 = 14'h268a == index ? 14'h387 : _GEN_9865;
  wire [13:0] _GEN_9867 = 14'h268b == index ? 14'h380 : _GEN_9866;
  wire [13:0] _GEN_9868 = 14'h268c == index ? 14'h305 : _GEN_9867;
  wire [13:0] _GEN_9869 = 14'h268d == index ? 14'h28c : _GEN_9868;
  wire [13:0] _GEN_9870 = 14'h268e == index ? 14'h287 : _GEN_9869;
  wire [13:0] _GEN_9871 = 14'h268f == index ? 14'h282 : _GEN_9870;
  wire [13:0] _GEN_9872 = 14'h2690 == index ? 14'h20d : _GEN_9871;
  wire [13:0] _GEN_9873 = 14'h2691 == index ? 14'h209 : _GEN_9872;
  wire [13:0] _GEN_9874 = 14'h2692 == index ? 14'h205 : _GEN_9873;
  wire [13:0] _GEN_9875 = 14'h2693 == index ? 14'h201 : _GEN_9874;
  wire [13:0] _GEN_9876 = 14'h2694 == index ? 14'h191 : _GEN_9875;
  wire [13:0] _GEN_9877 = 14'h2695 == index ? 14'h18e : _GEN_9876;
  wire [13:0] _GEN_9878 = 14'h2696 == index ? 14'h18b : _GEN_9877;
  wire [13:0] _GEN_9879 = 14'h2697 == index ? 14'h188 : _GEN_9878;
  wire [13:0] _GEN_9880 = 14'h2698 == index ? 14'h185 : _GEN_9879;
  wire [13:0] _GEN_9881 = 14'h2699 == index ? 14'h182 : _GEN_9880;
  wire [13:0] _GEN_9882 = 14'h269a == index ? 14'h119 : _GEN_9881;
  wire [13:0] _GEN_9883 = 14'h269b == index ? 14'h117 : _GEN_9882;
  wire [13:0] _GEN_9884 = 14'h269c == index ? 14'h115 : _GEN_9883;
  wire [13:0] _GEN_9885 = 14'h269d == index ? 14'h113 : _GEN_9884;
  wire [13:0] _GEN_9886 = 14'h269e == index ? 14'h111 : _GEN_9885;
  wire [13:0] _GEN_9887 = 14'h269f == index ? 14'h10f : _GEN_9886;
  wire [13:0] _GEN_9888 = 14'h26a0 == index ? 14'h10d : _GEN_9887;
  wire [13:0] _GEN_9889 = 14'h26a1 == index ? 14'h10b : _GEN_9888;
  wire [13:0] _GEN_9890 = 14'h26a2 == index ? 14'h109 : _GEN_9889;
  wire [13:0] _GEN_9891 = 14'h26a3 == index ? 14'h107 : _GEN_9890;
  wire [13:0] _GEN_9892 = 14'h26a4 == index ? 14'h105 : _GEN_9891;
  wire [13:0] _GEN_9893 = 14'h26a5 == index ? 14'h103 : _GEN_9892;
  wire [13:0] _GEN_9894 = 14'h26a6 == index ? 14'h101 : _GEN_9893;
  wire [13:0] _GEN_9895 = 14'h26a7 == index ? 14'ha6 : _GEN_9894;
  wire [13:0] _GEN_9896 = 14'h26a8 == index ? 14'ha5 : _GEN_9895;
  wire [13:0] _GEN_9897 = 14'h26a9 == index ? 14'ha4 : _GEN_9896;
  wire [13:0] _GEN_9898 = 14'h26aa == index ? 14'ha3 : _GEN_9897;
  wire [13:0] _GEN_9899 = 14'h26ab == index ? 14'ha2 : _GEN_9898;
  wire [13:0] _GEN_9900 = 14'h26ac == index ? 14'ha1 : _GEN_9899;
  wire [13:0] _GEN_9901 = 14'h26ad == index ? 14'ha0 : _GEN_9900;
  wire [13:0] _GEN_9902 = 14'h26ae == index ? 14'h9f : _GEN_9901;
  wire [13:0] _GEN_9903 = 14'h26af == index ? 14'h9e : _GEN_9902;
  wire [13:0] _GEN_9904 = 14'h26b0 == index ? 14'h9d : _GEN_9903;
  wire [13:0] _GEN_9905 = 14'h26b1 == index ? 14'h9c : _GEN_9904;
  wire [13:0] _GEN_9906 = 14'h26b2 == index ? 14'h9b : _GEN_9905;
  wire [13:0] _GEN_9907 = 14'h26b3 == index ? 14'h9a : _GEN_9906;
  wire [13:0] _GEN_9908 = 14'h26b4 == index ? 14'h99 : _GEN_9907;
  wire [13:0] _GEN_9909 = 14'h26b5 == index ? 14'h98 : _GEN_9908;
  wire [13:0] _GEN_9910 = 14'h26b6 == index ? 14'h97 : _GEN_9909;
  wire [13:0] _GEN_9911 = 14'h26b7 == index ? 14'h96 : _GEN_9910;
  wire [13:0] _GEN_9912 = 14'h26b8 == index ? 14'h95 : _GEN_9911;
  wire [13:0] _GEN_9913 = 14'h26b9 == index ? 14'h94 : _GEN_9912;
  wire [13:0] _GEN_9914 = 14'h26ba == index ? 14'h93 : _GEN_9913;
  wire [13:0] _GEN_9915 = 14'h26bb == index ? 14'h92 : _GEN_9914;
  wire [13:0] _GEN_9916 = 14'h26bc == index ? 14'h91 : _GEN_9915;
  wire [13:0] _GEN_9917 = 14'h26bd == index ? 14'h90 : _GEN_9916;
  wire [13:0] _GEN_9918 = 14'h26be == index ? 14'h8f : _GEN_9917;
  wire [13:0] _GEN_9919 = 14'h26bf == index ? 14'h8e : _GEN_9918;
  wire [13:0] _GEN_9920 = 14'h26c0 == index ? 14'h8d : _GEN_9919;
  wire [13:0] _GEN_9921 = 14'h26c1 == index ? 14'h8c : _GEN_9920;
  wire [13:0] _GEN_9922 = 14'h26c2 == index ? 14'h8b : _GEN_9921;
  wire [13:0] _GEN_9923 = 14'h26c3 == index ? 14'h8a : _GEN_9922;
  wire [13:0] _GEN_9924 = 14'h26c4 == index ? 14'h89 : _GEN_9923;
  wire [13:0] _GEN_9925 = 14'h26c5 == index ? 14'h88 : _GEN_9924;
  wire [13:0] _GEN_9926 = 14'h26c6 == index ? 14'h87 : _GEN_9925;
  wire [13:0] _GEN_9927 = 14'h26c7 == index ? 14'h86 : _GEN_9926;
  wire [13:0] _GEN_9928 = 14'h26c8 == index ? 14'h85 : _GEN_9927;
  wire [13:0] _GEN_9929 = 14'h26c9 == index ? 14'h84 : _GEN_9928;
  wire [13:0] _GEN_9930 = 14'h26ca == index ? 14'h83 : _GEN_9929;
  wire [13:0] _GEN_9931 = 14'h26cb == index ? 14'h82 : _GEN_9930;
  wire [13:0] _GEN_9932 = 14'h26cc == index ? 14'h81 : _GEN_9931;
  wire [13:0] _GEN_9933 = 14'h26cd == index ? 14'h80 : _GEN_9932;
  wire [13:0] _GEN_9934 = 14'h26ce == index ? 14'h4d : _GEN_9933;
  wire [13:0] _GEN_9935 = 14'h26cf == index ? 14'h4d : _GEN_9934;
  wire [13:0] _GEN_9936 = 14'h26d0 == index ? 14'h4d : _GEN_9935;
  wire [13:0] _GEN_9937 = 14'h26d1 == index ? 14'h4d : _GEN_9936;
  wire [13:0] _GEN_9938 = 14'h26d2 == index ? 14'h4d : _GEN_9937;
  wire [13:0] _GEN_9939 = 14'h26d3 == index ? 14'h4d : _GEN_9938;
  wire [13:0] _GEN_9940 = 14'h26d4 == index ? 14'h4d : _GEN_9939;
  wire [13:0] _GEN_9941 = 14'h26d5 == index ? 14'h4d : _GEN_9940;
  wire [13:0] _GEN_9942 = 14'h26d6 == index ? 14'h4d : _GEN_9941;
  wire [13:0] _GEN_9943 = 14'h26d7 == index ? 14'h4d : _GEN_9942;
  wire [13:0] _GEN_9944 = 14'h26d8 == index ? 14'h4d : _GEN_9943;
  wire [13:0] _GEN_9945 = 14'h26d9 == index ? 14'h4d : _GEN_9944;
  wire [13:0] _GEN_9946 = 14'h26da == index ? 14'h4d : _GEN_9945;
  wire [13:0] _GEN_9947 = 14'h26db == index ? 14'h4d : _GEN_9946;
  wire [13:0] _GEN_9948 = 14'h26dc == index ? 14'h4d : _GEN_9947;
  wire [13:0] _GEN_9949 = 14'h26dd == index ? 14'h4d : _GEN_9948;
  wire [13:0] _GEN_9950 = 14'h26de == index ? 14'h4d : _GEN_9949;
  wire [13:0] _GEN_9951 = 14'h26df == index ? 14'h4d : _GEN_9950;
  wire [13:0] _GEN_9952 = 14'h26e0 == index ? 14'h4d : _GEN_9951;
  wire [13:0] _GEN_9953 = 14'h26e1 == index ? 14'h4d : _GEN_9952;
  wire [13:0] _GEN_9954 = 14'h26e2 == index ? 14'h4d : _GEN_9953;
  wire [13:0] _GEN_9955 = 14'h26e3 == index ? 14'h4d : _GEN_9954;
  wire [13:0] _GEN_9956 = 14'h26e4 == index ? 14'h4d : _GEN_9955;
  wire [13:0] _GEN_9957 = 14'h26e5 == index ? 14'h4d : _GEN_9956;
  wire [13:0] _GEN_9958 = 14'h26e6 == index ? 14'h4d : _GEN_9957;
  wire [13:0] _GEN_9959 = 14'h26e7 == index ? 14'h4d : _GEN_9958;
  wire [13:0] _GEN_9960 = 14'h26e8 == index ? 14'h4d : _GEN_9959;
  wire [13:0] _GEN_9961 = 14'h26e9 == index ? 14'h4d : _GEN_9960;
  wire [13:0] _GEN_9962 = 14'h26ea == index ? 14'h4d : _GEN_9961;
  wire [13:0] _GEN_9963 = 14'h26eb == index ? 14'h4d : _GEN_9962;
  wire [13:0] _GEN_9964 = 14'h26ec == index ? 14'h4d : _GEN_9963;
  wire [13:0] _GEN_9965 = 14'h26ed == index ? 14'h4d : _GEN_9964;
  wire [13:0] _GEN_9966 = 14'h26ee == index ? 14'h4d : _GEN_9965;
  wire [13:0] _GEN_9967 = 14'h26ef == index ? 14'h4d : _GEN_9966;
  wire [13:0] _GEN_9968 = 14'h26f0 == index ? 14'h4d : _GEN_9967;
  wire [13:0] _GEN_9969 = 14'h26f1 == index ? 14'h4d : _GEN_9968;
  wire [13:0] _GEN_9970 = 14'h26f2 == index ? 14'h4d : _GEN_9969;
  wire [13:0] _GEN_9971 = 14'h26f3 == index ? 14'h4d : _GEN_9970;
  wire [13:0] _GEN_9972 = 14'h26f4 == index ? 14'h4d : _GEN_9971;
  wire [13:0] _GEN_9973 = 14'h26f5 == index ? 14'h4d : _GEN_9972;
  wire [13:0] _GEN_9974 = 14'h26f6 == index ? 14'h4d : _GEN_9973;
  wire [13:0] _GEN_9975 = 14'h26f7 == index ? 14'h4d : _GEN_9974;
  wire [13:0] _GEN_9976 = 14'h26f8 == index ? 14'h4d : _GEN_9975;
  wire [13:0] _GEN_9977 = 14'h26f9 == index ? 14'h4d : _GEN_9976;
  wire [13:0] _GEN_9978 = 14'h26fa == index ? 14'h4d : _GEN_9977;
  wire [13:0] _GEN_9979 = 14'h26fb == index ? 14'h4d : _GEN_9978;
  wire [13:0] _GEN_9980 = 14'h26fc == index ? 14'h4d : _GEN_9979;
  wire [13:0] _GEN_9981 = 14'h26fd == index ? 14'h4d : _GEN_9980;
  wire [13:0] _GEN_9982 = 14'h26fe == index ? 14'h4d : _GEN_9981;
  wire [13:0] _GEN_9983 = 14'h26ff == index ? 14'h4d : _GEN_9982;
  wire [13:0] _GEN_9984 = 14'h2700 == index ? 14'h0 : _GEN_9983;
  wire [13:0] _GEN_9985 = 14'h2701 == index ? 14'h2700 : _GEN_9984;
  wire [13:0] _GEN_9986 = 14'h2702 == index ? 14'h1380 : _GEN_9985;
  wire [13:0] _GEN_9987 = 14'h2703 == index ? 14'hd00 : _GEN_9986;
  wire [13:0] _GEN_9988 = 14'h2704 == index ? 14'h982 : _GEN_9987;
  wire [13:0] _GEN_9989 = 14'h2705 == index ? 14'h783 : _GEN_9988;
  wire [13:0] _GEN_9990 = 14'h2706 == index ? 14'h680 : _GEN_9989;
  wire [13:0] _GEN_9991 = 14'h2707 == index ? 14'h581 : _GEN_9990;
  wire [13:0] _GEN_9992 = 14'h2708 == index ? 14'h486 : _GEN_9991;
  wire [13:0] _GEN_9993 = 14'h2709 == index ? 14'h406 : _GEN_9992;
  wire [13:0] _GEN_9994 = 14'h270a == index ? 14'h388 : _GEN_9993;
  wire [13:0] _GEN_9995 = 14'h270b == index ? 14'h381 : _GEN_9994;
  wire [13:0] _GEN_9996 = 14'h270c == index ? 14'h306 : _GEN_9995;
  wire [13:0] _GEN_9997 = 14'h270d == index ? 14'h300 : _GEN_9996;
  wire [13:0] _GEN_9998 = 14'h270e == index ? 14'h288 : _GEN_9997;
  wire [13:0] _GEN_9999 = 14'h270f == index ? 14'h283 : _GEN_9998;
  wire [13:0] _GEN_10000 = 14'h2710 == index ? 14'h20e : _GEN_9999;
  wire [13:0] _GEN_10001 = 14'h2711 == index ? 14'h20a : _GEN_10000;
  wire [13:0] _GEN_10002 = 14'h2712 == index ? 14'h206 : _GEN_10001;
  wire [13:0] _GEN_10003 = 14'h2713 == index ? 14'h202 : _GEN_10002;
  wire [13:0] _GEN_10004 = 14'h2714 == index ? 14'h192 : _GEN_10003;
  wire [13:0] _GEN_10005 = 14'h2715 == index ? 14'h18f : _GEN_10004;
  wire [13:0] _GEN_10006 = 14'h2716 == index ? 14'h18c : _GEN_10005;
  wire [13:0] _GEN_10007 = 14'h2717 == index ? 14'h189 : _GEN_10006;
  wire [13:0] _GEN_10008 = 14'h2718 == index ? 14'h186 : _GEN_10007;
  wire [13:0] _GEN_10009 = 14'h2719 == index ? 14'h183 : _GEN_10008;
  wire [13:0] _GEN_10010 = 14'h271a == index ? 14'h180 : _GEN_10009;
  wire [13:0] _GEN_10011 = 14'h271b == index ? 14'h118 : _GEN_10010;
  wire [13:0] _GEN_10012 = 14'h271c == index ? 14'h116 : _GEN_10011;
  wire [13:0] _GEN_10013 = 14'h271d == index ? 14'h114 : _GEN_10012;
  wire [13:0] _GEN_10014 = 14'h271e == index ? 14'h112 : _GEN_10013;
  wire [13:0] _GEN_10015 = 14'h271f == index ? 14'h110 : _GEN_10014;
  wire [13:0] _GEN_10016 = 14'h2720 == index ? 14'h10e : _GEN_10015;
  wire [13:0] _GEN_10017 = 14'h2721 == index ? 14'h10c : _GEN_10016;
  wire [13:0] _GEN_10018 = 14'h2722 == index ? 14'h10a : _GEN_10017;
  wire [13:0] _GEN_10019 = 14'h2723 == index ? 14'h108 : _GEN_10018;
  wire [13:0] _GEN_10020 = 14'h2724 == index ? 14'h106 : _GEN_10019;
  wire [13:0] _GEN_10021 = 14'h2725 == index ? 14'h104 : _GEN_10020;
  wire [13:0] _GEN_10022 = 14'h2726 == index ? 14'h102 : _GEN_10021;
  wire [13:0] _GEN_10023 = 14'h2727 == index ? 14'h100 : _GEN_10022;
  wire [13:0] _GEN_10024 = 14'h2728 == index ? 14'ha6 : _GEN_10023;
  wire [13:0] _GEN_10025 = 14'h2729 == index ? 14'ha5 : _GEN_10024;
  wire [13:0] _GEN_10026 = 14'h272a == index ? 14'ha4 : _GEN_10025;
  wire [13:0] _GEN_10027 = 14'h272b == index ? 14'ha3 : _GEN_10026;
  wire [13:0] _GEN_10028 = 14'h272c == index ? 14'ha2 : _GEN_10027;
  wire [13:0] _GEN_10029 = 14'h272d == index ? 14'ha1 : _GEN_10028;
  wire [13:0] _GEN_10030 = 14'h272e == index ? 14'ha0 : _GEN_10029;
  wire [13:0] _GEN_10031 = 14'h272f == index ? 14'h9f : _GEN_10030;
  wire [13:0] _GEN_10032 = 14'h2730 == index ? 14'h9e : _GEN_10031;
  wire [13:0] _GEN_10033 = 14'h2731 == index ? 14'h9d : _GEN_10032;
  wire [13:0] _GEN_10034 = 14'h2732 == index ? 14'h9c : _GEN_10033;
  wire [13:0] _GEN_10035 = 14'h2733 == index ? 14'h9b : _GEN_10034;
  wire [13:0] _GEN_10036 = 14'h2734 == index ? 14'h9a : _GEN_10035;
  wire [13:0] _GEN_10037 = 14'h2735 == index ? 14'h99 : _GEN_10036;
  wire [13:0] _GEN_10038 = 14'h2736 == index ? 14'h98 : _GEN_10037;
  wire [13:0] _GEN_10039 = 14'h2737 == index ? 14'h97 : _GEN_10038;
  wire [13:0] _GEN_10040 = 14'h2738 == index ? 14'h96 : _GEN_10039;
  wire [13:0] _GEN_10041 = 14'h2739 == index ? 14'h95 : _GEN_10040;
  wire [13:0] _GEN_10042 = 14'h273a == index ? 14'h94 : _GEN_10041;
  wire [13:0] _GEN_10043 = 14'h273b == index ? 14'h93 : _GEN_10042;
  wire [13:0] _GEN_10044 = 14'h273c == index ? 14'h92 : _GEN_10043;
  wire [13:0] _GEN_10045 = 14'h273d == index ? 14'h91 : _GEN_10044;
  wire [13:0] _GEN_10046 = 14'h273e == index ? 14'h90 : _GEN_10045;
  wire [13:0] _GEN_10047 = 14'h273f == index ? 14'h8f : _GEN_10046;
  wire [13:0] _GEN_10048 = 14'h2740 == index ? 14'h8e : _GEN_10047;
  wire [13:0] _GEN_10049 = 14'h2741 == index ? 14'h8d : _GEN_10048;
  wire [13:0] _GEN_10050 = 14'h2742 == index ? 14'h8c : _GEN_10049;
  wire [13:0] _GEN_10051 = 14'h2743 == index ? 14'h8b : _GEN_10050;
  wire [13:0] _GEN_10052 = 14'h2744 == index ? 14'h8a : _GEN_10051;
  wire [13:0] _GEN_10053 = 14'h2745 == index ? 14'h89 : _GEN_10052;
  wire [13:0] _GEN_10054 = 14'h2746 == index ? 14'h88 : _GEN_10053;
  wire [13:0] _GEN_10055 = 14'h2747 == index ? 14'h87 : _GEN_10054;
  wire [13:0] _GEN_10056 = 14'h2748 == index ? 14'h86 : _GEN_10055;
  wire [13:0] _GEN_10057 = 14'h2749 == index ? 14'h85 : _GEN_10056;
  wire [13:0] _GEN_10058 = 14'h274a == index ? 14'h84 : _GEN_10057;
  wire [13:0] _GEN_10059 = 14'h274b == index ? 14'h83 : _GEN_10058;
  wire [13:0] _GEN_10060 = 14'h274c == index ? 14'h82 : _GEN_10059;
  wire [13:0] _GEN_10061 = 14'h274d == index ? 14'h81 : _GEN_10060;
  wire [13:0] _GEN_10062 = 14'h274e == index ? 14'h80 : _GEN_10061;
  wire [13:0] _GEN_10063 = 14'h274f == index ? 14'h4e : _GEN_10062;
  wire [13:0] _GEN_10064 = 14'h2750 == index ? 14'h4e : _GEN_10063;
  wire [13:0] _GEN_10065 = 14'h2751 == index ? 14'h4e : _GEN_10064;
  wire [13:0] _GEN_10066 = 14'h2752 == index ? 14'h4e : _GEN_10065;
  wire [13:0] _GEN_10067 = 14'h2753 == index ? 14'h4e : _GEN_10066;
  wire [13:0] _GEN_10068 = 14'h2754 == index ? 14'h4e : _GEN_10067;
  wire [13:0] _GEN_10069 = 14'h2755 == index ? 14'h4e : _GEN_10068;
  wire [13:0] _GEN_10070 = 14'h2756 == index ? 14'h4e : _GEN_10069;
  wire [13:0] _GEN_10071 = 14'h2757 == index ? 14'h4e : _GEN_10070;
  wire [13:0] _GEN_10072 = 14'h2758 == index ? 14'h4e : _GEN_10071;
  wire [13:0] _GEN_10073 = 14'h2759 == index ? 14'h4e : _GEN_10072;
  wire [13:0] _GEN_10074 = 14'h275a == index ? 14'h4e : _GEN_10073;
  wire [13:0] _GEN_10075 = 14'h275b == index ? 14'h4e : _GEN_10074;
  wire [13:0] _GEN_10076 = 14'h275c == index ? 14'h4e : _GEN_10075;
  wire [13:0] _GEN_10077 = 14'h275d == index ? 14'h4e : _GEN_10076;
  wire [13:0] _GEN_10078 = 14'h275e == index ? 14'h4e : _GEN_10077;
  wire [13:0] _GEN_10079 = 14'h275f == index ? 14'h4e : _GEN_10078;
  wire [13:0] _GEN_10080 = 14'h2760 == index ? 14'h4e : _GEN_10079;
  wire [13:0] _GEN_10081 = 14'h2761 == index ? 14'h4e : _GEN_10080;
  wire [13:0] _GEN_10082 = 14'h2762 == index ? 14'h4e : _GEN_10081;
  wire [13:0] _GEN_10083 = 14'h2763 == index ? 14'h4e : _GEN_10082;
  wire [13:0] _GEN_10084 = 14'h2764 == index ? 14'h4e : _GEN_10083;
  wire [13:0] _GEN_10085 = 14'h2765 == index ? 14'h4e : _GEN_10084;
  wire [13:0] _GEN_10086 = 14'h2766 == index ? 14'h4e : _GEN_10085;
  wire [13:0] _GEN_10087 = 14'h2767 == index ? 14'h4e : _GEN_10086;
  wire [13:0] _GEN_10088 = 14'h2768 == index ? 14'h4e : _GEN_10087;
  wire [13:0] _GEN_10089 = 14'h2769 == index ? 14'h4e : _GEN_10088;
  wire [13:0] _GEN_10090 = 14'h276a == index ? 14'h4e : _GEN_10089;
  wire [13:0] _GEN_10091 = 14'h276b == index ? 14'h4e : _GEN_10090;
  wire [13:0] _GEN_10092 = 14'h276c == index ? 14'h4e : _GEN_10091;
  wire [13:0] _GEN_10093 = 14'h276d == index ? 14'h4e : _GEN_10092;
  wire [13:0] _GEN_10094 = 14'h276e == index ? 14'h4e : _GEN_10093;
  wire [13:0] _GEN_10095 = 14'h276f == index ? 14'h4e : _GEN_10094;
  wire [13:0] _GEN_10096 = 14'h2770 == index ? 14'h4e : _GEN_10095;
  wire [13:0] _GEN_10097 = 14'h2771 == index ? 14'h4e : _GEN_10096;
  wire [13:0] _GEN_10098 = 14'h2772 == index ? 14'h4e : _GEN_10097;
  wire [13:0] _GEN_10099 = 14'h2773 == index ? 14'h4e : _GEN_10098;
  wire [13:0] _GEN_10100 = 14'h2774 == index ? 14'h4e : _GEN_10099;
  wire [13:0] _GEN_10101 = 14'h2775 == index ? 14'h4e : _GEN_10100;
  wire [13:0] _GEN_10102 = 14'h2776 == index ? 14'h4e : _GEN_10101;
  wire [13:0] _GEN_10103 = 14'h2777 == index ? 14'h4e : _GEN_10102;
  wire [13:0] _GEN_10104 = 14'h2778 == index ? 14'h4e : _GEN_10103;
  wire [13:0] _GEN_10105 = 14'h2779 == index ? 14'h4e : _GEN_10104;
  wire [13:0] _GEN_10106 = 14'h277a == index ? 14'h4e : _GEN_10105;
  wire [13:0] _GEN_10107 = 14'h277b == index ? 14'h4e : _GEN_10106;
  wire [13:0] _GEN_10108 = 14'h277c == index ? 14'h4e : _GEN_10107;
  wire [13:0] _GEN_10109 = 14'h277d == index ? 14'h4e : _GEN_10108;
  wire [13:0] _GEN_10110 = 14'h277e == index ? 14'h4e : _GEN_10109;
  wire [13:0] _GEN_10111 = 14'h277f == index ? 14'h4e : _GEN_10110;
  wire [13:0] _GEN_10112 = 14'h2780 == index ? 14'h0 : _GEN_10111;
  wire [13:0] _GEN_10113 = 14'h2781 == index ? 14'h2780 : _GEN_10112;
  wire [13:0] _GEN_10114 = 14'h2782 == index ? 14'h1381 : _GEN_10113;
  wire [13:0] _GEN_10115 = 14'h2783 == index ? 14'hd01 : _GEN_10114;
  wire [13:0] _GEN_10116 = 14'h2784 == index ? 14'h983 : _GEN_10115;
  wire [13:0] _GEN_10117 = 14'h2785 == index ? 14'h784 : _GEN_10116;
  wire [13:0] _GEN_10118 = 14'h2786 == index ? 14'h681 : _GEN_10117;
  wire [13:0] _GEN_10119 = 14'h2787 == index ? 14'h582 : _GEN_10118;
  wire [13:0] _GEN_10120 = 14'h2788 == index ? 14'h487 : _GEN_10119;
  wire [13:0] _GEN_10121 = 14'h2789 == index ? 14'h407 : _GEN_10120;
  wire [13:0] _GEN_10122 = 14'h278a == index ? 14'h389 : _GEN_10121;
  wire [13:0] _GEN_10123 = 14'h278b == index ? 14'h382 : _GEN_10122;
  wire [13:0] _GEN_10124 = 14'h278c == index ? 14'h307 : _GEN_10123;
  wire [13:0] _GEN_10125 = 14'h278d == index ? 14'h301 : _GEN_10124;
  wire [13:0] _GEN_10126 = 14'h278e == index ? 14'h289 : _GEN_10125;
  wire [13:0] _GEN_10127 = 14'h278f == index ? 14'h284 : _GEN_10126;
  wire [13:0] _GEN_10128 = 14'h2790 == index ? 14'h20f : _GEN_10127;
  wire [13:0] _GEN_10129 = 14'h2791 == index ? 14'h20b : _GEN_10128;
  wire [13:0] _GEN_10130 = 14'h2792 == index ? 14'h207 : _GEN_10129;
  wire [13:0] _GEN_10131 = 14'h2793 == index ? 14'h203 : _GEN_10130;
  wire [13:0] _GEN_10132 = 14'h2794 == index ? 14'h193 : _GEN_10131;
  wire [13:0] _GEN_10133 = 14'h2795 == index ? 14'h190 : _GEN_10132;
  wire [13:0] _GEN_10134 = 14'h2796 == index ? 14'h18d : _GEN_10133;
  wire [13:0] _GEN_10135 = 14'h2797 == index ? 14'h18a : _GEN_10134;
  wire [13:0] _GEN_10136 = 14'h2798 == index ? 14'h187 : _GEN_10135;
  wire [13:0] _GEN_10137 = 14'h2799 == index ? 14'h184 : _GEN_10136;
  wire [13:0] _GEN_10138 = 14'h279a == index ? 14'h181 : _GEN_10137;
  wire [13:0] _GEN_10139 = 14'h279b == index ? 14'h119 : _GEN_10138;
  wire [13:0] _GEN_10140 = 14'h279c == index ? 14'h117 : _GEN_10139;
  wire [13:0] _GEN_10141 = 14'h279d == index ? 14'h115 : _GEN_10140;
  wire [13:0] _GEN_10142 = 14'h279e == index ? 14'h113 : _GEN_10141;
  wire [13:0] _GEN_10143 = 14'h279f == index ? 14'h111 : _GEN_10142;
  wire [13:0] _GEN_10144 = 14'h27a0 == index ? 14'h10f : _GEN_10143;
  wire [13:0] _GEN_10145 = 14'h27a1 == index ? 14'h10d : _GEN_10144;
  wire [13:0] _GEN_10146 = 14'h27a2 == index ? 14'h10b : _GEN_10145;
  wire [13:0] _GEN_10147 = 14'h27a3 == index ? 14'h109 : _GEN_10146;
  wire [13:0] _GEN_10148 = 14'h27a4 == index ? 14'h107 : _GEN_10147;
  wire [13:0] _GEN_10149 = 14'h27a5 == index ? 14'h105 : _GEN_10148;
  wire [13:0] _GEN_10150 = 14'h27a6 == index ? 14'h103 : _GEN_10149;
  wire [13:0] _GEN_10151 = 14'h27a7 == index ? 14'h101 : _GEN_10150;
  wire [13:0] _GEN_10152 = 14'h27a8 == index ? 14'ha7 : _GEN_10151;
  wire [13:0] _GEN_10153 = 14'h27a9 == index ? 14'ha6 : _GEN_10152;
  wire [13:0] _GEN_10154 = 14'h27aa == index ? 14'ha5 : _GEN_10153;
  wire [13:0] _GEN_10155 = 14'h27ab == index ? 14'ha4 : _GEN_10154;
  wire [13:0] _GEN_10156 = 14'h27ac == index ? 14'ha3 : _GEN_10155;
  wire [13:0] _GEN_10157 = 14'h27ad == index ? 14'ha2 : _GEN_10156;
  wire [13:0] _GEN_10158 = 14'h27ae == index ? 14'ha1 : _GEN_10157;
  wire [13:0] _GEN_10159 = 14'h27af == index ? 14'ha0 : _GEN_10158;
  wire [13:0] _GEN_10160 = 14'h27b0 == index ? 14'h9f : _GEN_10159;
  wire [13:0] _GEN_10161 = 14'h27b1 == index ? 14'h9e : _GEN_10160;
  wire [13:0] _GEN_10162 = 14'h27b2 == index ? 14'h9d : _GEN_10161;
  wire [13:0] _GEN_10163 = 14'h27b3 == index ? 14'h9c : _GEN_10162;
  wire [13:0] _GEN_10164 = 14'h27b4 == index ? 14'h9b : _GEN_10163;
  wire [13:0] _GEN_10165 = 14'h27b5 == index ? 14'h9a : _GEN_10164;
  wire [13:0] _GEN_10166 = 14'h27b6 == index ? 14'h99 : _GEN_10165;
  wire [13:0] _GEN_10167 = 14'h27b7 == index ? 14'h98 : _GEN_10166;
  wire [13:0] _GEN_10168 = 14'h27b8 == index ? 14'h97 : _GEN_10167;
  wire [13:0] _GEN_10169 = 14'h27b9 == index ? 14'h96 : _GEN_10168;
  wire [13:0] _GEN_10170 = 14'h27ba == index ? 14'h95 : _GEN_10169;
  wire [13:0] _GEN_10171 = 14'h27bb == index ? 14'h94 : _GEN_10170;
  wire [13:0] _GEN_10172 = 14'h27bc == index ? 14'h93 : _GEN_10171;
  wire [13:0] _GEN_10173 = 14'h27bd == index ? 14'h92 : _GEN_10172;
  wire [13:0] _GEN_10174 = 14'h27be == index ? 14'h91 : _GEN_10173;
  wire [13:0] _GEN_10175 = 14'h27bf == index ? 14'h90 : _GEN_10174;
  wire [13:0] _GEN_10176 = 14'h27c0 == index ? 14'h8f : _GEN_10175;
  wire [13:0] _GEN_10177 = 14'h27c1 == index ? 14'h8e : _GEN_10176;
  wire [13:0] _GEN_10178 = 14'h27c2 == index ? 14'h8d : _GEN_10177;
  wire [13:0] _GEN_10179 = 14'h27c3 == index ? 14'h8c : _GEN_10178;
  wire [13:0] _GEN_10180 = 14'h27c4 == index ? 14'h8b : _GEN_10179;
  wire [13:0] _GEN_10181 = 14'h27c5 == index ? 14'h8a : _GEN_10180;
  wire [13:0] _GEN_10182 = 14'h27c6 == index ? 14'h89 : _GEN_10181;
  wire [13:0] _GEN_10183 = 14'h27c7 == index ? 14'h88 : _GEN_10182;
  wire [13:0] _GEN_10184 = 14'h27c8 == index ? 14'h87 : _GEN_10183;
  wire [13:0] _GEN_10185 = 14'h27c9 == index ? 14'h86 : _GEN_10184;
  wire [13:0] _GEN_10186 = 14'h27ca == index ? 14'h85 : _GEN_10185;
  wire [13:0] _GEN_10187 = 14'h27cb == index ? 14'h84 : _GEN_10186;
  wire [13:0] _GEN_10188 = 14'h27cc == index ? 14'h83 : _GEN_10187;
  wire [13:0] _GEN_10189 = 14'h27cd == index ? 14'h82 : _GEN_10188;
  wire [13:0] _GEN_10190 = 14'h27ce == index ? 14'h81 : _GEN_10189;
  wire [13:0] _GEN_10191 = 14'h27cf == index ? 14'h80 : _GEN_10190;
  wire [13:0] _GEN_10192 = 14'h27d0 == index ? 14'h4f : _GEN_10191;
  wire [13:0] _GEN_10193 = 14'h27d1 == index ? 14'h4f : _GEN_10192;
  wire [13:0] _GEN_10194 = 14'h27d2 == index ? 14'h4f : _GEN_10193;
  wire [13:0] _GEN_10195 = 14'h27d3 == index ? 14'h4f : _GEN_10194;
  wire [13:0] _GEN_10196 = 14'h27d4 == index ? 14'h4f : _GEN_10195;
  wire [13:0] _GEN_10197 = 14'h27d5 == index ? 14'h4f : _GEN_10196;
  wire [13:0] _GEN_10198 = 14'h27d6 == index ? 14'h4f : _GEN_10197;
  wire [13:0] _GEN_10199 = 14'h27d7 == index ? 14'h4f : _GEN_10198;
  wire [13:0] _GEN_10200 = 14'h27d8 == index ? 14'h4f : _GEN_10199;
  wire [13:0] _GEN_10201 = 14'h27d9 == index ? 14'h4f : _GEN_10200;
  wire [13:0] _GEN_10202 = 14'h27da == index ? 14'h4f : _GEN_10201;
  wire [13:0] _GEN_10203 = 14'h27db == index ? 14'h4f : _GEN_10202;
  wire [13:0] _GEN_10204 = 14'h27dc == index ? 14'h4f : _GEN_10203;
  wire [13:0] _GEN_10205 = 14'h27dd == index ? 14'h4f : _GEN_10204;
  wire [13:0] _GEN_10206 = 14'h27de == index ? 14'h4f : _GEN_10205;
  wire [13:0] _GEN_10207 = 14'h27df == index ? 14'h4f : _GEN_10206;
  wire [13:0] _GEN_10208 = 14'h27e0 == index ? 14'h4f : _GEN_10207;
  wire [13:0] _GEN_10209 = 14'h27e1 == index ? 14'h4f : _GEN_10208;
  wire [13:0] _GEN_10210 = 14'h27e2 == index ? 14'h4f : _GEN_10209;
  wire [13:0] _GEN_10211 = 14'h27e3 == index ? 14'h4f : _GEN_10210;
  wire [13:0] _GEN_10212 = 14'h27e4 == index ? 14'h4f : _GEN_10211;
  wire [13:0] _GEN_10213 = 14'h27e5 == index ? 14'h4f : _GEN_10212;
  wire [13:0] _GEN_10214 = 14'h27e6 == index ? 14'h4f : _GEN_10213;
  wire [13:0] _GEN_10215 = 14'h27e7 == index ? 14'h4f : _GEN_10214;
  wire [13:0] _GEN_10216 = 14'h27e8 == index ? 14'h4f : _GEN_10215;
  wire [13:0] _GEN_10217 = 14'h27e9 == index ? 14'h4f : _GEN_10216;
  wire [13:0] _GEN_10218 = 14'h27ea == index ? 14'h4f : _GEN_10217;
  wire [13:0] _GEN_10219 = 14'h27eb == index ? 14'h4f : _GEN_10218;
  wire [13:0] _GEN_10220 = 14'h27ec == index ? 14'h4f : _GEN_10219;
  wire [13:0] _GEN_10221 = 14'h27ed == index ? 14'h4f : _GEN_10220;
  wire [13:0] _GEN_10222 = 14'h27ee == index ? 14'h4f : _GEN_10221;
  wire [13:0] _GEN_10223 = 14'h27ef == index ? 14'h4f : _GEN_10222;
  wire [13:0] _GEN_10224 = 14'h27f0 == index ? 14'h4f : _GEN_10223;
  wire [13:0] _GEN_10225 = 14'h27f1 == index ? 14'h4f : _GEN_10224;
  wire [13:0] _GEN_10226 = 14'h27f2 == index ? 14'h4f : _GEN_10225;
  wire [13:0] _GEN_10227 = 14'h27f3 == index ? 14'h4f : _GEN_10226;
  wire [13:0] _GEN_10228 = 14'h27f4 == index ? 14'h4f : _GEN_10227;
  wire [13:0] _GEN_10229 = 14'h27f5 == index ? 14'h4f : _GEN_10228;
  wire [13:0] _GEN_10230 = 14'h27f6 == index ? 14'h4f : _GEN_10229;
  wire [13:0] _GEN_10231 = 14'h27f7 == index ? 14'h4f : _GEN_10230;
  wire [13:0] _GEN_10232 = 14'h27f8 == index ? 14'h4f : _GEN_10231;
  wire [13:0] _GEN_10233 = 14'h27f9 == index ? 14'h4f : _GEN_10232;
  wire [13:0] _GEN_10234 = 14'h27fa == index ? 14'h4f : _GEN_10233;
  wire [13:0] _GEN_10235 = 14'h27fb == index ? 14'h4f : _GEN_10234;
  wire [13:0] _GEN_10236 = 14'h27fc == index ? 14'h4f : _GEN_10235;
  wire [13:0] _GEN_10237 = 14'h27fd == index ? 14'h4f : _GEN_10236;
  wire [13:0] _GEN_10238 = 14'h27fe == index ? 14'h4f : _GEN_10237;
  wire [13:0] _GEN_10239 = 14'h27ff == index ? 14'h4f : _GEN_10238;
  wire [13:0] _GEN_10240 = 14'h2800 == index ? 14'h0 : _GEN_10239;
  wire [13:0] _GEN_10241 = 14'h2801 == index ? 14'h2800 : _GEN_10240;
  wire [13:0] _GEN_10242 = 14'h2802 == index ? 14'h1400 : _GEN_10241;
  wire [13:0] _GEN_10243 = 14'h2803 == index ? 14'hd02 : _GEN_10242;
  wire [13:0] _GEN_10244 = 14'h2804 == index ? 14'ha00 : _GEN_10243;
  wire [13:0] _GEN_10245 = 14'h2805 == index ? 14'h800 : _GEN_10244;
  wire [13:0] _GEN_10246 = 14'h2806 == index ? 14'h682 : _GEN_10245;
  wire [13:0] _GEN_10247 = 14'h2807 == index ? 14'h583 : _GEN_10246;
  wire [13:0] _GEN_10248 = 14'h2808 == index ? 14'h500 : _GEN_10247;
  wire [13:0] _GEN_10249 = 14'h2809 == index ? 14'h408 : _GEN_10248;
  wire [13:0] _GEN_10250 = 14'h280a == index ? 14'h400 : _GEN_10249;
  wire [13:0] _GEN_10251 = 14'h280b == index ? 14'h383 : _GEN_10250;
  wire [13:0] _GEN_10252 = 14'h280c == index ? 14'h308 : _GEN_10251;
  wire [13:0] _GEN_10253 = 14'h280d == index ? 14'h302 : _GEN_10252;
  wire [13:0] _GEN_10254 = 14'h280e == index ? 14'h28a : _GEN_10253;
  wire [13:0] _GEN_10255 = 14'h280f == index ? 14'h285 : _GEN_10254;
  wire [13:0] _GEN_10256 = 14'h2810 == index ? 14'h280 : _GEN_10255;
  wire [13:0] _GEN_10257 = 14'h2811 == index ? 14'h20c : _GEN_10256;
  wire [13:0] _GEN_10258 = 14'h2812 == index ? 14'h208 : _GEN_10257;
  wire [13:0] _GEN_10259 = 14'h2813 == index ? 14'h204 : _GEN_10258;
  wire [13:0] _GEN_10260 = 14'h2814 == index ? 14'h200 : _GEN_10259;
  wire [13:0] _GEN_10261 = 14'h2815 == index ? 14'h191 : _GEN_10260;
  wire [13:0] _GEN_10262 = 14'h2816 == index ? 14'h18e : _GEN_10261;
  wire [13:0] _GEN_10263 = 14'h2817 == index ? 14'h18b : _GEN_10262;
  wire [13:0] _GEN_10264 = 14'h2818 == index ? 14'h188 : _GEN_10263;
  wire [13:0] _GEN_10265 = 14'h2819 == index ? 14'h185 : _GEN_10264;
  wire [13:0] _GEN_10266 = 14'h281a == index ? 14'h182 : _GEN_10265;
  wire [13:0] _GEN_10267 = 14'h281b == index ? 14'h11a : _GEN_10266;
  wire [13:0] _GEN_10268 = 14'h281c == index ? 14'h118 : _GEN_10267;
  wire [13:0] _GEN_10269 = 14'h281d == index ? 14'h116 : _GEN_10268;
  wire [13:0] _GEN_10270 = 14'h281e == index ? 14'h114 : _GEN_10269;
  wire [13:0] _GEN_10271 = 14'h281f == index ? 14'h112 : _GEN_10270;
  wire [13:0] _GEN_10272 = 14'h2820 == index ? 14'h110 : _GEN_10271;
  wire [13:0] _GEN_10273 = 14'h2821 == index ? 14'h10e : _GEN_10272;
  wire [13:0] _GEN_10274 = 14'h2822 == index ? 14'h10c : _GEN_10273;
  wire [13:0] _GEN_10275 = 14'h2823 == index ? 14'h10a : _GEN_10274;
  wire [13:0] _GEN_10276 = 14'h2824 == index ? 14'h108 : _GEN_10275;
  wire [13:0] _GEN_10277 = 14'h2825 == index ? 14'h106 : _GEN_10276;
  wire [13:0] _GEN_10278 = 14'h2826 == index ? 14'h104 : _GEN_10277;
  wire [13:0] _GEN_10279 = 14'h2827 == index ? 14'h102 : _GEN_10278;
  wire [13:0] _GEN_10280 = 14'h2828 == index ? 14'h100 : _GEN_10279;
  wire [13:0] _GEN_10281 = 14'h2829 == index ? 14'ha7 : _GEN_10280;
  wire [13:0] _GEN_10282 = 14'h282a == index ? 14'ha6 : _GEN_10281;
  wire [13:0] _GEN_10283 = 14'h282b == index ? 14'ha5 : _GEN_10282;
  wire [13:0] _GEN_10284 = 14'h282c == index ? 14'ha4 : _GEN_10283;
  wire [13:0] _GEN_10285 = 14'h282d == index ? 14'ha3 : _GEN_10284;
  wire [13:0] _GEN_10286 = 14'h282e == index ? 14'ha2 : _GEN_10285;
  wire [13:0] _GEN_10287 = 14'h282f == index ? 14'ha1 : _GEN_10286;
  wire [13:0] _GEN_10288 = 14'h2830 == index ? 14'ha0 : _GEN_10287;
  wire [13:0] _GEN_10289 = 14'h2831 == index ? 14'h9f : _GEN_10288;
  wire [13:0] _GEN_10290 = 14'h2832 == index ? 14'h9e : _GEN_10289;
  wire [13:0] _GEN_10291 = 14'h2833 == index ? 14'h9d : _GEN_10290;
  wire [13:0] _GEN_10292 = 14'h2834 == index ? 14'h9c : _GEN_10291;
  wire [13:0] _GEN_10293 = 14'h2835 == index ? 14'h9b : _GEN_10292;
  wire [13:0] _GEN_10294 = 14'h2836 == index ? 14'h9a : _GEN_10293;
  wire [13:0] _GEN_10295 = 14'h2837 == index ? 14'h99 : _GEN_10294;
  wire [13:0] _GEN_10296 = 14'h2838 == index ? 14'h98 : _GEN_10295;
  wire [13:0] _GEN_10297 = 14'h2839 == index ? 14'h97 : _GEN_10296;
  wire [13:0] _GEN_10298 = 14'h283a == index ? 14'h96 : _GEN_10297;
  wire [13:0] _GEN_10299 = 14'h283b == index ? 14'h95 : _GEN_10298;
  wire [13:0] _GEN_10300 = 14'h283c == index ? 14'h94 : _GEN_10299;
  wire [13:0] _GEN_10301 = 14'h283d == index ? 14'h93 : _GEN_10300;
  wire [13:0] _GEN_10302 = 14'h283e == index ? 14'h92 : _GEN_10301;
  wire [13:0] _GEN_10303 = 14'h283f == index ? 14'h91 : _GEN_10302;
  wire [13:0] _GEN_10304 = 14'h2840 == index ? 14'h90 : _GEN_10303;
  wire [13:0] _GEN_10305 = 14'h2841 == index ? 14'h8f : _GEN_10304;
  wire [13:0] _GEN_10306 = 14'h2842 == index ? 14'h8e : _GEN_10305;
  wire [13:0] _GEN_10307 = 14'h2843 == index ? 14'h8d : _GEN_10306;
  wire [13:0] _GEN_10308 = 14'h2844 == index ? 14'h8c : _GEN_10307;
  wire [13:0] _GEN_10309 = 14'h2845 == index ? 14'h8b : _GEN_10308;
  wire [13:0] _GEN_10310 = 14'h2846 == index ? 14'h8a : _GEN_10309;
  wire [13:0] _GEN_10311 = 14'h2847 == index ? 14'h89 : _GEN_10310;
  wire [13:0] _GEN_10312 = 14'h2848 == index ? 14'h88 : _GEN_10311;
  wire [13:0] _GEN_10313 = 14'h2849 == index ? 14'h87 : _GEN_10312;
  wire [13:0] _GEN_10314 = 14'h284a == index ? 14'h86 : _GEN_10313;
  wire [13:0] _GEN_10315 = 14'h284b == index ? 14'h85 : _GEN_10314;
  wire [13:0] _GEN_10316 = 14'h284c == index ? 14'h84 : _GEN_10315;
  wire [13:0] _GEN_10317 = 14'h284d == index ? 14'h83 : _GEN_10316;
  wire [13:0] _GEN_10318 = 14'h284e == index ? 14'h82 : _GEN_10317;
  wire [13:0] _GEN_10319 = 14'h284f == index ? 14'h81 : _GEN_10318;
  wire [13:0] _GEN_10320 = 14'h2850 == index ? 14'h80 : _GEN_10319;
  wire [13:0] _GEN_10321 = 14'h2851 == index ? 14'h50 : _GEN_10320;
  wire [13:0] _GEN_10322 = 14'h2852 == index ? 14'h50 : _GEN_10321;
  wire [13:0] _GEN_10323 = 14'h2853 == index ? 14'h50 : _GEN_10322;
  wire [13:0] _GEN_10324 = 14'h2854 == index ? 14'h50 : _GEN_10323;
  wire [13:0] _GEN_10325 = 14'h2855 == index ? 14'h50 : _GEN_10324;
  wire [13:0] _GEN_10326 = 14'h2856 == index ? 14'h50 : _GEN_10325;
  wire [13:0] _GEN_10327 = 14'h2857 == index ? 14'h50 : _GEN_10326;
  wire [13:0] _GEN_10328 = 14'h2858 == index ? 14'h50 : _GEN_10327;
  wire [13:0] _GEN_10329 = 14'h2859 == index ? 14'h50 : _GEN_10328;
  wire [13:0] _GEN_10330 = 14'h285a == index ? 14'h50 : _GEN_10329;
  wire [13:0] _GEN_10331 = 14'h285b == index ? 14'h50 : _GEN_10330;
  wire [13:0] _GEN_10332 = 14'h285c == index ? 14'h50 : _GEN_10331;
  wire [13:0] _GEN_10333 = 14'h285d == index ? 14'h50 : _GEN_10332;
  wire [13:0] _GEN_10334 = 14'h285e == index ? 14'h50 : _GEN_10333;
  wire [13:0] _GEN_10335 = 14'h285f == index ? 14'h50 : _GEN_10334;
  wire [13:0] _GEN_10336 = 14'h2860 == index ? 14'h50 : _GEN_10335;
  wire [13:0] _GEN_10337 = 14'h2861 == index ? 14'h50 : _GEN_10336;
  wire [13:0] _GEN_10338 = 14'h2862 == index ? 14'h50 : _GEN_10337;
  wire [13:0] _GEN_10339 = 14'h2863 == index ? 14'h50 : _GEN_10338;
  wire [13:0] _GEN_10340 = 14'h2864 == index ? 14'h50 : _GEN_10339;
  wire [13:0] _GEN_10341 = 14'h2865 == index ? 14'h50 : _GEN_10340;
  wire [13:0] _GEN_10342 = 14'h2866 == index ? 14'h50 : _GEN_10341;
  wire [13:0] _GEN_10343 = 14'h2867 == index ? 14'h50 : _GEN_10342;
  wire [13:0] _GEN_10344 = 14'h2868 == index ? 14'h50 : _GEN_10343;
  wire [13:0] _GEN_10345 = 14'h2869 == index ? 14'h50 : _GEN_10344;
  wire [13:0] _GEN_10346 = 14'h286a == index ? 14'h50 : _GEN_10345;
  wire [13:0] _GEN_10347 = 14'h286b == index ? 14'h50 : _GEN_10346;
  wire [13:0] _GEN_10348 = 14'h286c == index ? 14'h50 : _GEN_10347;
  wire [13:0] _GEN_10349 = 14'h286d == index ? 14'h50 : _GEN_10348;
  wire [13:0] _GEN_10350 = 14'h286e == index ? 14'h50 : _GEN_10349;
  wire [13:0] _GEN_10351 = 14'h286f == index ? 14'h50 : _GEN_10350;
  wire [13:0] _GEN_10352 = 14'h2870 == index ? 14'h50 : _GEN_10351;
  wire [13:0] _GEN_10353 = 14'h2871 == index ? 14'h50 : _GEN_10352;
  wire [13:0] _GEN_10354 = 14'h2872 == index ? 14'h50 : _GEN_10353;
  wire [13:0] _GEN_10355 = 14'h2873 == index ? 14'h50 : _GEN_10354;
  wire [13:0] _GEN_10356 = 14'h2874 == index ? 14'h50 : _GEN_10355;
  wire [13:0] _GEN_10357 = 14'h2875 == index ? 14'h50 : _GEN_10356;
  wire [13:0] _GEN_10358 = 14'h2876 == index ? 14'h50 : _GEN_10357;
  wire [13:0] _GEN_10359 = 14'h2877 == index ? 14'h50 : _GEN_10358;
  wire [13:0] _GEN_10360 = 14'h2878 == index ? 14'h50 : _GEN_10359;
  wire [13:0] _GEN_10361 = 14'h2879 == index ? 14'h50 : _GEN_10360;
  wire [13:0] _GEN_10362 = 14'h287a == index ? 14'h50 : _GEN_10361;
  wire [13:0] _GEN_10363 = 14'h287b == index ? 14'h50 : _GEN_10362;
  wire [13:0] _GEN_10364 = 14'h287c == index ? 14'h50 : _GEN_10363;
  wire [13:0] _GEN_10365 = 14'h287d == index ? 14'h50 : _GEN_10364;
  wire [13:0] _GEN_10366 = 14'h287e == index ? 14'h50 : _GEN_10365;
  wire [13:0] _GEN_10367 = 14'h287f == index ? 14'h50 : _GEN_10366;
  wire [13:0] _GEN_10368 = 14'h2880 == index ? 14'h0 : _GEN_10367;
  wire [13:0] _GEN_10369 = 14'h2881 == index ? 14'h2880 : _GEN_10368;
  wire [13:0] _GEN_10370 = 14'h2882 == index ? 14'h1401 : _GEN_10369;
  wire [13:0] _GEN_10371 = 14'h2883 == index ? 14'hd80 : _GEN_10370;
  wire [13:0] _GEN_10372 = 14'h2884 == index ? 14'ha01 : _GEN_10371;
  wire [13:0] _GEN_10373 = 14'h2885 == index ? 14'h801 : _GEN_10372;
  wire [13:0] _GEN_10374 = 14'h2886 == index ? 14'h683 : _GEN_10373;
  wire [13:0] _GEN_10375 = 14'h2887 == index ? 14'h584 : _GEN_10374;
  wire [13:0] _GEN_10376 = 14'h2888 == index ? 14'h501 : _GEN_10375;
  wire [13:0] _GEN_10377 = 14'h2889 == index ? 14'h480 : _GEN_10376;
  wire [13:0] _GEN_10378 = 14'h288a == index ? 14'h401 : _GEN_10377;
  wire [13:0] _GEN_10379 = 14'h288b == index ? 14'h384 : _GEN_10378;
  wire [13:0] _GEN_10380 = 14'h288c == index ? 14'h309 : _GEN_10379;
  wire [13:0] _GEN_10381 = 14'h288d == index ? 14'h303 : _GEN_10380;
  wire [13:0] _GEN_10382 = 14'h288e == index ? 14'h28b : _GEN_10381;
  wire [13:0] _GEN_10383 = 14'h288f == index ? 14'h286 : _GEN_10382;
  wire [13:0] _GEN_10384 = 14'h2890 == index ? 14'h281 : _GEN_10383;
  wire [13:0] _GEN_10385 = 14'h2891 == index ? 14'h20d : _GEN_10384;
  wire [13:0] _GEN_10386 = 14'h2892 == index ? 14'h209 : _GEN_10385;
  wire [13:0] _GEN_10387 = 14'h2893 == index ? 14'h205 : _GEN_10386;
  wire [13:0] _GEN_10388 = 14'h2894 == index ? 14'h201 : _GEN_10387;
  wire [13:0] _GEN_10389 = 14'h2895 == index ? 14'h192 : _GEN_10388;
  wire [13:0] _GEN_10390 = 14'h2896 == index ? 14'h18f : _GEN_10389;
  wire [13:0] _GEN_10391 = 14'h2897 == index ? 14'h18c : _GEN_10390;
  wire [13:0] _GEN_10392 = 14'h2898 == index ? 14'h189 : _GEN_10391;
  wire [13:0] _GEN_10393 = 14'h2899 == index ? 14'h186 : _GEN_10392;
  wire [13:0] _GEN_10394 = 14'h289a == index ? 14'h183 : _GEN_10393;
  wire [13:0] _GEN_10395 = 14'h289b == index ? 14'h180 : _GEN_10394;
  wire [13:0] _GEN_10396 = 14'h289c == index ? 14'h119 : _GEN_10395;
  wire [13:0] _GEN_10397 = 14'h289d == index ? 14'h117 : _GEN_10396;
  wire [13:0] _GEN_10398 = 14'h289e == index ? 14'h115 : _GEN_10397;
  wire [13:0] _GEN_10399 = 14'h289f == index ? 14'h113 : _GEN_10398;
  wire [13:0] _GEN_10400 = 14'h28a0 == index ? 14'h111 : _GEN_10399;
  wire [13:0] _GEN_10401 = 14'h28a1 == index ? 14'h10f : _GEN_10400;
  wire [13:0] _GEN_10402 = 14'h28a2 == index ? 14'h10d : _GEN_10401;
  wire [13:0] _GEN_10403 = 14'h28a3 == index ? 14'h10b : _GEN_10402;
  wire [13:0] _GEN_10404 = 14'h28a4 == index ? 14'h109 : _GEN_10403;
  wire [13:0] _GEN_10405 = 14'h28a5 == index ? 14'h107 : _GEN_10404;
  wire [13:0] _GEN_10406 = 14'h28a6 == index ? 14'h105 : _GEN_10405;
  wire [13:0] _GEN_10407 = 14'h28a7 == index ? 14'h103 : _GEN_10406;
  wire [13:0] _GEN_10408 = 14'h28a8 == index ? 14'h101 : _GEN_10407;
  wire [13:0] _GEN_10409 = 14'h28a9 == index ? 14'ha8 : _GEN_10408;
  wire [13:0] _GEN_10410 = 14'h28aa == index ? 14'ha7 : _GEN_10409;
  wire [13:0] _GEN_10411 = 14'h28ab == index ? 14'ha6 : _GEN_10410;
  wire [13:0] _GEN_10412 = 14'h28ac == index ? 14'ha5 : _GEN_10411;
  wire [13:0] _GEN_10413 = 14'h28ad == index ? 14'ha4 : _GEN_10412;
  wire [13:0] _GEN_10414 = 14'h28ae == index ? 14'ha3 : _GEN_10413;
  wire [13:0] _GEN_10415 = 14'h28af == index ? 14'ha2 : _GEN_10414;
  wire [13:0] _GEN_10416 = 14'h28b0 == index ? 14'ha1 : _GEN_10415;
  wire [13:0] _GEN_10417 = 14'h28b1 == index ? 14'ha0 : _GEN_10416;
  wire [13:0] _GEN_10418 = 14'h28b2 == index ? 14'h9f : _GEN_10417;
  wire [13:0] _GEN_10419 = 14'h28b3 == index ? 14'h9e : _GEN_10418;
  wire [13:0] _GEN_10420 = 14'h28b4 == index ? 14'h9d : _GEN_10419;
  wire [13:0] _GEN_10421 = 14'h28b5 == index ? 14'h9c : _GEN_10420;
  wire [13:0] _GEN_10422 = 14'h28b6 == index ? 14'h9b : _GEN_10421;
  wire [13:0] _GEN_10423 = 14'h28b7 == index ? 14'h9a : _GEN_10422;
  wire [13:0] _GEN_10424 = 14'h28b8 == index ? 14'h99 : _GEN_10423;
  wire [13:0] _GEN_10425 = 14'h28b9 == index ? 14'h98 : _GEN_10424;
  wire [13:0] _GEN_10426 = 14'h28ba == index ? 14'h97 : _GEN_10425;
  wire [13:0] _GEN_10427 = 14'h28bb == index ? 14'h96 : _GEN_10426;
  wire [13:0] _GEN_10428 = 14'h28bc == index ? 14'h95 : _GEN_10427;
  wire [13:0] _GEN_10429 = 14'h28bd == index ? 14'h94 : _GEN_10428;
  wire [13:0] _GEN_10430 = 14'h28be == index ? 14'h93 : _GEN_10429;
  wire [13:0] _GEN_10431 = 14'h28bf == index ? 14'h92 : _GEN_10430;
  wire [13:0] _GEN_10432 = 14'h28c0 == index ? 14'h91 : _GEN_10431;
  wire [13:0] _GEN_10433 = 14'h28c1 == index ? 14'h90 : _GEN_10432;
  wire [13:0] _GEN_10434 = 14'h28c2 == index ? 14'h8f : _GEN_10433;
  wire [13:0] _GEN_10435 = 14'h28c3 == index ? 14'h8e : _GEN_10434;
  wire [13:0] _GEN_10436 = 14'h28c4 == index ? 14'h8d : _GEN_10435;
  wire [13:0] _GEN_10437 = 14'h28c5 == index ? 14'h8c : _GEN_10436;
  wire [13:0] _GEN_10438 = 14'h28c6 == index ? 14'h8b : _GEN_10437;
  wire [13:0] _GEN_10439 = 14'h28c7 == index ? 14'h8a : _GEN_10438;
  wire [13:0] _GEN_10440 = 14'h28c8 == index ? 14'h89 : _GEN_10439;
  wire [13:0] _GEN_10441 = 14'h28c9 == index ? 14'h88 : _GEN_10440;
  wire [13:0] _GEN_10442 = 14'h28ca == index ? 14'h87 : _GEN_10441;
  wire [13:0] _GEN_10443 = 14'h28cb == index ? 14'h86 : _GEN_10442;
  wire [13:0] _GEN_10444 = 14'h28cc == index ? 14'h85 : _GEN_10443;
  wire [13:0] _GEN_10445 = 14'h28cd == index ? 14'h84 : _GEN_10444;
  wire [13:0] _GEN_10446 = 14'h28ce == index ? 14'h83 : _GEN_10445;
  wire [13:0] _GEN_10447 = 14'h28cf == index ? 14'h82 : _GEN_10446;
  wire [13:0] _GEN_10448 = 14'h28d0 == index ? 14'h81 : _GEN_10447;
  wire [13:0] _GEN_10449 = 14'h28d1 == index ? 14'h80 : _GEN_10448;
  wire [13:0] _GEN_10450 = 14'h28d2 == index ? 14'h51 : _GEN_10449;
  wire [13:0] _GEN_10451 = 14'h28d3 == index ? 14'h51 : _GEN_10450;
  wire [13:0] _GEN_10452 = 14'h28d4 == index ? 14'h51 : _GEN_10451;
  wire [13:0] _GEN_10453 = 14'h28d5 == index ? 14'h51 : _GEN_10452;
  wire [13:0] _GEN_10454 = 14'h28d6 == index ? 14'h51 : _GEN_10453;
  wire [13:0] _GEN_10455 = 14'h28d7 == index ? 14'h51 : _GEN_10454;
  wire [13:0] _GEN_10456 = 14'h28d8 == index ? 14'h51 : _GEN_10455;
  wire [13:0] _GEN_10457 = 14'h28d9 == index ? 14'h51 : _GEN_10456;
  wire [13:0] _GEN_10458 = 14'h28da == index ? 14'h51 : _GEN_10457;
  wire [13:0] _GEN_10459 = 14'h28db == index ? 14'h51 : _GEN_10458;
  wire [13:0] _GEN_10460 = 14'h28dc == index ? 14'h51 : _GEN_10459;
  wire [13:0] _GEN_10461 = 14'h28dd == index ? 14'h51 : _GEN_10460;
  wire [13:0] _GEN_10462 = 14'h28de == index ? 14'h51 : _GEN_10461;
  wire [13:0] _GEN_10463 = 14'h28df == index ? 14'h51 : _GEN_10462;
  wire [13:0] _GEN_10464 = 14'h28e0 == index ? 14'h51 : _GEN_10463;
  wire [13:0] _GEN_10465 = 14'h28e1 == index ? 14'h51 : _GEN_10464;
  wire [13:0] _GEN_10466 = 14'h28e2 == index ? 14'h51 : _GEN_10465;
  wire [13:0] _GEN_10467 = 14'h28e3 == index ? 14'h51 : _GEN_10466;
  wire [13:0] _GEN_10468 = 14'h28e4 == index ? 14'h51 : _GEN_10467;
  wire [13:0] _GEN_10469 = 14'h28e5 == index ? 14'h51 : _GEN_10468;
  wire [13:0] _GEN_10470 = 14'h28e6 == index ? 14'h51 : _GEN_10469;
  wire [13:0] _GEN_10471 = 14'h28e7 == index ? 14'h51 : _GEN_10470;
  wire [13:0] _GEN_10472 = 14'h28e8 == index ? 14'h51 : _GEN_10471;
  wire [13:0] _GEN_10473 = 14'h28e9 == index ? 14'h51 : _GEN_10472;
  wire [13:0] _GEN_10474 = 14'h28ea == index ? 14'h51 : _GEN_10473;
  wire [13:0] _GEN_10475 = 14'h28eb == index ? 14'h51 : _GEN_10474;
  wire [13:0] _GEN_10476 = 14'h28ec == index ? 14'h51 : _GEN_10475;
  wire [13:0] _GEN_10477 = 14'h28ed == index ? 14'h51 : _GEN_10476;
  wire [13:0] _GEN_10478 = 14'h28ee == index ? 14'h51 : _GEN_10477;
  wire [13:0] _GEN_10479 = 14'h28ef == index ? 14'h51 : _GEN_10478;
  wire [13:0] _GEN_10480 = 14'h28f0 == index ? 14'h51 : _GEN_10479;
  wire [13:0] _GEN_10481 = 14'h28f1 == index ? 14'h51 : _GEN_10480;
  wire [13:0] _GEN_10482 = 14'h28f2 == index ? 14'h51 : _GEN_10481;
  wire [13:0] _GEN_10483 = 14'h28f3 == index ? 14'h51 : _GEN_10482;
  wire [13:0] _GEN_10484 = 14'h28f4 == index ? 14'h51 : _GEN_10483;
  wire [13:0] _GEN_10485 = 14'h28f5 == index ? 14'h51 : _GEN_10484;
  wire [13:0] _GEN_10486 = 14'h28f6 == index ? 14'h51 : _GEN_10485;
  wire [13:0] _GEN_10487 = 14'h28f7 == index ? 14'h51 : _GEN_10486;
  wire [13:0] _GEN_10488 = 14'h28f8 == index ? 14'h51 : _GEN_10487;
  wire [13:0] _GEN_10489 = 14'h28f9 == index ? 14'h51 : _GEN_10488;
  wire [13:0] _GEN_10490 = 14'h28fa == index ? 14'h51 : _GEN_10489;
  wire [13:0] _GEN_10491 = 14'h28fb == index ? 14'h51 : _GEN_10490;
  wire [13:0] _GEN_10492 = 14'h28fc == index ? 14'h51 : _GEN_10491;
  wire [13:0] _GEN_10493 = 14'h28fd == index ? 14'h51 : _GEN_10492;
  wire [13:0] _GEN_10494 = 14'h28fe == index ? 14'h51 : _GEN_10493;
  wire [13:0] _GEN_10495 = 14'h28ff == index ? 14'h51 : _GEN_10494;
  wire [13:0] _GEN_10496 = 14'h2900 == index ? 14'h0 : _GEN_10495;
  wire [13:0] _GEN_10497 = 14'h2901 == index ? 14'h2900 : _GEN_10496;
  wire [13:0] _GEN_10498 = 14'h2902 == index ? 14'h1480 : _GEN_10497;
  wire [13:0] _GEN_10499 = 14'h2903 == index ? 14'hd81 : _GEN_10498;
  wire [13:0] _GEN_10500 = 14'h2904 == index ? 14'ha02 : _GEN_10499;
  wire [13:0] _GEN_10501 = 14'h2905 == index ? 14'h802 : _GEN_10500;
  wire [13:0] _GEN_10502 = 14'h2906 == index ? 14'h684 : _GEN_10501;
  wire [13:0] _GEN_10503 = 14'h2907 == index ? 14'h585 : _GEN_10502;
  wire [13:0] _GEN_10504 = 14'h2908 == index ? 14'h502 : _GEN_10503;
  wire [13:0] _GEN_10505 = 14'h2909 == index ? 14'h481 : _GEN_10504;
  wire [13:0] _GEN_10506 = 14'h290a == index ? 14'h402 : _GEN_10505;
  wire [13:0] _GEN_10507 = 14'h290b == index ? 14'h385 : _GEN_10506;
  wire [13:0] _GEN_10508 = 14'h290c == index ? 14'h30a : _GEN_10507;
  wire [13:0] _GEN_10509 = 14'h290d == index ? 14'h304 : _GEN_10508;
  wire [13:0] _GEN_10510 = 14'h290e == index ? 14'h28c : _GEN_10509;
  wire [13:0] _GEN_10511 = 14'h290f == index ? 14'h287 : _GEN_10510;
  wire [13:0] _GEN_10512 = 14'h2910 == index ? 14'h282 : _GEN_10511;
  wire [13:0] _GEN_10513 = 14'h2911 == index ? 14'h20e : _GEN_10512;
  wire [13:0] _GEN_10514 = 14'h2912 == index ? 14'h20a : _GEN_10513;
  wire [13:0] _GEN_10515 = 14'h2913 == index ? 14'h206 : _GEN_10514;
  wire [13:0] _GEN_10516 = 14'h2914 == index ? 14'h202 : _GEN_10515;
  wire [13:0] _GEN_10517 = 14'h2915 == index ? 14'h193 : _GEN_10516;
  wire [13:0] _GEN_10518 = 14'h2916 == index ? 14'h190 : _GEN_10517;
  wire [13:0] _GEN_10519 = 14'h2917 == index ? 14'h18d : _GEN_10518;
  wire [13:0] _GEN_10520 = 14'h2918 == index ? 14'h18a : _GEN_10519;
  wire [13:0] _GEN_10521 = 14'h2919 == index ? 14'h187 : _GEN_10520;
  wire [13:0] _GEN_10522 = 14'h291a == index ? 14'h184 : _GEN_10521;
  wire [13:0] _GEN_10523 = 14'h291b == index ? 14'h181 : _GEN_10522;
  wire [13:0] _GEN_10524 = 14'h291c == index ? 14'h11a : _GEN_10523;
  wire [13:0] _GEN_10525 = 14'h291d == index ? 14'h118 : _GEN_10524;
  wire [13:0] _GEN_10526 = 14'h291e == index ? 14'h116 : _GEN_10525;
  wire [13:0] _GEN_10527 = 14'h291f == index ? 14'h114 : _GEN_10526;
  wire [13:0] _GEN_10528 = 14'h2920 == index ? 14'h112 : _GEN_10527;
  wire [13:0] _GEN_10529 = 14'h2921 == index ? 14'h110 : _GEN_10528;
  wire [13:0] _GEN_10530 = 14'h2922 == index ? 14'h10e : _GEN_10529;
  wire [13:0] _GEN_10531 = 14'h2923 == index ? 14'h10c : _GEN_10530;
  wire [13:0] _GEN_10532 = 14'h2924 == index ? 14'h10a : _GEN_10531;
  wire [13:0] _GEN_10533 = 14'h2925 == index ? 14'h108 : _GEN_10532;
  wire [13:0] _GEN_10534 = 14'h2926 == index ? 14'h106 : _GEN_10533;
  wire [13:0] _GEN_10535 = 14'h2927 == index ? 14'h104 : _GEN_10534;
  wire [13:0] _GEN_10536 = 14'h2928 == index ? 14'h102 : _GEN_10535;
  wire [13:0] _GEN_10537 = 14'h2929 == index ? 14'h100 : _GEN_10536;
  wire [13:0] _GEN_10538 = 14'h292a == index ? 14'ha8 : _GEN_10537;
  wire [13:0] _GEN_10539 = 14'h292b == index ? 14'ha7 : _GEN_10538;
  wire [13:0] _GEN_10540 = 14'h292c == index ? 14'ha6 : _GEN_10539;
  wire [13:0] _GEN_10541 = 14'h292d == index ? 14'ha5 : _GEN_10540;
  wire [13:0] _GEN_10542 = 14'h292e == index ? 14'ha4 : _GEN_10541;
  wire [13:0] _GEN_10543 = 14'h292f == index ? 14'ha3 : _GEN_10542;
  wire [13:0] _GEN_10544 = 14'h2930 == index ? 14'ha2 : _GEN_10543;
  wire [13:0] _GEN_10545 = 14'h2931 == index ? 14'ha1 : _GEN_10544;
  wire [13:0] _GEN_10546 = 14'h2932 == index ? 14'ha0 : _GEN_10545;
  wire [13:0] _GEN_10547 = 14'h2933 == index ? 14'h9f : _GEN_10546;
  wire [13:0] _GEN_10548 = 14'h2934 == index ? 14'h9e : _GEN_10547;
  wire [13:0] _GEN_10549 = 14'h2935 == index ? 14'h9d : _GEN_10548;
  wire [13:0] _GEN_10550 = 14'h2936 == index ? 14'h9c : _GEN_10549;
  wire [13:0] _GEN_10551 = 14'h2937 == index ? 14'h9b : _GEN_10550;
  wire [13:0] _GEN_10552 = 14'h2938 == index ? 14'h9a : _GEN_10551;
  wire [13:0] _GEN_10553 = 14'h2939 == index ? 14'h99 : _GEN_10552;
  wire [13:0] _GEN_10554 = 14'h293a == index ? 14'h98 : _GEN_10553;
  wire [13:0] _GEN_10555 = 14'h293b == index ? 14'h97 : _GEN_10554;
  wire [13:0] _GEN_10556 = 14'h293c == index ? 14'h96 : _GEN_10555;
  wire [13:0] _GEN_10557 = 14'h293d == index ? 14'h95 : _GEN_10556;
  wire [13:0] _GEN_10558 = 14'h293e == index ? 14'h94 : _GEN_10557;
  wire [13:0] _GEN_10559 = 14'h293f == index ? 14'h93 : _GEN_10558;
  wire [13:0] _GEN_10560 = 14'h2940 == index ? 14'h92 : _GEN_10559;
  wire [13:0] _GEN_10561 = 14'h2941 == index ? 14'h91 : _GEN_10560;
  wire [13:0] _GEN_10562 = 14'h2942 == index ? 14'h90 : _GEN_10561;
  wire [13:0] _GEN_10563 = 14'h2943 == index ? 14'h8f : _GEN_10562;
  wire [13:0] _GEN_10564 = 14'h2944 == index ? 14'h8e : _GEN_10563;
  wire [13:0] _GEN_10565 = 14'h2945 == index ? 14'h8d : _GEN_10564;
  wire [13:0] _GEN_10566 = 14'h2946 == index ? 14'h8c : _GEN_10565;
  wire [13:0] _GEN_10567 = 14'h2947 == index ? 14'h8b : _GEN_10566;
  wire [13:0] _GEN_10568 = 14'h2948 == index ? 14'h8a : _GEN_10567;
  wire [13:0] _GEN_10569 = 14'h2949 == index ? 14'h89 : _GEN_10568;
  wire [13:0] _GEN_10570 = 14'h294a == index ? 14'h88 : _GEN_10569;
  wire [13:0] _GEN_10571 = 14'h294b == index ? 14'h87 : _GEN_10570;
  wire [13:0] _GEN_10572 = 14'h294c == index ? 14'h86 : _GEN_10571;
  wire [13:0] _GEN_10573 = 14'h294d == index ? 14'h85 : _GEN_10572;
  wire [13:0] _GEN_10574 = 14'h294e == index ? 14'h84 : _GEN_10573;
  wire [13:0] _GEN_10575 = 14'h294f == index ? 14'h83 : _GEN_10574;
  wire [13:0] _GEN_10576 = 14'h2950 == index ? 14'h82 : _GEN_10575;
  wire [13:0] _GEN_10577 = 14'h2951 == index ? 14'h81 : _GEN_10576;
  wire [13:0] _GEN_10578 = 14'h2952 == index ? 14'h80 : _GEN_10577;
  wire [13:0] _GEN_10579 = 14'h2953 == index ? 14'h52 : _GEN_10578;
  wire [13:0] _GEN_10580 = 14'h2954 == index ? 14'h52 : _GEN_10579;
  wire [13:0] _GEN_10581 = 14'h2955 == index ? 14'h52 : _GEN_10580;
  wire [13:0] _GEN_10582 = 14'h2956 == index ? 14'h52 : _GEN_10581;
  wire [13:0] _GEN_10583 = 14'h2957 == index ? 14'h52 : _GEN_10582;
  wire [13:0] _GEN_10584 = 14'h2958 == index ? 14'h52 : _GEN_10583;
  wire [13:0] _GEN_10585 = 14'h2959 == index ? 14'h52 : _GEN_10584;
  wire [13:0] _GEN_10586 = 14'h295a == index ? 14'h52 : _GEN_10585;
  wire [13:0] _GEN_10587 = 14'h295b == index ? 14'h52 : _GEN_10586;
  wire [13:0] _GEN_10588 = 14'h295c == index ? 14'h52 : _GEN_10587;
  wire [13:0] _GEN_10589 = 14'h295d == index ? 14'h52 : _GEN_10588;
  wire [13:0] _GEN_10590 = 14'h295e == index ? 14'h52 : _GEN_10589;
  wire [13:0] _GEN_10591 = 14'h295f == index ? 14'h52 : _GEN_10590;
  wire [13:0] _GEN_10592 = 14'h2960 == index ? 14'h52 : _GEN_10591;
  wire [13:0] _GEN_10593 = 14'h2961 == index ? 14'h52 : _GEN_10592;
  wire [13:0] _GEN_10594 = 14'h2962 == index ? 14'h52 : _GEN_10593;
  wire [13:0] _GEN_10595 = 14'h2963 == index ? 14'h52 : _GEN_10594;
  wire [13:0] _GEN_10596 = 14'h2964 == index ? 14'h52 : _GEN_10595;
  wire [13:0] _GEN_10597 = 14'h2965 == index ? 14'h52 : _GEN_10596;
  wire [13:0] _GEN_10598 = 14'h2966 == index ? 14'h52 : _GEN_10597;
  wire [13:0] _GEN_10599 = 14'h2967 == index ? 14'h52 : _GEN_10598;
  wire [13:0] _GEN_10600 = 14'h2968 == index ? 14'h52 : _GEN_10599;
  wire [13:0] _GEN_10601 = 14'h2969 == index ? 14'h52 : _GEN_10600;
  wire [13:0] _GEN_10602 = 14'h296a == index ? 14'h52 : _GEN_10601;
  wire [13:0] _GEN_10603 = 14'h296b == index ? 14'h52 : _GEN_10602;
  wire [13:0] _GEN_10604 = 14'h296c == index ? 14'h52 : _GEN_10603;
  wire [13:0] _GEN_10605 = 14'h296d == index ? 14'h52 : _GEN_10604;
  wire [13:0] _GEN_10606 = 14'h296e == index ? 14'h52 : _GEN_10605;
  wire [13:0] _GEN_10607 = 14'h296f == index ? 14'h52 : _GEN_10606;
  wire [13:0] _GEN_10608 = 14'h2970 == index ? 14'h52 : _GEN_10607;
  wire [13:0] _GEN_10609 = 14'h2971 == index ? 14'h52 : _GEN_10608;
  wire [13:0] _GEN_10610 = 14'h2972 == index ? 14'h52 : _GEN_10609;
  wire [13:0] _GEN_10611 = 14'h2973 == index ? 14'h52 : _GEN_10610;
  wire [13:0] _GEN_10612 = 14'h2974 == index ? 14'h52 : _GEN_10611;
  wire [13:0] _GEN_10613 = 14'h2975 == index ? 14'h52 : _GEN_10612;
  wire [13:0] _GEN_10614 = 14'h2976 == index ? 14'h52 : _GEN_10613;
  wire [13:0] _GEN_10615 = 14'h2977 == index ? 14'h52 : _GEN_10614;
  wire [13:0] _GEN_10616 = 14'h2978 == index ? 14'h52 : _GEN_10615;
  wire [13:0] _GEN_10617 = 14'h2979 == index ? 14'h52 : _GEN_10616;
  wire [13:0] _GEN_10618 = 14'h297a == index ? 14'h52 : _GEN_10617;
  wire [13:0] _GEN_10619 = 14'h297b == index ? 14'h52 : _GEN_10618;
  wire [13:0] _GEN_10620 = 14'h297c == index ? 14'h52 : _GEN_10619;
  wire [13:0] _GEN_10621 = 14'h297d == index ? 14'h52 : _GEN_10620;
  wire [13:0] _GEN_10622 = 14'h297e == index ? 14'h52 : _GEN_10621;
  wire [13:0] _GEN_10623 = 14'h297f == index ? 14'h52 : _GEN_10622;
  wire [13:0] _GEN_10624 = 14'h2980 == index ? 14'h0 : _GEN_10623;
  wire [13:0] _GEN_10625 = 14'h2981 == index ? 14'h2980 : _GEN_10624;
  wire [13:0] _GEN_10626 = 14'h2982 == index ? 14'h1481 : _GEN_10625;
  wire [13:0] _GEN_10627 = 14'h2983 == index ? 14'hd82 : _GEN_10626;
  wire [13:0] _GEN_10628 = 14'h2984 == index ? 14'ha03 : _GEN_10627;
  wire [13:0] _GEN_10629 = 14'h2985 == index ? 14'h803 : _GEN_10628;
  wire [13:0] _GEN_10630 = 14'h2986 == index ? 14'h685 : _GEN_10629;
  wire [13:0] _GEN_10631 = 14'h2987 == index ? 14'h586 : _GEN_10630;
  wire [13:0] _GEN_10632 = 14'h2988 == index ? 14'h503 : _GEN_10631;
  wire [13:0] _GEN_10633 = 14'h2989 == index ? 14'h482 : _GEN_10632;
  wire [13:0] _GEN_10634 = 14'h298a == index ? 14'h403 : _GEN_10633;
  wire [13:0] _GEN_10635 = 14'h298b == index ? 14'h386 : _GEN_10634;
  wire [13:0] _GEN_10636 = 14'h298c == index ? 14'h30b : _GEN_10635;
  wire [13:0] _GEN_10637 = 14'h298d == index ? 14'h305 : _GEN_10636;
  wire [13:0] _GEN_10638 = 14'h298e == index ? 14'h28d : _GEN_10637;
  wire [13:0] _GEN_10639 = 14'h298f == index ? 14'h288 : _GEN_10638;
  wire [13:0] _GEN_10640 = 14'h2990 == index ? 14'h283 : _GEN_10639;
  wire [13:0] _GEN_10641 = 14'h2991 == index ? 14'h20f : _GEN_10640;
  wire [13:0] _GEN_10642 = 14'h2992 == index ? 14'h20b : _GEN_10641;
  wire [13:0] _GEN_10643 = 14'h2993 == index ? 14'h207 : _GEN_10642;
  wire [13:0] _GEN_10644 = 14'h2994 == index ? 14'h203 : _GEN_10643;
  wire [13:0] _GEN_10645 = 14'h2995 == index ? 14'h194 : _GEN_10644;
  wire [13:0] _GEN_10646 = 14'h2996 == index ? 14'h191 : _GEN_10645;
  wire [13:0] _GEN_10647 = 14'h2997 == index ? 14'h18e : _GEN_10646;
  wire [13:0] _GEN_10648 = 14'h2998 == index ? 14'h18b : _GEN_10647;
  wire [13:0] _GEN_10649 = 14'h2999 == index ? 14'h188 : _GEN_10648;
  wire [13:0] _GEN_10650 = 14'h299a == index ? 14'h185 : _GEN_10649;
  wire [13:0] _GEN_10651 = 14'h299b == index ? 14'h182 : _GEN_10650;
  wire [13:0] _GEN_10652 = 14'h299c == index ? 14'h11b : _GEN_10651;
  wire [13:0] _GEN_10653 = 14'h299d == index ? 14'h119 : _GEN_10652;
  wire [13:0] _GEN_10654 = 14'h299e == index ? 14'h117 : _GEN_10653;
  wire [13:0] _GEN_10655 = 14'h299f == index ? 14'h115 : _GEN_10654;
  wire [13:0] _GEN_10656 = 14'h29a0 == index ? 14'h113 : _GEN_10655;
  wire [13:0] _GEN_10657 = 14'h29a1 == index ? 14'h111 : _GEN_10656;
  wire [13:0] _GEN_10658 = 14'h29a2 == index ? 14'h10f : _GEN_10657;
  wire [13:0] _GEN_10659 = 14'h29a3 == index ? 14'h10d : _GEN_10658;
  wire [13:0] _GEN_10660 = 14'h29a4 == index ? 14'h10b : _GEN_10659;
  wire [13:0] _GEN_10661 = 14'h29a5 == index ? 14'h109 : _GEN_10660;
  wire [13:0] _GEN_10662 = 14'h29a6 == index ? 14'h107 : _GEN_10661;
  wire [13:0] _GEN_10663 = 14'h29a7 == index ? 14'h105 : _GEN_10662;
  wire [13:0] _GEN_10664 = 14'h29a8 == index ? 14'h103 : _GEN_10663;
  wire [13:0] _GEN_10665 = 14'h29a9 == index ? 14'h101 : _GEN_10664;
  wire [13:0] _GEN_10666 = 14'h29aa == index ? 14'ha9 : _GEN_10665;
  wire [13:0] _GEN_10667 = 14'h29ab == index ? 14'ha8 : _GEN_10666;
  wire [13:0] _GEN_10668 = 14'h29ac == index ? 14'ha7 : _GEN_10667;
  wire [13:0] _GEN_10669 = 14'h29ad == index ? 14'ha6 : _GEN_10668;
  wire [13:0] _GEN_10670 = 14'h29ae == index ? 14'ha5 : _GEN_10669;
  wire [13:0] _GEN_10671 = 14'h29af == index ? 14'ha4 : _GEN_10670;
  wire [13:0] _GEN_10672 = 14'h29b0 == index ? 14'ha3 : _GEN_10671;
  wire [13:0] _GEN_10673 = 14'h29b1 == index ? 14'ha2 : _GEN_10672;
  wire [13:0] _GEN_10674 = 14'h29b2 == index ? 14'ha1 : _GEN_10673;
  wire [13:0] _GEN_10675 = 14'h29b3 == index ? 14'ha0 : _GEN_10674;
  wire [13:0] _GEN_10676 = 14'h29b4 == index ? 14'h9f : _GEN_10675;
  wire [13:0] _GEN_10677 = 14'h29b5 == index ? 14'h9e : _GEN_10676;
  wire [13:0] _GEN_10678 = 14'h29b6 == index ? 14'h9d : _GEN_10677;
  wire [13:0] _GEN_10679 = 14'h29b7 == index ? 14'h9c : _GEN_10678;
  wire [13:0] _GEN_10680 = 14'h29b8 == index ? 14'h9b : _GEN_10679;
  wire [13:0] _GEN_10681 = 14'h29b9 == index ? 14'h9a : _GEN_10680;
  wire [13:0] _GEN_10682 = 14'h29ba == index ? 14'h99 : _GEN_10681;
  wire [13:0] _GEN_10683 = 14'h29bb == index ? 14'h98 : _GEN_10682;
  wire [13:0] _GEN_10684 = 14'h29bc == index ? 14'h97 : _GEN_10683;
  wire [13:0] _GEN_10685 = 14'h29bd == index ? 14'h96 : _GEN_10684;
  wire [13:0] _GEN_10686 = 14'h29be == index ? 14'h95 : _GEN_10685;
  wire [13:0] _GEN_10687 = 14'h29bf == index ? 14'h94 : _GEN_10686;
  wire [13:0] _GEN_10688 = 14'h29c0 == index ? 14'h93 : _GEN_10687;
  wire [13:0] _GEN_10689 = 14'h29c1 == index ? 14'h92 : _GEN_10688;
  wire [13:0] _GEN_10690 = 14'h29c2 == index ? 14'h91 : _GEN_10689;
  wire [13:0] _GEN_10691 = 14'h29c3 == index ? 14'h90 : _GEN_10690;
  wire [13:0] _GEN_10692 = 14'h29c4 == index ? 14'h8f : _GEN_10691;
  wire [13:0] _GEN_10693 = 14'h29c5 == index ? 14'h8e : _GEN_10692;
  wire [13:0] _GEN_10694 = 14'h29c6 == index ? 14'h8d : _GEN_10693;
  wire [13:0] _GEN_10695 = 14'h29c7 == index ? 14'h8c : _GEN_10694;
  wire [13:0] _GEN_10696 = 14'h29c8 == index ? 14'h8b : _GEN_10695;
  wire [13:0] _GEN_10697 = 14'h29c9 == index ? 14'h8a : _GEN_10696;
  wire [13:0] _GEN_10698 = 14'h29ca == index ? 14'h89 : _GEN_10697;
  wire [13:0] _GEN_10699 = 14'h29cb == index ? 14'h88 : _GEN_10698;
  wire [13:0] _GEN_10700 = 14'h29cc == index ? 14'h87 : _GEN_10699;
  wire [13:0] _GEN_10701 = 14'h29cd == index ? 14'h86 : _GEN_10700;
  wire [13:0] _GEN_10702 = 14'h29ce == index ? 14'h85 : _GEN_10701;
  wire [13:0] _GEN_10703 = 14'h29cf == index ? 14'h84 : _GEN_10702;
  wire [13:0] _GEN_10704 = 14'h29d0 == index ? 14'h83 : _GEN_10703;
  wire [13:0] _GEN_10705 = 14'h29d1 == index ? 14'h82 : _GEN_10704;
  wire [13:0] _GEN_10706 = 14'h29d2 == index ? 14'h81 : _GEN_10705;
  wire [13:0] _GEN_10707 = 14'h29d3 == index ? 14'h80 : _GEN_10706;
  wire [13:0] _GEN_10708 = 14'h29d4 == index ? 14'h53 : _GEN_10707;
  wire [13:0] _GEN_10709 = 14'h29d5 == index ? 14'h53 : _GEN_10708;
  wire [13:0] _GEN_10710 = 14'h29d6 == index ? 14'h53 : _GEN_10709;
  wire [13:0] _GEN_10711 = 14'h29d7 == index ? 14'h53 : _GEN_10710;
  wire [13:0] _GEN_10712 = 14'h29d8 == index ? 14'h53 : _GEN_10711;
  wire [13:0] _GEN_10713 = 14'h29d9 == index ? 14'h53 : _GEN_10712;
  wire [13:0] _GEN_10714 = 14'h29da == index ? 14'h53 : _GEN_10713;
  wire [13:0] _GEN_10715 = 14'h29db == index ? 14'h53 : _GEN_10714;
  wire [13:0] _GEN_10716 = 14'h29dc == index ? 14'h53 : _GEN_10715;
  wire [13:0] _GEN_10717 = 14'h29dd == index ? 14'h53 : _GEN_10716;
  wire [13:0] _GEN_10718 = 14'h29de == index ? 14'h53 : _GEN_10717;
  wire [13:0] _GEN_10719 = 14'h29df == index ? 14'h53 : _GEN_10718;
  wire [13:0] _GEN_10720 = 14'h29e0 == index ? 14'h53 : _GEN_10719;
  wire [13:0] _GEN_10721 = 14'h29e1 == index ? 14'h53 : _GEN_10720;
  wire [13:0] _GEN_10722 = 14'h29e2 == index ? 14'h53 : _GEN_10721;
  wire [13:0] _GEN_10723 = 14'h29e3 == index ? 14'h53 : _GEN_10722;
  wire [13:0] _GEN_10724 = 14'h29e4 == index ? 14'h53 : _GEN_10723;
  wire [13:0] _GEN_10725 = 14'h29e5 == index ? 14'h53 : _GEN_10724;
  wire [13:0] _GEN_10726 = 14'h29e6 == index ? 14'h53 : _GEN_10725;
  wire [13:0] _GEN_10727 = 14'h29e7 == index ? 14'h53 : _GEN_10726;
  wire [13:0] _GEN_10728 = 14'h29e8 == index ? 14'h53 : _GEN_10727;
  wire [13:0] _GEN_10729 = 14'h29e9 == index ? 14'h53 : _GEN_10728;
  wire [13:0] _GEN_10730 = 14'h29ea == index ? 14'h53 : _GEN_10729;
  wire [13:0] _GEN_10731 = 14'h29eb == index ? 14'h53 : _GEN_10730;
  wire [13:0] _GEN_10732 = 14'h29ec == index ? 14'h53 : _GEN_10731;
  wire [13:0] _GEN_10733 = 14'h29ed == index ? 14'h53 : _GEN_10732;
  wire [13:0] _GEN_10734 = 14'h29ee == index ? 14'h53 : _GEN_10733;
  wire [13:0] _GEN_10735 = 14'h29ef == index ? 14'h53 : _GEN_10734;
  wire [13:0] _GEN_10736 = 14'h29f0 == index ? 14'h53 : _GEN_10735;
  wire [13:0] _GEN_10737 = 14'h29f1 == index ? 14'h53 : _GEN_10736;
  wire [13:0] _GEN_10738 = 14'h29f2 == index ? 14'h53 : _GEN_10737;
  wire [13:0] _GEN_10739 = 14'h29f3 == index ? 14'h53 : _GEN_10738;
  wire [13:0] _GEN_10740 = 14'h29f4 == index ? 14'h53 : _GEN_10739;
  wire [13:0] _GEN_10741 = 14'h29f5 == index ? 14'h53 : _GEN_10740;
  wire [13:0] _GEN_10742 = 14'h29f6 == index ? 14'h53 : _GEN_10741;
  wire [13:0] _GEN_10743 = 14'h29f7 == index ? 14'h53 : _GEN_10742;
  wire [13:0] _GEN_10744 = 14'h29f8 == index ? 14'h53 : _GEN_10743;
  wire [13:0] _GEN_10745 = 14'h29f9 == index ? 14'h53 : _GEN_10744;
  wire [13:0] _GEN_10746 = 14'h29fa == index ? 14'h53 : _GEN_10745;
  wire [13:0] _GEN_10747 = 14'h29fb == index ? 14'h53 : _GEN_10746;
  wire [13:0] _GEN_10748 = 14'h29fc == index ? 14'h53 : _GEN_10747;
  wire [13:0] _GEN_10749 = 14'h29fd == index ? 14'h53 : _GEN_10748;
  wire [13:0] _GEN_10750 = 14'h29fe == index ? 14'h53 : _GEN_10749;
  wire [13:0] _GEN_10751 = 14'h29ff == index ? 14'h53 : _GEN_10750;
  wire [13:0] _GEN_10752 = 14'h2a00 == index ? 14'h0 : _GEN_10751;
  wire [13:0] _GEN_10753 = 14'h2a01 == index ? 14'h2a00 : _GEN_10752;
  wire [13:0] _GEN_10754 = 14'h2a02 == index ? 14'h1500 : _GEN_10753;
  wire [13:0] _GEN_10755 = 14'h2a03 == index ? 14'he00 : _GEN_10754;
  wire [13:0] _GEN_10756 = 14'h2a04 == index ? 14'ha80 : _GEN_10755;
  wire [13:0] _GEN_10757 = 14'h2a05 == index ? 14'h804 : _GEN_10756;
  wire [13:0] _GEN_10758 = 14'h2a06 == index ? 14'h700 : _GEN_10757;
  wire [13:0] _GEN_10759 = 14'h2a07 == index ? 14'h600 : _GEN_10758;
  wire [13:0] _GEN_10760 = 14'h2a08 == index ? 14'h504 : _GEN_10759;
  wire [13:0] _GEN_10761 = 14'h2a09 == index ? 14'h483 : _GEN_10760;
  wire [13:0] _GEN_10762 = 14'h2a0a == index ? 14'h404 : _GEN_10761;
  wire [13:0] _GEN_10763 = 14'h2a0b == index ? 14'h387 : _GEN_10762;
  wire [13:0] _GEN_10764 = 14'h2a0c == index ? 14'h380 : _GEN_10763;
  wire [13:0] _GEN_10765 = 14'h2a0d == index ? 14'h306 : _GEN_10764;
  wire [13:0] _GEN_10766 = 14'h2a0e == index ? 14'h300 : _GEN_10765;
  wire [13:0] _GEN_10767 = 14'h2a0f == index ? 14'h289 : _GEN_10766;
  wire [13:0] _GEN_10768 = 14'h2a10 == index ? 14'h284 : _GEN_10767;
  wire [13:0] _GEN_10769 = 14'h2a11 == index ? 14'h210 : _GEN_10768;
  wire [13:0] _GEN_10770 = 14'h2a12 == index ? 14'h20c : _GEN_10769;
  wire [13:0] _GEN_10771 = 14'h2a13 == index ? 14'h208 : _GEN_10770;
  wire [13:0] _GEN_10772 = 14'h2a14 == index ? 14'h204 : _GEN_10771;
  wire [13:0] _GEN_10773 = 14'h2a15 == index ? 14'h200 : _GEN_10772;
  wire [13:0] _GEN_10774 = 14'h2a16 == index ? 14'h192 : _GEN_10773;
  wire [13:0] _GEN_10775 = 14'h2a17 == index ? 14'h18f : _GEN_10774;
  wire [13:0] _GEN_10776 = 14'h2a18 == index ? 14'h18c : _GEN_10775;
  wire [13:0] _GEN_10777 = 14'h2a19 == index ? 14'h189 : _GEN_10776;
  wire [13:0] _GEN_10778 = 14'h2a1a == index ? 14'h186 : _GEN_10777;
  wire [13:0] _GEN_10779 = 14'h2a1b == index ? 14'h183 : _GEN_10778;
  wire [13:0] _GEN_10780 = 14'h2a1c == index ? 14'h180 : _GEN_10779;
  wire [13:0] _GEN_10781 = 14'h2a1d == index ? 14'h11a : _GEN_10780;
  wire [13:0] _GEN_10782 = 14'h2a1e == index ? 14'h118 : _GEN_10781;
  wire [13:0] _GEN_10783 = 14'h2a1f == index ? 14'h116 : _GEN_10782;
  wire [13:0] _GEN_10784 = 14'h2a20 == index ? 14'h114 : _GEN_10783;
  wire [13:0] _GEN_10785 = 14'h2a21 == index ? 14'h112 : _GEN_10784;
  wire [13:0] _GEN_10786 = 14'h2a22 == index ? 14'h110 : _GEN_10785;
  wire [13:0] _GEN_10787 = 14'h2a23 == index ? 14'h10e : _GEN_10786;
  wire [13:0] _GEN_10788 = 14'h2a24 == index ? 14'h10c : _GEN_10787;
  wire [13:0] _GEN_10789 = 14'h2a25 == index ? 14'h10a : _GEN_10788;
  wire [13:0] _GEN_10790 = 14'h2a26 == index ? 14'h108 : _GEN_10789;
  wire [13:0] _GEN_10791 = 14'h2a27 == index ? 14'h106 : _GEN_10790;
  wire [13:0] _GEN_10792 = 14'h2a28 == index ? 14'h104 : _GEN_10791;
  wire [13:0] _GEN_10793 = 14'h2a29 == index ? 14'h102 : _GEN_10792;
  wire [13:0] _GEN_10794 = 14'h2a2a == index ? 14'h100 : _GEN_10793;
  wire [13:0] _GEN_10795 = 14'h2a2b == index ? 14'ha9 : _GEN_10794;
  wire [13:0] _GEN_10796 = 14'h2a2c == index ? 14'ha8 : _GEN_10795;
  wire [13:0] _GEN_10797 = 14'h2a2d == index ? 14'ha7 : _GEN_10796;
  wire [13:0] _GEN_10798 = 14'h2a2e == index ? 14'ha6 : _GEN_10797;
  wire [13:0] _GEN_10799 = 14'h2a2f == index ? 14'ha5 : _GEN_10798;
  wire [13:0] _GEN_10800 = 14'h2a30 == index ? 14'ha4 : _GEN_10799;
  wire [13:0] _GEN_10801 = 14'h2a31 == index ? 14'ha3 : _GEN_10800;
  wire [13:0] _GEN_10802 = 14'h2a32 == index ? 14'ha2 : _GEN_10801;
  wire [13:0] _GEN_10803 = 14'h2a33 == index ? 14'ha1 : _GEN_10802;
  wire [13:0] _GEN_10804 = 14'h2a34 == index ? 14'ha0 : _GEN_10803;
  wire [13:0] _GEN_10805 = 14'h2a35 == index ? 14'h9f : _GEN_10804;
  wire [13:0] _GEN_10806 = 14'h2a36 == index ? 14'h9e : _GEN_10805;
  wire [13:0] _GEN_10807 = 14'h2a37 == index ? 14'h9d : _GEN_10806;
  wire [13:0] _GEN_10808 = 14'h2a38 == index ? 14'h9c : _GEN_10807;
  wire [13:0] _GEN_10809 = 14'h2a39 == index ? 14'h9b : _GEN_10808;
  wire [13:0] _GEN_10810 = 14'h2a3a == index ? 14'h9a : _GEN_10809;
  wire [13:0] _GEN_10811 = 14'h2a3b == index ? 14'h99 : _GEN_10810;
  wire [13:0] _GEN_10812 = 14'h2a3c == index ? 14'h98 : _GEN_10811;
  wire [13:0] _GEN_10813 = 14'h2a3d == index ? 14'h97 : _GEN_10812;
  wire [13:0] _GEN_10814 = 14'h2a3e == index ? 14'h96 : _GEN_10813;
  wire [13:0] _GEN_10815 = 14'h2a3f == index ? 14'h95 : _GEN_10814;
  wire [13:0] _GEN_10816 = 14'h2a40 == index ? 14'h94 : _GEN_10815;
  wire [13:0] _GEN_10817 = 14'h2a41 == index ? 14'h93 : _GEN_10816;
  wire [13:0] _GEN_10818 = 14'h2a42 == index ? 14'h92 : _GEN_10817;
  wire [13:0] _GEN_10819 = 14'h2a43 == index ? 14'h91 : _GEN_10818;
  wire [13:0] _GEN_10820 = 14'h2a44 == index ? 14'h90 : _GEN_10819;
  wire [13:0] _GEN_10821 = 14'h2a45 == index ? 14'h8f : _GEN_10820;
  wire [13:0] _GEN_10822 = 14'h2a46 == index ? 14'h8e : _GEN_10821;
  wire [13:0] _GEN_10823 = 14'h2a47 == index ? 14'h8d : _GEN_10822;
  wire [13:0] _GEN_10824 = 14'h2a48 == index ? 14'h8c : _GEN_10823;
  wire [13:0] _GEN_10825 = 14'h2a49 == index ? 14'h8b : _GEN_10824;
  wire [13:0] _GEN_10826 = 14'h2a4a == index ? 14'h8a : _GEN_10825;
  wire [13:0] _GEN_10827 = 14'h2a4b == index ? 14'h89 : _GEN_10826;
  wire [13:0] _GEN_10828 = 14'h2a4c == index ? 14'h88 : _GEN_10827;
  wire [13:0] _GEN_10829 = 14'h2a4d == index ? 14'h87 : _GEN_10828;
  wire [13:0] _GEN_10830 = 14'h2a4e == index ? 14'h86 : _GEN_10829;
  wire [13:0] _GEN_10831 = 14'h2a4f == index ? 14'h85 : _GEN_10830;
  wire [13:0] _GEN_10832 = 14'h2a50 == index ? 14'h84 : _GEN_10831;
  wire [13:0] _GEN_10833 = 14'h2a51 == index ? 14'h83 : _GEN_10832;
  wire [13:0] _GEN_10834 = 14'h2a52 == index ? 14'h82 : _GEN_10833;
  wire [13:0] _GEN_10835 = 14'h2a53 == index ? 14'h81 : _GEN_10834;
  wire [13:0] _GEN_10836 = 14'h2a54 == index ? 14'h80 : _GEN_10835;
  wire [13:0] _GEN_10837 = 14'h2a55 == index ? 14'h54 : _GEN_10836;
  wire [13:0] _GEN_10838 = 14'h2a56 == index ? 14'h54 : _GEN_10837;
  wire [13:0] _GEN_10839 = 14'h2a57 == index ? 14'h54 : _GEN_10838;
  wire [13:0] _GEN_10840 = 14'h2a58 == index ? 14'h54 : _GEN_10839;
  wire [13:0] _GEN_10841 = 14'h2a59 == index ? 14'h54 : _GEN_10840;
  wire [13:0] _GEN_10842 = 14'h2a5a == index ? 14'h54 : _GEN_10841;
  wire [13:0] _GEN_10843 = 14'h2a5b == index ? 14'h54 : _GEN_10842;
  wire [13:0] _GEN_10844 = 14'h2a5c == index ? 14'h54 : _GEN_10843;
  wire [13:0] _GEN_10845 = 14'h2a5d == index ? 14'h54 : _GEN_10844;
  wire [13:0] _GEN_10846 = 14'h2a5e == index ? 14'h54 : _GEN_10845;
  wire [13:0] _GEN_10847 = 14'h2a5f == index ? 14'h54 : _GEN_10846;
  wire [13:0] _GEN_10848 = 14'h2a60 == index ? 14'h54 : _GEN_10847;
  wire [13:0] _GEN_10849 = 14'h2a61 == index ? 14'h54 : _GEN_10848;
  wire [13:0] _GEN_10850 = 14'h2a62 == index ? 14'h54 : _GEN_10849;
  wire [13:0] _GEN_10851 = 14'h2a63 == index ? 14'h54 : _GEN_10850;
  wire [13:0] _GEN_10852 = 14'h2a64 == index ? 14'h54 : _GEN_10851;
  wire [13:0] _GEN_10853 = 14'h2a65 == index ? 14'h54 : _GEN_10852;
  wire [13:0] _GEN_10854 = 14'h2a66 == index ? 14'h54 : _GEN_10853;
  wire [13:0] _GEN_10855 = 14'h2a67 == index ? 14'h54 : _GEN_10854;
  wire [13:0] _GEN_10856 = 14'h2a68 == index ? 14'h54 : _GEN_10855;
  wire [13:0] _GEN_10857 = 14'h2a69 == index ? 14'h54 : _GEN_10856;
  wire [13:0] _GEN_10858 = 14'h2a6a == index ? 14'h54 : _GEN_10857;
  wire [13:0] _GEN_10859 = 14'h2a6b == index ? 14'h54 : _GEN_10858;
  wire [13:0] _GEN_10860 = 14'h2a6c == index ? 14'h54 : _GEN_10859;
  wire [13:0] _GEN_10861 = 14'h2a6d == index ? 14'h54 : _GEN_10860;
  wire [13:0] _GEN_10862 = 14'h2a6e == index ? 14'h54 : _GEN_10861;
  wire [13:0] _GEN_10863 = 14'h2a6f == index ? 14'h54 : _GEN_10862;
  wire [13:0] _GEN_10864 = 14'h2a70 == index ? 14'h54 : _GEN_10863;
  wire [13:0] _GEN_10865 = 14'h2a71 == index ? 14'h54 : _GEN_10864;
  wire [13:0] _GEN_10866 = 14'h2a72 == index ? 14'h54 : _GEN_10865;
  wire [13:0] _GEN_10867 = 14'h2a73 == index ? 14'h54 : _GEN_10866;
  wire [13:0] _GEN_10868 = 14'h2a74 == index ? 14'h54 : _GEN_10867;
  wire [13:0] _GEN_10869 = 14'h2a75 == index ? 14'h54 : _GEN_10868;
  wire [13:0] _GEN_10870 = 14'h2a76 == index ? 14'h54 : _GEN_10869;
  wire [13:0] _GEN_10871 = 14'h2a77 == index ? 14'h54 : _GEN_10870;
  wire [13:0] _GEN_10872 = 14'h2a78 == index ? 14'h54 : _GEN_10871;
  wire [13:0] _GEN_10873 = 14'h2a79 == index ? 14'h54 : _GEN_10872;
  wire [13:0] _GEN_10874 = 14'h2a7a == index ? 14'h54 : _GEN_10873;
  wire [13:0] _GEN_10875 = 14'h2a7b == index ? 14'h54 : _GEN_10874;
  wire [13:0] _GEN_10876 = 14'h2a7c == index ? 14'h54 : _GEN_10875;
  wire [13:0] _GEN_10877 = 14'h2a7d == index ? 14'h54 : _GEN_10876;
  wire [13:0] _GEN_10878 = 14'h2a7e == index ? 14'h54 : _GEN_10877;
  wire [13:0] _GEN_10879 = 14'h2a7f == index ? 14'h54 : _GEN_10878;
  wire [13:0] _GEN_10880 = 14'h2a80 == index ? 14'h0 : _GEN_10879;
  wire [13:0] _GEN_10881 = 14'h2a81 == index ? 14'h2a80 : _GEN_10880;
  wire [13:0] _GEN_10882 = 14'h2a82 == index ? 14'h1501 : _GEN_10881;
  wire [13:0] _GEN_10883 = 14'h2a83 == index ? 14'he01 : _GEN_10882;
  wire [13:0] _GEN_10884 = 14'h2a84 == index ? 14'ha81 : _GEN_10883;
  wire [13:0] _GEN_10885 = 14'h2a85 == index ? 14'h880 : _GEN_10884;
  wire [13:0] _GEN_10886 = 14'h2a86 == index ? 14'h701 : _GEN_10885;
  wire [13:0] _GEN_10887 = 14'h2a87 == index ? 14'h601 : _GEN_10886;
  wire [13:0] _GEN_10888 = 14'h2a88 == index ? 14'h505 : _GEN_10887;
  wire [13:0] _GEN_10889 = 14'h2a89 == index ? 14'h484 : _GEN_10888;
  wire [13:0] _GEN_10890 = 14'h2a8a == index ? 14'h405 : _GEN_10889;
  wire [13:0] _GEN_10891 = 14'h2a8b == index ? 14'h388 : _GEN_10890;
  wire [13:0] _GEN_10892 = 14'h2a8c == index ? 14'h381 : _GEN_10891;
  wire [13:0] _GEN_10893 = 14'h2a8d == index ? 14'h307 : _GEN_10892;
  wire [13:0] _GEN_10894 = 14'h2a8e == index ? 14'h301 : _GEN_10893;
  wire [13:0] _GEN_10895 = 14'h2a8f == index ? 14'h28a : _GEN_10894;
  wire [13:0] _GEN_10896 = 14'h2a90 == index ? 14'h285 : _GEN_10895;
  wire [13:0] _GEN_10897 = 14'h2a91 == index ? 14'h280 : _GEN_10896;
  wire [13:0] _GEN_10898 = 14'h2a92 == index ? 14'h20d : _GEN_10897;
  wire [13:0] _GEN_10899 = 14'h2a93 == index ? 14'h209 : _GEN_10898;
  wire [13:0] _GEN_10900 = 14'h2a94 == index ? 14'h205 : _GEN_10899;
  wire [13:0] _GEN_10901 = 14'h2a95 == index ? 14'h201 : _GEN_10900;
  wire [13:0] _GEN_10902 = 14'h2a96 == index ? 14'h193 : _GEN_10901;
  wire [13:0] _GEN_10903 = 14'h2a97 == index ? 14'h190 : _GEN_10902;
  wire [13:0] _GEN_10904 = 14'h2a98 == index ? 14'h18d : _GEN_10903;
  wire [13:0] _GEN_10905 = 14'h2a99 == index ? 14'h18a : _GEN_10904;
  wire [13:0] _GEN_10906 = 14'h2a9a == index ? 14'h187 : _GEN_10905;
  wire [13:0] _GEN_10907 = 14'h2a9b == index ? 14'h184 : _GEN_10906;
  wire [13:0] _GEN_10908 = 14'h2a9c == index ? 14'h181 : _GEN_10907;
  wire [13:0] _GEN_10909 = 14'h2a9d == index ? 14'h11b : _GEN_10908;
  wire [13:0] _GEN_10910 = 14'h2a9e == index ? 14'h119 : _GEN_10909;
  wire [13:0] _GEN_10911 = 14'h2a9f == index ? 14'h117 : _GEN_10910;
  wire [13:0] _GEN_10912 = 14'h2aa0 == index ? 14'h115 : _GEN_10911;
  wire [13:0] _GEN_10913 = 14'h2aa1 == index ? 14'h113 : _GEN_10912;
  wire [13:0] _GEN_10914 = 14'h2aa2 == index ? 14'h111 : _GEN_10913;
  wire [13:0] _GEN_10915 = 14'h2aa3 == index ? 14'h10f : _GEN_10914;
  wire [13:0] _GEN_10916 = 14'h2aa4 == index ? 14'h10d : _GEN_10915;
  wire [13:0] _GEN_10917 = 14'h2aa5 == index ? 14'h10b : _GEN_10916;
  wire [13:0] _GEN_10918 = 14'h2aa6 == index ? 14'h109 : _GEN_10917;
  wire [13:0] _GEN_10919 = 14'h2aa7 == index ? 14'h107 : _GEN_10918;
  wire [13:0] _GEN_10920 = 14'h2aa8 == index ? 14'h105 : _GEN_10919;
  wire [13:0] _GEN_10921 = 14'h2aa9 == index ? 14'h103 : _GEN_10920;
  wire [13:0] _GEN_10922 = 14'h2aaa == index ? 14'h101 : _GEN_10921;
  wire [13:0] _GEN_10923 = 14'h2aab == index ? 14'haa : _GEN_10922;
  wire [13:0] _GEN_10924 = 14'h2aac == index ? 14'ha9 : _GEN_10923;
  wire [13:0] _GEN_10925 = 14'h2aad == index ? 14'ha8 : _GEN_10924;
  wire [13:0] _GEN_10926 = 14'h2aae == index ? 14'ha7 : _GEN_10925;
  wire [13:0] _GEN_10927 = 14'h2aaf == index ? 14'ha6 : _GEN_10926;
  wire [13:0] _GEN_10928 = 14'h2ab0 == index ? 14'ha5 : _GEN_10927;
  wire [13:0] _GEN_10929 = 14'h2ab1 == index ? 14'ha4 : _GEN_10928;
  wire [13:0] _GEN_10930 = 14'h2ab2 == index ? 14'ha3 : _GEN_10929;
  wire [13:0] _GEN_10931 = 14'h2ab3 == index ? 14'ha2 : _GEN_10930;
  wire [13:0] _GEN_10932 = 14'h2ab4 == index ? 14'ha1 : _GEN_10931;
  wire [13:0] _GEN_10933 = 14'h2ab5 == index ? 14'ha0 : _GEN_10932;
  wire [13:0] _GEN_10934 = 14'h2ab6 == index ? 14'h9f : _GEN_10933;
  wire [13:0] _GEN_10935 = 14'h2ab7 == index ? 14'h9e : _GEN_10934;
  wire [13:0] _GEN_10936 = 14'h2ab8 == index ? 14'h9d : _GEN_10935;
  wire [13:0] _GEN_10937 = 14'h2ab9 == index ? 14'h9c : _GEN_10936;
  wire [13:0] _GEN_10938 = 14'h2aba == index ? 14'h9b : _GEN_10937;
  wire [13:0] _GEN_10939 = 14'h2abb == index ? 14'h9a : _GEN_10938;
  wire [13:0] _GEN_10940 = 14'h2abc == index ? 14'h99 : _GEN_10939;
  wire [13:0] _GEN_10941 = 14'h2abd == index ? 14'h98 : _GEN_10940;
  wire [13:0] _GEN_10942 = 14'h2abe == index ? 14'h97 : _GEN_10941;
  wire [13:0] _GEN_10943 = 14'h2abf == index ? 14'h96 : _GEN_10942;
  wire [13:0] _GEN_10944 = 14'h2ac0 == index ? 14'h95 : _GEN_10943;
  wire [13:0] _GEN_10945 = 14'h2ac1 == index ? 14'h94 : _GEN_10944;
  wire [13:0] _GEN_10946 = 14'h2ac2 == index ? 14'h93 : _GEN_10945;
  wire [13:0] _GEN_10947 = 14'h2ac3 == index ? 14'h92 : _GEN_10946;
  wire [13:0] _GEN_10948 = 14'h2ac4 == index ? 14'h91 : _GEN_10947;
  wire [13:0] _GEN_10949 = 14'h2ac5 == index ? 14'h90 : _GEN_10948;
  wire [13:0] _GEN_10950 = 14'h2ac6 == index ? 14'h8f : _GEN_10949;
  wire [13:0] _GEN_10951 = 14'h2ac7 == index ? 14'h8e : _GEN_10950;
  wire [13:0] _GEN_10952 = 14'h2ac8 == index ? 14'h8d : _GEN_10951;
  wire [13:0] _GEN_10953 = 14'h2ac9 == index ? 14'h8c : _GEN_10952;
  wire [13:0] _GEN_10954 = 14'h2aca == index ? 14'h8b : _GEN_10953;
  wire [13:0] _GEN_10955 = 14'h2acb == index ? 14'h8a : _GEN_10954;
  wire [13:0] _GEN_10956 = 14'h2acc == index ? 14'h89 : _GEN_10955;
  wire [13:0] _GEN_10957 = 14'h2acd == index ? 14'h88 : _GEN_10956;
  wire [13:0] _GEN_10958 = 14'h2ace == index ? 14'h87 : _GEN_10957;
  wire [13:0] _GEN_10959 = 14'h2acf == index ? 14'h86 : _GEN_10958;
  wire [13:0] _GEN_10960 = 14'h2ad0 == index ? 14'h85 : _GEN_10959;
  wire [13:0] _GEN_10961 = 14'h2ad1 == index ? 14'h84 : _GEN_10960;
  wire [13:0] _GEN_10962 = 14'h2ad2 == index ? 14'h83 : _GEN_10961;
  wire [13:0] _GEN_10963 = 14'h2ad3 == index ? 14'h82 : _GEN_10962;
  wire [13:0] _GEN_10964 = 14'h2ad4 == index ? 14'h81 : _GEN_10963;
  wire [13:0] _GEN_10965 = 14'h2ad5 == index ? 14'h80 : _GEN_10964;
  wire [13:0] _GEN_10966 = 14'h2ad6 == index ? 14'h55 : _GEN_10965;
  wire [13:0] _GEN_10967 = 14'h2ad7 == index ? 14'h55 : _GEN_10966;
  wire [13:0] _GEN_10968 = 14'h2ad8 == index ? 14'h55 : _GEN_10967;
  wire [13:0] _GEN_10969 = 14'h2ad9 == index ? 14'h55 : _GEN_10968;
  wire [13:0] _GEN_10970 = 14'h2ada == index ? 14'h55 : _GEN_10969;
  wire [13:0] _GEN_10971 = 14'h2adb == index ? 14'h55 : _GEN_10970;
  wire [13:0] _GEN_10972 = 14'h2adc == index ? 14'h55 : _GEN_10971;
  wire [13:0] _GEN_10973 = 14'h2add == index ? 14'h55 : _GEN_10972;
  wire [13:0] _GEN_10974 = 14'h2ade == index ? 14'h55 : _GEN_10973;
  wire [13:0] _GEN_10975 = 14'h2adf == index ? 14'h55 : _GEN_10974;
  wire [13:0] _GEN_10976 = 14'h2ae0 == index ? 14'h55 : _GEN_10975;
  wire [13:0] _GEN_10977 = 14'h2ae1 == index ? 14'h55 : _GEN_10976;
  wire [13:0] _GEN_10978 = 14'h2ae2 == index ? 14'h55 : _GEN_10977;
  wire [13:0] _GEN_10979 = 14'h2ae3 == index ? 14'h55 : _GEN_10978;
  wire [13:0] _GEN_10980 = 14'h2ae4 == index ? 14'h55 : _GEN_10979;
  wire [13:0] _GEN_10981 = 14'h2ae5 == index ? 14'h55 : _GEN_10980;
  wire [13:0] _GEN_10982 = 14'h2ae6 == index ? 14'h55 : _GEN_10981;
  wire [13:0] _GEN_10983 = 14'h2ae7 == index ? 14'h55 : _GEN_10982;
  wire [13:0] _GEN_10984 = 14'h2ae8 == index ? 14'h55 : _GEN_10983;
  wire [13:0] _GEN_10985 = 14'h2ae9 == index ? 14'h55 : _GEN_10984;
  wire [13:0] _GEN_10986 = 14'h2aea == index ? 14'h55 : _GEN_10985;
  wire [13:0] _GEN_10987 = 14'h2aeb == index ? 14'h55 : _GEN_10986;
  wire [13:0] _GEN_10988 = 14'h2aec == index ? 14'h55 : _GEN_10987;
  wire [13:0] _GEN_10989 = 14'h2aed == index ? 14'h55 : _GEN_10988;
  wire [13:0] _GEN_10990 = 14'h2aee == index ? 14'h55 : _GEN_10989;
  wire [13:0] _GEN_10991 = 14'h2aef == index ? 14'h55 : _GEN_10990;
  wire [13:0] _GEN_10992 = 14'h2af0 == index ? 14'h55 : _GEN_10991;
  wire [13:0] _GEN_10993 = 14'h2af1 == index ? 14'h55 : _GEN_10992;
  wire [13:0] _GEN_10994 = 14'h2af2 == index ? 14'h55 : _GEN_10993;
  wire [13:0] _GEN_10995 = 14'h2af3 == index ? 14'h55 : _GEN_10994;
  wire [13:0] _GEN_10996 = 14'h2af4 == index ? 14'h55 : _GEN_10995;
  wire [13:0] _GEN_10997 = 14'h2af5 == index ? 14'h55 : _GEN_10996;
  wire [13:0] _GEN_10998 = 14'h2af6 == index ? 14'h55 : _GEN_10997;
  wire [13:0] _GEN_10999 = 14'h2af7 == index ? 14'h55 : _GEN_10998;
  wire [13:0] _GEN_11000 = 14'h2af8 == index ? 14'h55 : _GEN_10999;
  wire [13:0] _GEN_11001 = 14'h2af9 == index ? 14'h55 : _GEN_11000;
  wire [13:0] _GEN_11002 = 14'h2afa == index ? 14'h55 : _GEN_11001;
  wire [13:0] _GEN_11003 = 14'h2afb == index ? 14'h55 : _GEN_11002;
  wire [13:0] _GEN_11004 = 14'h2afc == index ? 14'h55 : _GEN_11003;
  wire [13:0] _GEN_11005 = 14'h2afd == index ? 14'h55 : _GEN_11004;
  wire [13:0] _GEN_11006 = 14'h2afe == index ? 14'h55 : _GEN_11005;
  wire [13:0] _GEN_11007 = 14'h2aff == index ? 14'h55 : _GEN_11006;
  wire [13:0] _GEN_11008 = 14'h2b00 == index ? 14'h0 : _GEN_11007;
  wire [13:0] _GEN_11009 = 14'h2b01 == index ? 14'h2b00 : _GEN_11008;
  wire [13:0] _GEN_11010 = 14'h2b02 == index ? 14'h1580 : _GEN_11009;
  wire [13:0] _GEN_11011 = 14'h2b03 == index ? 14'he02 : _GEN_11010;
  wire [13:0] _GEN_11012 = 14'h2b04 == index ? 14'ha82 : _GEN_11011;
  wire [13:0] _GEN_11013 = 14'h2b05 == index ? 14'h881 : _GEN_11012;
  wire [13:0] _GEN_11014 = 14'h2b06 == index ? 14'h702 : _GEN_11013;
  wire [13:0] _GEN_11015 = 14'h2b07 == index ? 14'h602 : _GEN_11014;
  wire [13:0] _GEN_11016 = 14'h2b08 == index ? 14'h506 : _GEN_11015;
  wire [13:0] _GEN_11017 = 14'h2b09 == index ? 14'h485 : _GEN_11016;
  wire [13:0] _GEN_11018 = 14'h2b0a == index ? 14'h406 : _GEN_11017;
  wire [13:0] _GEN_11019 = 14'h2b0b == index ? 14'h389 : _GEN_11018;
  wire [13:0] _GEN_11020 = 14'h2b0c == index ? 14'h382 : _GEN_11019;
  wire [13:0] _GEN_11021 = 14'h2b0d == index ? 14'h308 : _GEN_11020;
  wire [13:0] _GEN_11022 = 14'h2b0e == index ? 14'h302 : _GEN_11021;
  wire [13:0] _GEN_11023 = 14'h2b0f == index ? 14'h28b : _GEN_11022;
  wire [13:0] _GEN_11024 = 14'h2b10 == index ? 14'h286 : _GEN_11023;
  wire [13:0] _GEN_11025 = 14'h2b11 == index ? 14'h281 : _GEN_11024;
  wire [13:0] _GEN_11026 = 14'h2b12 == index ? 14'h20e : _GEN_11025;
  wire [13:0] _GEN_11027 = 14'h2b13 == index ? 14'h20a : _GEN_11026;
  wire [13:0] _GEN_11028 = 14'h2b14 == index ? 14'h206 : _GEN_11027;
  wire [13:0] _GEN_11029 = 14'h2b15 == index ? 14'h202 : _GEN_11028;
  wire [13:0] _GEN_11030 = 14'h2b16 == index ? 14'h194 : _GEN_11029;
  wire [13:0] _GEN_11031 = 14'h2b17 == index ? 14'h191 : _GEN_11030;
  wire [13:0] _GEN_11032 = 14'h2b18 == index ? 14'h18e : _GEN_11031;
  wire [13:0] _GEN_11033 = 14'h2b19 == index ? 14'h18b : _GEN_11032;
  wire [13:0] _GEN_11034 = 14'h2b1a == index ? 14'h188 : _GEN_11033;
  wire [13:0] _GEN_11035 = 14'h2b1b == index ? 14'h185 : _GEN_11034;
  wire [13:0] _GEN_11036 = 14'h2b1c == index ? 14'h182 : _GEN_11035;
  wire [13:0] _GEN_11037 = 14'h2b1d == index ? 14'h11c : _GEN_11036;
  wire [13:0] _GEN_11038 = 14'h2b1e == index ? 14'h11a : _GEN_11037;
  wire [13:0] _GEN_11039 = 14'h2b1f == index ? 14'h118 : _GEN_11038;
  wire [13:0] _GEN_11040 = 14'h2b20 == index ? 14'h116 : _GEN_11039;
  wire [13:0] _GEN_11041 = 14'h2b21 == index ? 14'h114 : _GEN_11040;
  wire [13:0] _GEN_11042 = 14'h2b22 == index ? 14'h112 : _GEN_11041;
  wire [13:0] _GEN_11043 = 14'h2b23 == index ? 14'h110 : _GEN_11042;
  wire [13:0] _GEN_11044 = 14'h2b24 == index ? 14'h10e : _GEN_11043;
  wire [13:0] _GEN_11045 = 14'h2b25 == index ? 14'h10c : _GEN_11044;
  wire [13:0] _GEN_11046 = 14'h2b26 == index ? 14'h10a : _GEN_11045;
  wire [13:0] _GEN_11047 = 14'h2b27 == index ? 14'h108 : _GEN_11046;
  wire [13:0] _GEN_11048 = 14'h2b28 == index ? 14'h106 : _GEN_11047;
  wire [13:0] _GEN_11049 = 14'h2b29 == index ? 14'h104 : _GEN_11048;
  wire [13:0] _GEN_11050 = 14'h2b2a == index ? 14'h102 : _GEN_11049;
  wire [13:0] _GEN_11051 = 14'h2b2b == index ? 14'h100 : _GEN_11050;
  wire [13:0] _GEN_11052 = 14'h2b2c == index ? 14'haa : _GEN_11051;
  wire [13:0] _GEN_11053 = 14'h2b2d == index ? 14'ha9 : _GEN_11052;
  wire [13:0] _GEN_11054 = 14'h2b2e == index ? 14'ha8 : _GEN_11053;
  wire [13:0] _GEN_11055 = 14'h2b2f == index ? 14'ha7 : _GEN_11054;
  wire [13:0] _GEN_11056 = 14'h2b30 == index ? 14'ha6 : _GEN_11055;
  wire [13:0] _GEN_11057 = 14'h2b31 == index ? 14'ha5 : _GEN_11056;
  wire [13:0] _GEN_11058 = 14'h2b32 == index ? 14'ha4 : _GEN_11057;
  wire [13:0] _GEN_11059 = 14'h2b33 == index ? 14'ha3 : _GEN_11058;
  wire [13:0] _GEN_11060 = 14'h2b34 == index ? 14'ha2 : _GEN_11059;
  wire [13:0] _GEN_11061 = 14'h2b35 == index ? 14'ha1 : _GEN_11060;
  wire [13:0] _GEN_11062 = 14'h2b36 == index ? 14'ha0 : _GEN_11061;
  wire [13:0] _GEN_11063 = 14'h2b37 == index ? 14'h9f : _GEN_11062;
  wire [13:0] _GEN_11064 = 14'h2b38 == index ? 14'h9e : _GEN_11063;
  wire [13:0] _GEN_11065 = 14'h2b39 == index ? 14'h9d : _GEN_11064;
  wire [13:0] _GEN_11066 = 14'h2b3a == index ? 14'h9c : _GEN_11065;
  wire [13:0] _GEN_11067 = 14'h2b3b == index ? 14'h9b : _GEN_11066;
  wire [13:0] _GEN_11068 = 14'h2b3c == index ? 14'h9a : _GEN_11067;
  wire [13:0] _GEN_11069 = 14'h2b3d == index ? 14'h99 : _GEN_11068;
  wire [13:0] _GEN_11070 = 14'h2b3e == index ? 14'h98 : _GEN_11069;
  wire [13:0] _GEN_11071 = 14'h2b3f == index ? 14'h97 : _GEN_11070;
  wire [13:0] _GEN_11072 = 14'h2b40 == index ? 14'h96 : _GEN_11071;
  wire [13:0] _GEN_11073 = 14'h2b41 == index ? 14'h95 : _GEN_11072;
  wire [13:0] _GEN_11074 = 14'h2b42 == index ? 14'h94 : _GEN_11073;
  wire [13:0] _GEN_11075 = 14'h2b43 == index ? 14'h93 : _GEN_11074;
  wire [13:0] _GEN_11076 = 14'h2b44 == index ? 14'h92 : _GEN_11075;
  wire [13:0] _GEN_11077 = 14'h2b45 == index ? 14'h91 : _GEN_11076;
  wire [13:0] _GEN_11078 = 14'h2b46 == index ? 14'h90 : _GEN_11077;
  wire [13:0] _GEN_11079 = 14'h2b47 == index ? 14'h8f : _GEN_11078;
  wire [13:0] _GEN_11080 = 14'h2b48 == index ? 14'h8e : _GEN_11079;
  wire [13:0] _GEN_11081 = 14'h2b49 == index ? 14'h8d : _GEN_11080;
  wire [13:0] _GEN_11082 = 14'h2b4a == index ? 14'h8c : _GEN_11081;
  wire [13:0] _GEN_11083 = 14'h2b4b == index ? 14'h8b : _GEN_11082;
  wire [13:0] _GEN_11084 = 14'h2b4c == index ? 14'h8a : _GEN_11083;
  wire [13:0] _GEN_11085 = 14'h2b4d == index ? 14'h89 : _GEN_11084;
  wire [13:0] _GEN_11086 = 14'h2b4e == index ? 14'h88 : _GEN_11085;
  wire [13:0] _GEN_11087 = 14'h2b4f == index ? 14'h87 : _GEN_11086;
  wire [13:0] _GEN_11088 = 14'h2b50 == index ? 14'h86 : _GEN_11087;
  wire [13:0] _GEN_11089 = 14'h2b51 == index ? 14'h85 : _GEN_11088;
  wire [13:0] _GEN_11090 = 14'h2b52 == index ? 14'h84 : _GEN_11089;
  wire [13:0] _GEN_11091 = 14'h2b53 == index ? 14'h83 : _GEN_11090;
  wire [13:0] _GEN_11092 = 14'h2b54 == index ? 14'h82 : _GEN_11091;
  wire [13:0] _GEN_11093 = 14'h2b55 == index ? 14'h81 : _GEN_11092;
  wire [13:0] _GEN_11094 = 14'h2b56 == index ? 14'h80 : _GEN_11093;
  wire [13:0] _GEN_11095 = 14'h2b57 == index ? 14'h56 : _GEN_11094;
  wire [13:0] _GEN_11096 = 14'h2b58 == index ? 14'h56 : _GEN_11095;
  wire [13:0] _GEN_11097 = 14'h2b59 == index ? 14'h56 : _GEN_11096;
  wire [13:0] _GEN_11098 = 14'h2b5a == index ? 14'h56 : _GEN_11097;
  wire [13:0] _GEN_11099 = 14'h2b5b == index ? 14'h56 : _GEN_11098;
  wire [13:0] _GEN_11100 = 14'h2b5c == index ? 14'h56 : _GEN_11099;
  wire [13:0] _GEN_11101 = 14'h2b5d == index ? 14'h56 : _GEN_11100;
  wire [13:0] _GEN_11102 = 14'h2b5e == index ? 14'h56 : _GEN_11101;
  wire [13:0] _GEN_11103 = 14'h2b5f == index ? 14'h56 : _GEN_11102;
  wire [13:0] _GEN_11104 = 14'h2b60 == index ? 14'h56 : _GEN_11103;
  wire [13:0] _GEN_11105 = 14'h2b61 == index ? 14'h56 : _GEN_11104;
  wire [13:0] _GEN_11106 = 14'h2b62 == index ? 14'h56 : _GEN_11105;
  wire [13:0] _GEN_11107 = 14'h2b63 == index ? 14'h56 : _GEN_11106;
  wire [13:0] _GEN_11108 = 14'h2b64 == index ? 14'h56 : _GEN_11107;
  wire [13:0] _GEN_11109 = 14'h2b65 == index ? 14'h56 : _GEN_11108;
  wire [13:0] _GEN_11110 = 14'h2b66 == index ? 14'h56 : _GEN_11109;
  wire [13:0] _GEN_11111 = 14'h2b67 == index ? 14'h56 : _GEN_11110;
  wire [13:0] _GEN_11112 = 14'h2b68 == index ? 14'h56 : _GEN_11111;
  wire [13:0] _GEN_11113 = 14'h2b69 == index ? 14'h56 : _GEN_11112;
  wire [13:0] _GEN_11114 = 14'h2b6a == index ? 14'h56 : _GEN_11113;
  wire [13:0] _GEN_11115 = 14'h2b6b == index ? 14'h56 : _GEN_11114;
  wire [13:0] _GEN_11116 = 14'h2b6c == index ? 14'h56 : _GEN_11115;
  wire [13:0] _GEN_11117 = 14'h2b6d == index ? 14'h56 : _GEN_11116;
  wire [13:0] _GEN_11118 = 14'h2b6e == index ? 14'h56 : _GEN_11117;
  wire [13:0] _GEN_11119 = 14'h2b6f == index ? 14'h56 : _GEN_11118;
  wire [13:0] _GEN_11120 = 14'h2b70 == index ? 14'h56 : _GEN_11119;
  wire [13:0] _GEN_11121 = 14'h2b71 == index ? 14'h56 : _GEN_11120;
  wire [13:0] _GEN_11122 = 14'h2b72 == index ? 14'h56 : _GEN_11121;
  wire [13:0] _GEN_11123 = 14'h2b73 == index ? 14'h56 : _GEN_11122;
  wire [13:0] _GEN_11124 = 14'h2b74 == index ? 14'h56 : _GEN_11123;
  wire [13:0] _GEN_11125 = 14'h2b75 == index ? 14'h56 : _GEN_11124;
  wire [13:0] _GEN_11126 = 14'h2b76 == index ? 14'h56 : _GEN_11125;
  wire [13:0] _GEN_11127 = 14'h2b77 == index ? 14'h56 : _GEN_11126;
  wire [13:0] _GEN_11128 = 14'h2b78 == index ? 14'h56 : _GEN_11127;
  wire [13:0] _GEN_11129 = 14'h2b79 == index ? 14'h56 : _GEN_11128;
  wire [13:0] _GEN_11130 = 14'h2b7a == index ? 14'h56 : _GEN_11129;
  wire [13:0] _GEN_11131 = 14'h2b7b == index ? 14'h56 : _GEN_11130;
  wire [13:0] _GEN_11132 = 14'h2b7c == index ? 14'h56 : _GEN_11131;
  wire [13:0] _GEN_11133 = 14'h2b7d == index ? 14'h56 : _GEN_11132;
  wire [13:0] _GEN_11134 = 14'h2b7e == index ? 14'h56 : _GEN_11133;
  wire [13:0] _GEN_11135 = 14'h2b7f == index ? 14'h56 : _GEN_11134;
  wire [13:0] _GEN_11136 = 14'h2b80 == index ? 14'h0 : _GEN_11135;
  wire [13:0] _GEN_11137 = 14'h2b81 == index ? 14'h2b80 : _GEN_11136;
  wire [13:0] _GEN_11138 = 14'h2b82 == index ? 14'h1581 : _GEN_11137;
  wire [13:0] _GEN_11139 = 14'h2b83 == index ? 14'he80 : _GEN_11138;
  wire [13:0] _GEN_11140 = 14'h2b84 == index ? 14'ha83 : _GEN_11139;
  wire [13:0] _GEN_11141 = 14'h2b85 == index ? 14'h882 : _GEN_11140;
  wire [13:0] _GEN_11142 = 14'h2b86 == index ? 14'h703 : _GEN_11141;
  wire [13:0] _GEN_11143 = 14'h2b87 == index ? 14'h603 : _GEN_11142;
  wire [13:0] _GEN_11144 = 14'h2b88 == index ? 14'h507 : _GEN_11143;
  wire [13:0] _GEN_11145 = 14'h2b89 == index ? 14'h486 : _GEN_11144;
  wire [13:0] _GEN_11146 = 14'h2b8a == index ? 14'h407 : _GEN_11145;
  wire [13:0] _GEN_11147 = 14'h2b8b == index ? 14'h38a : _GEN_11146;
  wire [13:0] _GEN_11148 = 14'h2b8c == index ? 14'h383 : _GEN_11147;
  wire [13:0] _GEN_11149 = 14'h2b8d == index ? 14'h309 : _GEN_11148;
  wire [13:0] _GEN_11150 = 14'h2b8e == index ? 14'h303 : _GEN_11149;
  wire [13:0] _GEN_11151 = 14'h2b8f == index ? 14'h28c : _GEN_11150;
  wire [13:0] _GEN_11152 = 14'h2b90 == index ? 14'h287 : _GEN_11151;
  wire [13:0] _GEN_11153 = 14'h2b91 == index ? 14'h282 : _GEN_11152;
  wire [13:0] _GEN_11154 = 14'h2b92 == index ? 14'h20f : _GEN_11153;
  wire [13:0] _GEN_11155 = 14'h2b93 == index ? 14'h20b : _GEN_11154;
  wire [13:0] _GEN_11156 = 14'h2b94 == index ? 14'h207 : _GEN_11155;
  wire [13:0] _GEN_11157 = 14'h2b95 == index ? 14'h203 : _GEN_11156;
  wire [13:0] _GEN_11158 = 14'h2b96 == index ? 14'h195 : _GEN_11157;
  wire [13:0] _GEN_11159 = 14'h2b97 == index ? 14'h192 : _GEN_11158;
  wire [13:0] _GEN_11160 = 14'h2b98 == index ? 14'h18f : _GEN_11159;
  wire [13:0] _GEN_11161 = 14'h2b99 == index ? 14'h18c : _GEN_11160;
  wire [13:0] _GEN_11162 = 14'h2b9a == index ? 14'h189 : _GEN_11161;
  wire [13:0] _GEN_11163 = 14'h2b9b == index ? 14'h186 : _GEN_11162;
  wire [13:0] _GEN_11164 = 14'h2b9c == index ? 14'h183 : _GEN_11163;
  wire [13:0] _GEN_11165 = 14'h2b9d == index ? 14'h180 : _GEN_11164;
  wire [13:0] _GEN_11166 = 14'h2b9e == index ? 14'h11b : _GEN_11165;
  wire [13:0] _GEN_11167 = 14'h2b9f == index ? 14'h119 : _GEN_11166;
  wire [13:0] _GEN_11168 = 14'h2ba0 == index ? 14'h117 : _GEN_11167;
  wire [13:0] _GEN_11169 = 14'h2ba1 == index ? 14'h115 : _GEN_11168;
  wire [13:0] _GEN_11170 = 14'h2ba2 == index ? 14'h113 : _GEN_11169;
  wire [13:0] _GEN_11171 = 14'h2ba3 == index ? 14'h111 : _GEN_11170;
  wire [13:0] _GEN_11172 = 14'h2ba4 == index ? 14'h10f : _GEN_11171;
  wire [13:0] _GEN_11173 = 14'h2ba5 == index ? 14'h10d : _GEN_11172;
  wire [13:0] _GEN_11174 = 14'h2ba6 == index ? 14'h10b : _GEN_11173;
  wire [13:0] _GEN_11175 = 14'h2ba7 == index ? 14'h109 : _GEN_11174;
  wire [13:0] _GEN_11176 = 14'h2ba8 == index ? 14'h107 : _GEN_11175;
  wire [13:0] _GEN_11177 = 14'h2ba9 == index ? 14'h105 : _GEN_11176;
  wire [13:0] _GEN_11178 = 14'h2baa == index ? 14'h103 : _GEN_11177;
  wire [13:0] _GEN_11179 = 14'h2bab == index ? 14'h101 : _GEN_11178;
  wire [13:0] _GEN_11180 = 14'h2bac == index ? 14'hab : _GEN_11179;
  wire [13:0] _GEN_11181 = 14'h2bad == index ? 14'haa : _GEN_11180;
  wire [13:0] _GEN_11182 = 14'h2bae == index ? 14'ha9 : _GEN_11181;
  wire [13:0] _GEN_11183 = 14'h2baf == index ? 14'ha8 : _GEN_11182;
  wire [13:0] _GEN_11184 = 14'h2bb0 == index ? 14'ha7 : _GEN_11183;
  wire [13:0] _GEN_11185 = 14'h2bb1 == index ? 14'ha6 : _GEN_11184;
  wire [13:0] _GEN_11186 = 14'h2bb2 == index ? 14'ha5 : _GEN_11185;
  wire [13:0] _GEN_11187 = 14'h2bb3 == index ? 14'ha4 : _GEN_11186;
  wire [13:0] _GEN_11188 = 14'h2bb4 == index ? 14'ha3 : _GEN_11187;
  wire [13:0] _GEN_11189 = 14'h2bb5 == index ? 14'ha2 : _GEN_11188;
  wire [13:0] _GEN_11190 = 14'h2bb6 == index ? 14'ha1 : _GEN_11189;
  wire [13:0] _GEN_11191 = 14'h2bb7 == index ? 14'ha0 : _GEN_11190;
  wire [13:0] _GEN_11192 = 14'h2bb8 == index ? 14'h9f : _GEN_11191;
  wire [13:0] _GEN_11193 = 14'h2bb9 == index ? 14'h9e : _GEN_11192;
  wire [13:0] _GEN_11194 = 14'h2bba == index ? 14'h9d : _GEN_11193;
  wire [13:0] _GEN_11195 = 14'h2bbb == index ? 14'h9c : _GEN_11194;
  wire [13:0] _GEN_11196 = 14'h2bbc == index ? 14'h9b : _GEN_11195;
  wire [13:0] _GEN_11197 = 14'h2bbd == index ? 14'h9a : _GEN_11196;
  wire [13:0] _GEN_11198 = 14'h2bbe == index ? 14'h99 : _GEN_11197;
  wire [13:0] _GEN_11199 = 14'h2bbf == index ? 14'h98 : _GEN_11198;
  wire [13:0] _GEN_11200 = 14'h2bc0 == index ? 14'h97 : _GEN_11199;
  wire [13:0] _GEN_11201 = 14'h2bc1 == index ? 14'h96 : _GEN_11200;
  wire [13:0] _GEN_11202 = 14'h2bc2 == index ? 14'h95 : _GEN_11201;
  wire [13:0] _GEN_11203 = 14'h2bc3 == index ? 14'h94 : _GEN_11202;
  wire [13:0] _GEN_11204 = 14'h2bc4 == index ? 14'h93 : _GEN_11203;
  wire [13:0] _GEN_11205 = 14'h2bc5 == index ? 14'h92 : _GEN_11204;
  wire [13:0] _GEN_11206 = 14'h2bc6 == index ? 14'h91 : _GEN_11205;
  wire [13:0] _GEN_11207 = 14'h2bc7 == index ? 14'h90 : _GEN_11206;
  wire [13:0] _GEN_11208 = 14'h2bc8 == index ? 14'h8f : _GEN_11207;
  wire [13:0] _GEN_11209 = 14'h2bc9 == index ? 14'h8e : _GEN_11208;
  wire [13:0] _GEN_11210 = 14'h2bca == index ? 14'h8d : _GEN_11209;
  wire [13:0] _GEN_11211 = 14'h2bcb == index ? 14'h8c : _GEN_11210;
  wire [13:0] _GEN_11212 = 14'h2bcc == index ? 14'h8b : _GEN_11211;
  wire [13:0] _GEN_11213 = 14'h2bcd == index ? 14'h8a : _GEN_11212;
  wire [13:0] _GEN_11214 = 14'h2bce == index ? 14'h89 : _GEN_11213;
  wire [13:0] _GEN_11215 = 14'h2bcf == index ? 14'h88 : _GEN_11214;
  wire [13:0] _GEN_11216 = 14'h2bd0 == index ? 14'h87 : _GEN_11215;
  wire [13:0] _GEN_11217 = 14'h2bd1 == index ? 14'h86 : _GEN_11216;
  wire [13:0] _GEN_11218 = 14'h2bd2 == index ? 14'h85 : _GEN_11217;
  wire [13:0] _GEN_11219 = 14'h2bd3 == index ? 14'h84 : _GEN_11218;
  wire [13:0] _GEN_11220 = 14'h2bd4 == index ? 14'h83 : _GEN_11219;
  wire [13:0] _GEN_11221 = 14'h2bd5 == index ? 14'h82 : _GEN_11220;
  wire [13:0] _GEN_11222 = 14'h2bd6 == index ? 14'h81 : _GEN_11221;
  wire [13:0] _GEN_11223 = 14'h2bd7 == index ? 14'h80 : _GEN_11222;
  wire [13:0] _GEN_11224 = 14'h2bd8 == index ? 14'h57 : _GEN_11223;
  wire [13:0] _GEN_11225 = 14'h2bd9 == index ? 14'h57 : _GEN_11224;
  wire [13:0] _GEN_11226 = 14'h2bda == index ? 14'h57 : _GEN_11225;
  wire [13:0] _GEN_11227 = 14'h2bdb == index ? 14'h57 : _GEN_11226;
  wire [13:0] _GEN_11228 = 14'h2bdc == index ? 14'h57 : _GEN_11227;
  wire [13:0] _GEN_11229 = 14'h2bdd == index ? 14'h57 : _GEN_11228;
  wire [13:0] _GEN_11230 = 14'h2bde == index ? 14'h57 : _GEN_11229;
  wire [13:0] _GEN_11231 = 14'h2bdf == index ? 14'h57 : _GEN_11230;
  wire [13:0] _GEN_11232 = 14'h2be0 == index ? 14'h57 : _GEN_11231;
  wire [13:0] _GEN_11233 = 14'h2be1 == index ? 14'h57 : _GEN_11232;
  wire [13:0] _GEN_11234 = 14'h2be2 == index ? 14'h57 : _GEN_11233;
  wire [13:0] _GEN_11235 = 14'h2be3 == index ? 14'h57 : _GEN_11234;
  wire [13:0] _GEN_11236 = 14'h2be4 == index ? 14'h57 : _GEN_11235;
  wire [13:0] _GEN_11237 = 14'h2be5 == index ? 14'h57 : _GEN_11236;
  wire [13:0] _GEN_11238 = 14'h2be6 == index ? 14'h57 : _GEN_11237;
  wire [13:0] _GEN_11239 = 14'h2be7 == index ? 14'h57 : _GEN_11238;
  wire [13:0] _GEN_11240 = 14'h2be8 == index ? 14'h57 : _GEN_11239;
  wire [13:0] _GEN_11241 = 14'h2be9 == index ? 14'h57 : _GEN_11240;
  wire [13:0] _GEN_11242 = 14'h2bea == index ? 14'h57 : _GEN_11241;
  wire [13:0] _GEN_11243 = 14'h2beb == index ? 14'h57 : _GEN_11242;
  wire [13:0] _GEN_11244 = 14'h2bec == index ? 14'h57 : _GEN_11243;
  wire [13:0] _GEN_11245 = 14'h2bed == index ? 14'h57 : _GEN_11244;
  wire [13:0] _GEN_11246 = 14'h2bee == index ? 14'h57 : _GEN_11245;
  wire [13:0] _GEN_11247 = 14'h2bef == index ? 14'h57 : _GEN_11246;
  wire [13:0] _GEN_11248 = 14'h2bf0 == index ? 14'h57 : _GEN_11247;
  wire [13:0] _GEN_11249 = 14'h2bf1 == index ? 14'h57 : _GEN_11248;
  wire [13:0] _GEN_11250 = 14'h2bf2 == index ? 14'h57 : _GEN_11249;
  wire [13:0] _GEN_11251 = 14'h2bf3 == index ? 14'h57 : _GEN_11250;
  wire [13:0] _GEN_11252 = 14'h2bf4 == index ? 14'h57 : _GEN_11251;
  wire [13:0] _GEN_11253 = 14'h2bf5 == index ? 14'h57 : _GEN_11252;
  wire [13:0] _GEN_11254 = 14'h2bf6 == index ? 14'h57 : _GEN_11253;
  wire [13:0] _GEN_11255 = 14'h2bf7 == index ? 14'h57 : _GEN_11254;
  wire [13:0] _GEN_11256 = 14'h2bf8 == index ? 14'h57 : _GEN_11255;
  wire [13:0] _GEN_11257 = 14'h2bf9 == index ? 14'h57 : _GEN_11256;
  wire [13:0] _GEN_11258 = 14'h2bfa == index ? 14'h57 : _GEN_11257;
  wire [13:0] _GEN_11259 = 14'h2bfb == index ? 14'h57 : _GEN_11258;
  wire [13:0] _GEN_11260 = 14'h2bfc == index ? 14'h57 : _GEN_11259;
  wire [13:0] _GEN_11261 = 14'h2bfd == index ? 14'h57 : _GEN_11260;
  wire [13:0] _GEN_11262 = 14'h2bfe == index ? 14'h57 : _GEN_11261;
  wire [13:0] _GEN_11263 = 14'h2bff == index ? 14'h57 : _GEN_11262;
  wire [13:0] _GEN_11264 = 14'h2c00 == index ? 14'h0 : _GEN_11263;
  wire [13:0] _GEN_11265 = 14'h2c01 == index ? 14'h2c00 : _GEN_11264;
  wire [13:0] _GEN_11266 = 14'h2c02 == index ? 14'h1600 : _GEN_11265;
  wire [13:0] _GEN_11267 = 14'h2c03 == index ? 14'he81 : _GEN_11266;
  wire [13:0] _GEN_11268 = 14'h2c04 == index ? 14'hb00 : _GEN_11267;
  wire [13:0] _GEN_11269 = 14'h2c05 == index ? 14'h883 : _GEN_11268;
  wire [13:0] _GEN_11270 = 14'h2c06 == index ? 14'h704 : _GEN_11269;
  wire [13:0] _GEN_11271 = 14'h2c07 == index ? 14'h604 : _GEN_11270;
  wire [13:0] _GEN_11272 = 14'h2c08 == index ? 14'h580 : _GEN_11271;
  wire [13:0] _GEN_11273 = 14'h2c09 == index ? 14'h487 : _GEN_11272;
  wire [13:0] _GEN_11274 = 14'h2c0a == index ? 14'h408 : _GEN_11273;
  wire [13:0] _GEN_11275 = 14'h2c0b == index ? 14'h400 : _GEN_11274;
  wire [13:0] _GEN_11276 = 14'h2c0c == index ? 14'h384 : _GEN_11275;
  wire [13:0] _GEN_11277 = 14'h2c0d == index ? 14'h30a : _GEN_11276;
  wire [13:0] _GEN_11278 = 14'h2c0e == index ? 14'h304 : _GEN_11277;
  wire [13:0] _GEN_11279 = 14'h2c0f == index ? 14'h28d : _GEN_11278;
  wire [13:0] _GEN_11280 = 14'h2c10 == index ? 14'h288 : _GEN_11279;
  wire [13:0] _GEN_11281 = 14'h2c11 == index ? 14'h283 : _GEN_11280;
  wire [13:0] _GEN_11282 = 14'h2c12 == index ? 14'h210 : _GEN_11281;
  wire [13:0] _GEN_11283 = 14'h2c13 == index ? 14'h20c : _GEN_11282;
  wire [13:0] _GEN_11284 = 14'h2c14 == index ? 14'h208 : _GEN_11283;
  wire [13:0] _GEN_11285 = 14'h2c15 == index ? 14'h204 : _GEN_11284;
  wire [13:0] _GEN_11286 = 14'h2c16 == index ? 14'h200 : _GEN_11285;
  wire [13:0] _GEN_11287 = 14'h2c17 == index ? 14'h193 : _GEN_11286;
  wire [13:0] _GEN_11288 = 14'h2c18 == index ? 14'h190 : _GEN_11287;
  wire [13:0] _GEN_11289 = 14'h2c19 == index ? 14'h18d : _GEN_11288;
  wire [13:0] _GEN_11290 = 14'h2c1a == index ? 14'h18a : _GEN_11289;
  wire [13:0] _GEN_11291 = 14'h2c1b == index ? 14'h187 : _GEN_11290;
  wire [13:0] _GEN_11292 = 14'h2c1c == index ? 14'h184 : _GEN_11291;
  wire [13:0] _GEN_11293 = 14'h2c1d == index ? 14'h181 : _GEN_11292;
  wire [13:0] _GEN_11294 = 14'h2c1e == index ? 14'h11c : _GEN_11293;
  wire [13:0] _GEN_11295 = 14'h2c1f == index ? 14'h11a : _GEN_11294;
  wire [13:0] _GEN_11296 = 14'h2c20 == index ? 14'h118 : _GEN_11295;
  wire [13:0] _GEN_11297 = 14'h2c21 == index ? 14'h116 : _GEN_11296;
  wire [13:0] _GEN_11298 = 14'h2c22 == index ? 14'h114 : _GEN_11297;
  wire [13:0] _GEN_11299 = 14'h2c23 == index ? 14'h112 : _GEN_11298;
  wire [13:0] _GEN_11300 = 14'h2c24 == index ? 14'h110 : _GEN_11299;
  wire [13:0] _GEN_11301 = 14'h2c25 == index ? 14'h10e : _GEN_11300;
  wire [13:0] _GEN_11302 = 14'h2c26 == index ? 14'h10c : _GEN_11301;
  wire [13:0] _GEN_11303 = 14'h2c27 == index ? 14'h10a : _GEN_11302;
  wire [13:0] _GEN_11304 = 14'h2c28 == index ? 14'h108 : _GEN_11303;
  wire [13:0] _GEN_11305 = 14'h2c29 == index ? 14'h106 : _GEN_11304;
  wire [13:0] _GEN_11306 = 14'h2c2a == index ? 14'h104 : _GEN_11305;
  wire [13:0] _GEN_11307 = 14'h2c2b == index ? 14'h102 : _GEN_11306;
  wire [13:0] _GEN_11308 = 14'h2c2c == index ? 14'h100 : _GEN_11307;
  wire [13:0] _GEN_11309 = 14'h2c2d == index ? 14'hab : _GEN_11308;
  wire [13:0] _GEN_11310 = 14'h2c2e == index ? 14'haa : _GEN_11309;
  wire [13:0] _GEN_11311 = 14'h2c2f == index ? 14'ha9 : _GEN_11310;
  wire [13:0] _GEN_11312 = 14'h2c30 == index ? 14'ha8 : _GEN_11311;
  wire [13:0] _GEN_11313 = 14'h2c31 == index ? 14'ha7 : _GEN_11312;
  wire [13:0] _GEN_11314 = 14'h2c32 == index ? 14'ha6 : _GEN_11313;
  wire [13:0] _GEN_11315 = 14'h2c33 == index ? 14'ha5 : _GEN_11314;
  wire [13:0] _GEN_11316 = 14'h2c34 == index ? 14'ha4 : _GEN_11315;
  wire [13:0] _GEN_11317 = 14'h2c35 == index ? 14'ha3 : _GEN_11316;
  wire [13:0] _GEN_11318 = 14'h2c36 == index ? 14'ha2 : _GEN_11317;
  wire [13:0] _GEN_11319 = 14'h2c37 == index ? 14'ha1 : _GEN_11318;
  wire [13:0] _GEN_11320 = 14'h2c38 == index ? 14'ha0 : _GEN_11319;
  wire [13:0] _GEN_11321 = 14'h2c39 == index ? 14'h9f : _GEN_11320;
  wire [13:0] _GEN_11322 = 14'h2c3a == index ? 14'h9e : _GEN_11321;
  wire [13:0] _GEN_11323 = 14'h2c3b == index ? 14'h9d : _GEN_11322;
  wire [13:0] _GEN_11324 = 14'h2c3c == index ? 14'h9c : _GEN_11323;
  wire [13:0] _GEN_11325 = 14'h2c3d == index ? 14'h9b : _GEN_11324;
  wire [13:0] _GEN_11326 = 14'h2c3e == index ? 14'h9a : _GEN_11325;
  wire [13:0] _GEN_11327 = 14'h2c3f == index ? 14'h99 : _GEN_11326;
  wire [13:0] _GEN_11328 = 14'h2c40 == index ? 14'h98 : _GEN_11327;
  wire [13:0] _GEN_11329 = 14'h2c41 == index ? 14'h97 : _GEN_11328;
  wire [13:0] _GEN_11330 = 14'h2c42 == index ? 14'h96 : _GEN_11329;
  wire [13:0] _GEN_11331 = 14'h2c43 == index ? 14'h95 : _GEN_11330;
  wire [13:0] _GEN_11332 = 14'h2c44 == index ? 14'h94 : _GEN_11331;
  wire [13:0] _GEN_11333 = 14'h2c45 == index ? 14'h93 : _GEN_11332;
  wire [13:0] _GEN_11334 = 14'h2c46 == index ? 14'h92 : _GEN_11333;
  wire [13:0] _GEN_11335 = 14'h2c47 == index ? 14'h91 : _GEN_11334;
  wire [13:0] _GEN_11336 = 14'h2c48 == index ? 14'h90 : _GEN_11335;
  wire [13:0] _GEN_11337 = 14'h2c49 == index ? 14'h8f : _GEN_11336;
  wire [13:0] _GEN_11338 = 14'h2c4a == index ? 14'h8e : _GEN_11337;
  wire [13:0] _GEN_11339 = 14'h2c4b == index ? 14'h8d : _GEN_11338;
  wire [13:0] _GEN_11340 = 14'h2c4c == index ? 14'h8c : _GEN_11339;
  wire [13:0] _GEN_11341 = 14'h2c4d == index ? 14'h8b : _GEN_11340;
  wire [13:0] _GEN_11342 = 14'h2c4e == index ? 14'h8a : _GEN_11341;
  wire [13:0] _GEN_11343 = 14'h2c4f == index ? 14'h89 : _GEN_11342;
  wire [13:0] _GEN_11344 = 14'h2c50 == index ? 14'h88 : _GEN_11343;
  wire [13:0] _GEN_11345 = 14'h2c51 == index ? 14'h87 : _GEN_11344;
  wire [13:0] _GEN_11346 = 14'h2c52 == index ? 14'h86 : _GEN_11345;
  wire [13:0] _GEN_11347 = 14'h2c53 == index ? 14'h85 : _GEN_11346;
  wire [13:0] _GEN_11348 = 14'h2c54 == index ? 14'h84 : _GEN_11347;
  wire [13:0] _GEN_11349 = 14'h2c55 == index ? 14'h83 : _GEN_11348;
  wire [13:0] _GEN_11350 = 14'h2c56 == index ? 14'h82 : _GEN_11349;
  wire [13:0] _GEN_11351 = 14'h2c57 == index ? 14'h81 : _GEN_11350;
  wire [13:0] _GEN_11352 = 14'h2c58 == index ? 14'h80 : _GEN_11351;
  wire [13:0] _GEN_11353 = 14'h2c59 == index ? 14'h58 : _GEN_11352;
  wire [13:0] _GEN_11354 = 14'h2c5a == index ? 14'h58 : _GEN_11353;
  wire [13:0] _GEN_11355 = 14'h2c5b == index ? 14'h58 : _GEN_11354;
  wire [13:0] _GEN_11356 = 14'h2c5c == index ? 14'h58 : _GEN_11355;
  wire [13:0] _GEN_11357 = 14'h2c5d == index ? 14'h58 : _GEN_11356;
  wire [13:0] _GEN_11358 = 14'h2c5e == index ? 14'h58 : _GEN_11357;
  wire [13:0] _GEN_11359 = 14'h2c5f == index ? 14'h58 : _GEN_11358;
  wire [13:0] _GEN_11360 = 14'h2c60 == index ? 14'h58 : _GEN_11359;
  wire [13:0] _GEN_11361 = 14'h2c61 == index ? 14'h58 : _GEN_11360;
  wire [13:0] _GEN_11362 = 14'h2c62 == index ? 14'h58 : _GEN_11361;
  wire [13:0] _GEN_11363 = 14'h2c63 == index ? 14'h58 : _GEN_11362;
  wire [13:0] _GEN_11364 = 14'h2c64 == index ? 14'h58 : _GEN_11363;
  wire [13:0] _GEN_11365 = 14'h2c65 == index ? 14'h58 : _GEN_11364;
  wire [13:0] _GEN_11366 = 14'h2c66 == index ? 14'h58 : _GEN_11365;
  wire [13:0] _GEN_11367 = 14'h2c67 == index ? 14'h58 : _GEN_11366;
  wire [13:0] _GEN_11368 = 14'h2c68 == index ? 14'h58 : _GEN_11367;
  wire [13:0] _GEN_11369 = 14'h2c69 == index ? 14'h58 : _GEN_11368;
  wire [13:0] _GEN_11370 = 14'h2c6a == index ? 14'h58 : _GEN_11369;
  wire [13:0] _GEN_11371 = 14'h2c6b == index ? 14'h58 : _GEN_11370;
  wire [13:0] _GEN_11372 = 14'h2c6c == index ? 14'h58 : _GEN_11371;
  wire [13:0] _GEN_11373 = 14'h2c6d == index ? 14'h58 : _GEN_11372;
  wire [13:0] _GEN_11374 = 14'h2c6e == index ? 14'h58 : _GEN_11373;
  wire [13:0] _GEN_11375 = 14'h2c6f == index ? 14'h58 : _GEN_11374;
  wire [13:0] _GEN_11376 = 14'h2c70 == index ? 14'h58 : _GEN_11375;
  wire [13:0] _GEN_11377 = 14'h2c71 == index ? 14'h58 : _GEN_11376;
  wire [13:0] _GEN_11378 = 14'h2c72 == index ? 14'h58 : _GEN_11377;
  wire [13:0] _GEN_11379 = 14'h2c73 == index ? 14'h58 : _GEN_11378;
  wire [13:0] _GEN_11380 = 14'h2c74 == index ? 14'h58 : _GEN_11379;
  wire [13:0] _GEN_11381 = 14'h2c75 == index ? 14'h58 : _GEN_11380;
  wire [13:0] _GEN_11382 = 14'h2c76 == index ? 14'h58 : _GEN_11381;
  wire [13:0] _GEN_11383 = 14'h2c77 == index ? 14'h58 : _GEN_11382;
  wire [13:0] _GEN_11384 = 14'h2c78 == index ? 14'h58 : _GEN_11383;
  wire [13:0] _GEN_11385 = 14'h2c79 == index ? 14'h58 : _GEN_11384;
  wire [13:0] _GEN_11386 = 14'h2c7a == index ? 14'h58 : _GEN_11385;
  wire [13:0] _GEN_11387 = 14'h2c7b == index ? 14'h58 : _GEN_11386;
  wire [13:0] _GEN_11388 = 14'h2c7c == index ? 14'h58 : _GEN_11387;
  wire [13:0] _GEN_11389 = 14'h2c7d == index ? 14'h58 : _GEN_11388;
  wire [13:0] _GEN_11390 = 14'h2c7e == index ? 14'h58 : _GEN_11389;
  wire [13:0] _GEN_11391 = 14'h2c7f == index ? 14'h58 : _GEN_11390;
  wire [13:0] _GEN_11392 = 14'h2c80 == index ? 14'h0 : _GEN_11391;
  wire [13:0] _GEN_11393 = 14'h2c81 == index ? 14'h2c80 : _GEN_11392;
  wire [13:0] _GEN_11394 = 14'h2c82 == index ? 14'h1601 : _GEN_11393;
  wire [13:0] _GEN_11395 = 14'h2c83 == index ? 14'he82 : _GEN_11394;
  wire [13:0] _GEN_11396 = 14'h2c84 == index ? 14'hb01 : _GEN_11395;
  wire [13:0] _GEN_11397 = 14'h2c85 == index ? 14'h884 : _GEN_11396;
  wire [13:0] _GEN_11398 = 14'h2c86 == index ? 14'h705 : _GEN_11397;
  wire [13:0] _GEN_11399 = 14'h2c87 == index ? 14'h605 : _GEN_11398;
  wire [13:0] _GEN_11400 = 14'h2c88 == index ? 14'h581 : _GEN_11399;
  wire [13:0] _GEN_11401 = 14'h2c89 == index ? 14'h488 : _GEN_11400;
  wire [13:0] _GEN_11402 = 14'h2c8a == index ? 14'h409 : _GEN_11401;
  wire [13:0] _GEN_11403 = 14'h2c8b == index ? 14'h401 : _GEN_11402;
  wire [13:0] _GEN_11404 = 14'h2c8c == index ? 14'h385 : _GEN_11403;
  wire [13:0] _GEN_11405 = 14'h2c8d == index ? 14'h30b : _GEN_11404;
  wire [13:0] _GEN_11406 = 14'h2c8e == index ? 14'h305 : _GEN_11405;
  wire [13:0] _GEN_11407 = 14'h2c8f == index ? 14'h28e : _GEN_11406;
  wire [13:0] _GEN_11408 = 14'h2c90 == index ? 14'h289 : _GEN_11407;
  wire [13:0] _GEN_11409 = 14'h2c91 == index ? 14'h284 : _GEN_11408;
  wire [13:0] _GEN_11410 = 14'h2c92 == index ? 14'h211 : _GEN_11409;
  wire [13:0] _GEN_11411 = 14'h2c93 == index ? 14'h20d : _GEN_11410;
  wire [13:0] _GEN_11412 = 14'h2c94 == index ? 14'h209 : _GEN_11411;
  wire [13:0] _GEN_11413 = 14'h2c95 == index ? 14'h205 : _GEN_11412;
  wire [13:0] _GEN_11414 = 14'h2c96 == index ? 14'h201 : _GEN_11413;
  wire [13:0] _GEN_11415 = 14'h2c97 == index ? 14'h194 : _GEN_11414;
  wire [13:0] _GEN_11416 = 14'h2c98 == index ? 14'h191 : _GEN_11415;
  wire [13:0] _GEN_11417 = 14'h2c99 == index ? 14'h18e : _GEN_11416;
  wire [13:0] _GEN_11418 = 14'h2c9a == index ? 14'h18b : _GEN_11417;
  wire [13:0] _GEN_11419 = 14'h2c9b == index ? 14'h188 : _GEN_11418;
  wire [13:0] _GEN_11420 = 14'h2c9c == index ? 14'h185 : _GEN_11419;
  wire [13:0] _GEN_11421 = 14'h2c9d == index ? 14'h182 : _GEN_11420;
  wire [13:0] _GEN_11422 = 14'h2c9e == index ? 14'h11d : _GEN_11421;
  wire [13:0] _GEN_11423 = 14'h2c9f == index ? 14'h11b : _GEN_11422;
  wire [13:0] _GEN_11424 = 14'h2ca0 == index ? 14'h119 : _GEN_11423;
  wire [13:0] _GEN_11425 = 14'h2ca1 == index ? 14'h117 : _GEN_11424;
  wire [13:0] _GEN_11426 = 14'h2ca2 == index ? 14'h115 : _GEN_11425;
  wire [13:0] _GEN_11427 = 14'h2ca3 == index ? 14'h113 : _GEN_11426;
  wire [13:0] _GEN_11428 = 14'h2ca4 == index ? 14'h111 : _GEN_11427;
  wire [13:0] _GEN_11429 = 14'h2ca5 == index ? 14'h10f : _GEN_11428;
  wire [13:0] _GEN_11430 = 14'h2ca6 == index ? 14'h10d : _GEN_11429;
  wire [13:0] _GEN_11431 = 14'h2ca7 == index ? 14'h10b : _GEN_11430;
  wire [13:0] _GEN_11432 = 14'h2ca8 == index ? 14'h109 : _GEN_11431;
  wire [13:0] _GEN_11433 = 14'h2ca9 == index ? 14'h107 : _GEN_11432;
  wire [13:0] _GEN_11434 = 14'h2caa == index ? 14'h105 : _GEN_11433;
  wire [13:0] _GEN_11435 = 14'h2cab == index ? 14'h103 : _GEN_11434;
  wire [13:0] _GEN_11436 = 14'h2cac == index ? 14'h101 : _GEN_11435;
  wire [13:0] _GEN_11437 = 14'h2cad == index ? 14'hac : _GEN_11436;
  wire [13:0] _GEN_11438 = 14'h2cae == index ? 14'hab : _GEN_11437;
  wire [13:0] _GEN_11439 = 14'h2caf == index ? 14'haa : _GEN_11438;
  wire [13:0] _GEN_11440 = 14'h2cb0 == index ? 14'ha9 : _GEN_11439;
  wire [13:0] _GEN_11441 = 14'h2cb1 == index ? 14'ha8 : _GEN_11440;
  wire [13:0] _GEN_11442 = 14'h2cb2 == index ? 14'ha7 : _GEN_11441;
  wire [13:0] _GEN_11443 = 14'h2cb3 == index ? 14'ha6 : _GEN_11442;
  wire [13:0] _GEN_11444 = 14'h2cb4 == index ? 14'ha5 : _GEN_11443;
  wire [13:0] _GEN_11445 = 14'h2cb5 == index ? 14'ha4 : _GEN_11444;
  wire [13:0] _GEN_11446 = 14'h2cb6 == index ? 14'ha3 : _GEN_11445;
  wire [13:0] _GEN_11447 = 14'h2cb7 == index ? 14'ha2 : _GEN_11446;
  wire [13:0] _GEN_11448 = 14'h2cb8 == index ? 14'ha1 : _GEN_11447;
  wire [13:0] _GEN_11449 = 14'h2cb9 == index ? 14'ha0 : _GEN_11448;
  wire [13:0] _GEN_11450 = 14'h2cba == index ? 14'h9f : _GEN_11449;
  wire [13:0] _GEN_11451 = 14'h2cbb == index ? 14'h9e : _GEN_11450;
  wire [13:0] _GEN_11452 = 14'h2cbc == index ? 14'h9d : _GEN_11451;
  wire [13:0] _GEN_11453 = 14'h2cbd == index ? 14'h9c : _GEN_11452;
  wire [13:0] _GEN_11454 = 14'h2cbe == index ? 14'h9b : _GEN_11453;
  wire [13:0] _GEN_11455 = 14'h2cbf == index ? 14'h9a : _GEN_11454;
  wire [13:0] _GEN_11456 = 14'h2cc0 == index ? 14'h99 : _GEN_11455;
  wire [13:0] _GEN_11457 = 14'h2cc1 == index ? 14'h98 : _GEN_11456;
  wire [13:0] _GEN_11458 = 14'h2cc2 == index ? 14'h97 : _GEN_11457;
  wire [13:0] _GEN_11459 = 14'h2cc3 == index ? 14'h96 : _GEN_11458;
  wire [13:0] _GEN_11460 = 14'h2cc4 == index ? 14'h95 : _GEN_11459;
  wire [13:0] _GEN_11461 = 14'h2cc5 == index ? 14'h94 : _GEN_11460;
  wire [13:0] _GEN_11462 = 14'h2cc6 == index ? 14'h93 : _GEN_11461;
  wire [13:0] _GEN_11463 = 14'h2cc7 == index ? 14'h92 : _GEN_11462;
  wire [13:0] _GEN_11464 = 14'h2cc8 == index ? 14'h91 : _GEN_11463;
  wire [13:0] _GEN_11465 = 14'h2cc9 == index ? 14'h90 : _GEN_11464;
  wire [13:0] _GEN_11466 = 14'h2cca == index ? 14'h8f : _GEN_11465;
  wire [13:0] _GEN_11467 = 14'h2ccb == index ? 14'h8e : _GEN_11466;
  wire [13:0] _GEN_11468 = 14'h2ccc == index ? 14'h8d : _GEN_11467;
  wire [13:0] _GEN_11469 = 14'h2ccd == index ? 14'h8c : _GEN_11468;
  wire [13:0] _GEN_11470 = 14'h2cce == index ? 14'h8b : _GEN_11469;
  wire [13:0] _GEN_11471 = 14'h2ccf == index ? 14'h8a : _GEN_11470;
  wire [13:0] _GEN_11472 = 14'h2cd0 == index ? 14'h89 : _GEN_11471;
  wire [13:0] _GEN_11473 = 14'h2cd1 == index ? 14'h88 : _GEN_11472;
  wire [13:0] _GEN_11474 = 14'h2cd2 == index ? 14'h87 : _GEN_11473;
  wire [13:0] _GEN_11475 = 14'h2cd3 == index ? 14'h86 : _GEN_11474;
  wire [13:0] _GEN_11476 = 14'h2cd4 == index ? 14'h85 : _GEN_11475;
  wire [13:0] _GEN_11477 = 14'h2cd5 == index ? 14'h84 : _GEN_11476;
  wire [13:0] _GEN_11478 = 14'h2cd6 == index ? 14'h83 : _GEN_11477;
  wire [13:0] _GEN_11479 = 14'h2cd7 == index ? 14'h82 : _GEN_11478;
  wire [13:0] _GEN_11480 = 14'h2cd8 == index ? 14'h81 : _GEN_11479;
  wire [13:0] _GEN_11481 = 14'h2cd9 == index ? 14'h80 : _GEN_11480;
  wire [13:0] _GEN_11482 = 14'h2cda == index ? 14'h59 : _GEN_11481;
  wire [13:0] _GEN_11483 = 14'h2cdb == index ? 14'h59 : _GEN_11482;
  wire [13:0] _GEN_11484 = 14'h2cdc == index ? 14'h59 : _GEN_11483;
  wire [13:0] _GEN_11485 = 14'h2cdd == index ? 14'h59 : _GEN_11484;
  wire [13:0] _GEN_11486 = 14'h2cde == index ? 14'h59 : _GEN_11485;
  wire [13:0] _GEN_11487 = 14'h2cdf == index ? 14'h59 : _GEN_11486;
  wire [13:0] _GEN_11488 = 14'h2ce0 == index ? 14'h59 : _GEN_11487;
  wire [13:0] _GEN_11489 = 14'h2ce1 == index ? 14'h59 : _GEN_11488;
  wire [13:0] _GEN_11490 = 14'h2ce2 == index ? 14'h59 : _GEN_11489;
  wire [13:0] _GEN_11491 = 14'h2ce3 == index ? 14'h59 : _GEN_11490;
  wire [13:0] _GEN_11492 = 14'h2ce4 == index ? 14'h59 : _GEN_11491;
  wire [13:0] _GEN_11493 = 14'h2ce5 == index ? 14'h59 : _GEN_11492;
  wire [13:0] _GEN_11494 = 14'h2ce6 == index ? 14'h59 : _GEN_11493;
  wire [13:0] _GEN_11495 = 14'h2ce7 == index ? 14'h59 : _GEN_11494;
  wire [13:0] _GEN_11496 = 14'h2ce8 == index ? 14'h59 : _GEN_11495;
  wire [13:0] _GEN_11497 = 14'h2ce9 == index ? 14'h59 : _GEN_11496;
  wire [13:0] _GEN_11498 = 14'h2cea == index ? 14'h59 : _GEN_11497;
  wire [13:0] _GEN_11499 = 14'h2ceb == index ? 14'h59 : _GEN_11498;
  wire [13:0] _GEN_11500 = 14'h2cec == index ? 14'h59 : _GEN_11499;
  wire [13:0] _GEN_11501 = 14'h2ced == index ? 14'h59 : _GEN_11500;
  wire [13:0] _GEN_11502 = 14'h2cee == index ? 14'h59 : _GEN_11501;
  wire [13:0] _GEN_11503 = 14'h2cef == index ? 14'h59 : _GEN_11502;
  wire [13:0] _GEN_11504 = 14'h2cf0 == index ? 14'h59 : _GEN_11503;
  wire [13:0] _GEN_11505 = 14'h2cf1 == index ? 14'h59 : _GEN_11504;
  wire [13:0] _GEN_11506 = 14'h2cf2 == index ? 14'h59 : _GEN_11505;
  wire [13:0] _GEN_11507 = 14'h2cf3 == index ? 14'h59 : _GEN_11506;
  wire [13:0] _GEN_11508 = 14'h2cf4 == index ? 14'h59 : _GEN_11507;
  wire [13:0] _GEN_11509 = 14'h2cf5 == index ? 14'h59 : _GEN_11508;
  wire [13:0] _GEN_11510 = 14'h2cf6 == index ? 14'h59 : _GEN_11509;
  wire [13:0] _GEN_11511 = 14'h2cf7 == index ? 14'h59 : _GEN_11510;
  wire [13:0] _GEN_11512 = 14'h2cf8 == index ? 14'h59 : _GEN_11511;
  wire [13:0] _GEN_11513 = 14'h2cf9 == index ? 14'h59 : _GEN_11512;
  wire [13:0] _GEN_11514 = 14'h2cfa == index ? 14'h59 : _GEN_11513;
  wire [13:0] _GEN_11515 = 14'h2cfb == index ? 14'h59 : _GEN_11514;
  wire [13:0] _GEN_11516 = 14'h2cfc == index ? 14'h59 : _GEN_11515;
  wire [13:0] _GEN_11517 = 14'h2cfd == index ? 14'h59 : _GEN_11516;
  wire [13:0] _GEN_11518 = 14'h2cfe == index ? 14'h59 : _GEN_11517;
  wire [13:0] _GEN_11519 = 14'h2cff == index ? 14'h59 : _GEN_11518;
  wire [13:0] _GEN_11520 = 14'h2d00 == index ? 14'h0 : _GEN_11519;
  wire [13:0] _GEN_11521 = 14'h2d01 == index ? 14'h2d00 : _GEN_11520;
  wire [13:0] _GEN_11522 = 14'h2d02 == index ? 14'h1680 : _GEN_11521;
  wire [13:0] _GEN_11523 = 14'h2d03 == index ? 14'hf00 : _GEN_11522;
  wire [13:0] _GEN_11524 = 14'h2d04 == index ? 14'hb02 : _GEN_11523;
  wire [13:0] _GEN_11525 = 14'h2d05 == index ? 14'h900 : _GEN_11524;
  wire [13:0] _GEN_11526 = 14'h2d06 == index ? 14'h780 : _GEN_11525;
  wire [13:0] _GEN_11527 = 14'h2d07 == index ? 14'h606 : _GEN_11526;
  wire [13:0] _GEN_11528 = 14'h2d08 == index ? 14'h582 : _GEN_11527;
  wire [13:0] _GEN_11529 = 14'h2d09 == index ? 14'h500 : _GEN_11528;
  wire [13:0] _GEN_11530 = 14'h2d0a == index ? 14'h480 : _GEN_11529;
  wire [13:0] _GEN_11531 = 14'h2d0b == index ? 14'h402 : _GEN_11530;
  wire [13:0] _GEN_11532 = 14'h2d0c == index ? 14'h386 : _GEN_11531;
  wire [13:0] _GEN_11533 = 14'h2d0d == index ? 14'h30c : _GEN_11532;
  wire [13:0] _GEN_11534 = 14'h2d0e == index ? 14'h306 : _GEN_11533;
  wire [13:0] _GEN_11535 = 14'h2d0f == index ? 14'h300 : _GEN_11534;
  wire [13:0] _GEN_11536 = 14'h2d10 == index ? 14'h28a : _GEN_11535;
  wire [13:0] _GEN_11537 = 14'h2d11 == index ? 14'h285 : _GEN_11536;
  wire [13:0] _GEN_11538 = 14'h2d12 == index ? 14'h280 : _GEN_11537;
  wire [13:0] _GEN_11539 = 14'h2d13 == index ? 14'h20e : _GEN_11538;
  wire [13:0] _GEN_11540 = 14'h2d14 == index ? 14'h20a : _GEN_11539;
  wire [13:0] _GEN_11541 = 14'h2d15 == index ? 14'h206 : _GEN_11540;
  wire [13:0] _GEN_11542 = 14'h2d16 == index ? 14'h202 : _GEN_11541;
  wire [13:0] _GEN_11543 = 14'h2d17 == index ? 14'h195 : _GEN_11542;
  wire [13:0] _GEN_11544 = 14'h2d18 == index ? 14'h192 : _GEN_11543;
  wire [13:0] _GEN_11545 = 14'h2d19 == index ? 14'h18f : _GEN_11544;
  wire [13:0] _GEN_11546 = 14'h2d1a == index ? 14'h18c : _GEN_11545;
  wire [13:0] _GEN_11547 = 14'h2d1b == index ? 14'h189 : _GEN_11546;
  wire [13:0] _GEN_11548 = 14'h2d1c == index ? 14'h186 : _GEN_11547;
  wire [13:0] _GEN_11549 = 14'h2d1d == index ? 14'h183 : _GEN_11548;
  wire [13:0] _GEN_11550 = 14'h2d1e == index ? 14'h180 : _GEN_11549;
  wire [13:0] _GEN_11551 = 14'h2d1f == index ? 14'h11c : _GEN_11550;
  wire [13:0] _GEN_11552 = 14'h2d20 == index ? 14'h11a : _GEN_11551;
  wire [13:0] _GEN_11553 = 14'h2d21 == index ? 14'h118 : _GEN_11552;
  wire [13:0] _GEN_11554 = 14'h2d22 == index ? 14'h116 : _GEN_11553;
  wire [13:0] _GEN_11555 = 14'h2d23 == index ? 14'h114 : _GEN_11554;
  wire [13:0] _GEN_11556 = 14'h2d24 == index ? 14'h112 : _GEN_11555;
  wire [13:0] _GEN_11557 = 14'h2d25 == index ? 14'h110 : _GEN_11556;
  wire [13:0] _GEN_11558 = 14'h2d26 == index ? 14'h10e : _GEN_11557;
  wire [13:0] _GEN_11559 = 14'h2d27 == index ? 14'h10c : _GEN_11558;
  wire [13:0] _GEN_11560 = 14'h2d28 == index ? 14'h10a : _GEN_11559;
  wire [13:0] _GEN_11561 = 14'h2d29 == index ? 14'h108 : _GEN_11560;
  wire [13:0] _GEN_11562 = 14'h2d2a == index ? 14'h106 : _GEN_11561;
  wire [13:0] _GEN_11563 = 14'h2d2b == index ? 14'h104 : _GEN_11562;
  wire [13:0] _GEN_11564 = 14'h2d2c == index ? 14'h102 : _GEN_11563;
  wire [13:0] _GEN_11565 = 14'h2d2d == index ? 14'h100 : _GEN_11564;
  wire [13:0] _GEN_11566 = 14'h2d2e == index ? 14'hac : _GEN_11565;
  wire [13:0] _GEN_11567 = 14'h2d2f == index ? 14'hab : _GEN_11566;
  wire [13:0] _GEN_11568 = 14'h2d30 == index ? 14'haa : _GEN_11567;
  wire [13:0] _GEN_11569 = 14'h2d31 == index ? 14'ha9 : _GEN_11568;
  wire [13:0] _GEN_11570 = 14'h2d32 == index ? 14'ha8 : _GEN_11569;
  wire [13:0] _GEN_11571 = 14'h2d33 == index ? 14'ha7 : _GEN_11570;
  wire [13:0] _GEN_11572 = 14'h2d34 == index ? 14'ha6 : _GEN_11571;
  wire [13:0] _GEN_11573 = 14'h2d35 == index ? 14'ha5 : _GEN_11572;
  wire [13:0] _GEN_11574 = 14'h2d36 == index ? 14'ha4 : _GEN_11573;
  wire [13:0] _GEN_11575 = 14'h2d37 == index ? 14'ha3 : _GEN_11574;
  wire [13:0] _GEN_11576 = 14'h2d38 == index ? 14'ha2 : _GEN_11575;
  wire [13:0] _GEN_11577 = 14'h2d39 == index ? 14'ha1 : _GEN_11576;
  wire [13:0] _GEN_11578 = 14'h2d3a == index ? 14'ha0 : _GEN_11577;
  wire [13:0] _GEN_11579 = 14'h2d3b == index ? 14'h9f : _GEN_11578;
  wire [13:0] _GEN_11580 = 14'h2d3c == index ? 14'h9e : _GEN_11579;
  wire [13:0] _GEN_11581 = 14'h2d3d == index ? 14'h9d : _GEN_11580;
  wire [13:0] _GEN_11582 = 14'h2d3e == index ? 14'h9c : _GEN_11581;
  wire [13:0] _GEN_11583 = 14'h2d3f == index ? 14'h9b : _GEN_11582;
  wire [13:0] _GEN_11584 = 14'h2d40 == index ? 14'h9a : _GEN_11583;
  wire [13:0] _GEN_11585 = 14'h2d41 == index ? 14'h99 : _GEN_11584;
  wire [13:0] _GEN_11586 = 14'h2d42 == index ? 14'h98 : _GEN_11585;
  wire [13:0] _GEN_11587 = 14'h2d43 == index ? 14'h97 : _GEN_11586;
  wire [13:0] _GEN_11588 = 14'h2d44 == index ? 14'h96 : _GEN_11587;
  wire [13:0] _GEN_11589 = 14'h2d45 == index ? 14'h95 : _GEN_11588;
  wire [13:0] _GEN_11590 = 14'h2d46 == index ? 14'h94 : _GEN_11589;
  wire [13:0] _GEN_11591 = 14'h2d47 == index ? 14'h93 : _GEN_11590;
  wire [13:0] _GEN_11592 = 14'h2d48 == index ? 14'h92 : _GEN_11591;
  wire [13:0] _GEN_11593 = 14'h2d49 == index ? 14'h91 : _GEN_11592;
  wire [13:0] _GEN_11594 = 14'h2d4a == index ? 14'h90 : _GEN_11593;
  wire [13:0] _GEN_11595 = 14'h2d4b == index ? 14'h8f : _GEN_11594;
  wire [13:0] _GEN_11596 = 14'h2d4c == index ? 14'h8e : _GEN_11595;
  wire [13:0] _GEN_11597 = 14'h2d4d == index ? 14'h8d : _GEN_11596;
  wire [13:0] _GEN_11598 = 14'h2d4e == index ? 14'h8c : _GEN_11597;
  wire [13:0] _GEN_11599 = 14'h2d4f == index ? 14'h8b : _GEN_11598;
  wire [13:0] _GEN_11600 = 14'h2d50 == index ? 14'h8a : _GEN_11599;
  wire [13:0] _GEN_11601 = 14'h2d51 == index ? 14'h89 : _GEN_11600;
  wire [13:0] _GEN_11602 = 14'h2d52 == index ? 14'h88 : _GEN_11601;
  wire [13:0] _GEN_11603 = 14'h2d53 == index ? 14'h87 : _GEN_11602;
  wire [13:0] _GEN_11604 = 14'h2d54 == index ? 14'h86 : _GEN_11603;
  wire [13:0] _GEN_11605 = 14'h2d55 == index ? 14'h85 : _GEN_11604;
  wire [13:0] _GEN_11606 = 14'h2d56 == index ? 14'h84 : _GEN_11605;
  wire [13:0] _GEN_11607 = 14'h2d57 == index ? 14'h83 : _GEN_11606;
  wire [13:0] _GEN_11608 = 14'h2d58 == index ? 14'h82 : _GEN_11607;
  wire [13:0] _GEN_11609 = 14'h2d59 == index ? 14'h81 : _GEN_11608;
  wire [13:0] _GEN_11610 = 14'h2d5a == index ? 14'h80 : _GEN_11609;
  wire [13:0] _GEN_11611 = 14'h2d5b == index ? 14'h5a : _GEN_11610;
  wire [13:0] _GEN_11612 = 14'h2d5c == index ? 14'h5a : _GEN_11611;
  wire [13:0] _GEN_11613 = 14'h2d5d == index ? 14'h5a : _GEN_11612;
  wire [13:0] _GEN_11614 = 14'h2d5e == index ? 14'h5a : _GEN_11613;
  wire [13:0] _GEN_11615 = 14'h2d5f == index ? 14'h5a : _GEN_11614;
  wire [13:0] _GEN_11616 = 14'h2d60 == index ? 14'h5a : _GEN_11615;
  wire [13:0] _GEN_11617 = 14'h2d61 == index ? 14'h5a : _GEN_11616;
  wire [13:0] _GEN_11618 = 14'h2d62 == index ? 14'h5a : _GEN_11617;
  wire [13:0] _GEN_11619 = 14'h2d63 == index ? 14'h5a : _GEN_11618;
  wire [13:0] _GEN_11620 = 14'h2d64 == index ? 14'h5a : _GEN_11619;
  wire [13:0] _GEN_11621 = 14'h2d65 == index ? 14'h5a : _GEN_11620;
  wire [13:0] _GEN_11622 = 14'h2d66 == index ? 14'h5a : _GEN_11621;
  wire [13:0] _GEN_11623 = 14'h2d67 == index ? 14'h5a : _GEN_11622;
  wire [13:0] _GEN_11624 = 14'h2d68 == index ? 14'h5a : _GEN_11623;
  wire [13:0] _GEN_11625 = 14'h2d69 == index ? 14'h5a : _GEN_11624;
  wire [13:0] _GEN_11626 = 14'h2d6a == index ? 14'h5a : _GEN_11625;
  wire [13:0] _GEN_11627 = 14'h2d6b == index ? 14'h5a : _GEN_11626;
  wire [13:0] _GEN_11628 = 14'h2d6c == index ? 14'h5a : _GEN_11627;
  wire [13:0] _GEN_11629 = 14'h2d6d == index ? 14'h5a : _GEN_11628;
  wire [13:0] _GEN_11630 = 14'h2d6e == index ? 14'h5a : _GEN_11629;
  wire [13:0] _GEN_11631 = 14'h2d6f == index ? 14'h5a : _GEN_11630;
  wire [13:0] _GEN_11632 = 14'h2d70 == index ? 14'h5a : _GEN_11631;
  wire [13:0] _GEN_11633 = 14'h2d71 == index ? 14'h5a : _GEN_11632;
  wire [13:0] _GEN_11634 = 14'h2d72 == index ? 14'h5a : _GEN_11633;
  wire [13:0] _GEN_11635 = 14'h2d73 == index ? 14'h5a : _GEN_11634;
  wire [13:0] _GEN_11636 = 14'h2d74 == index ? 14'h5a : _GEN_11635;
  wire [13:0] _GEN_11637 = 14'h2d75 == index ? 14'h5a : _GEN_11636;
  wire [13:0] _GEN_11638 = 14'h2d76 == index ? 14'h5a : _GEN_11637;
  wire [13:0] _GEN_11639 = 14'h2d77 == index ? 14'h5a : _GEN_11638;
  wire [13:0] _GEN_11640 = 14'h2d78 == index ? 14'h5a : _GEN_11639;
  wire [13:0] _GEN_11641 = 14'h2d79 == index ? 14'h5a : _GEN_11640;
  wire [13:0] _GEN_11642 = 14'h2d7a == index ? 14'h5a : _GEN_11641;
  wire [13:0] _GEN_11643 = 14'h2d7b == index ? 14'h5a : _GEN_11642;
  wire [13:0] _GEN_11644 = 14'h2d7c == index ? 14'h5a : _GEN_11643;
  wire [13:0] _GEN_11645 = 14'h2d7d == index ? 14'h5a : _GEN_11644;
  wire [13:0] _GEN_11646 = 14'h2d7e == index ? 14'h5a : _GEN_11645;
  wire [13:0] _GEN_11647 = 14'h2d7f == index ? 14'h5a : _GEN_11646;
  wire [13:0] _GEN_11648 = 14'h2d80 == index ? 14'h0 : _GEN_11647;
  wire [13:0] _GEN_11649 = 14'h2d81 == index ? 14'h2d80 : _GEN_11648;
  wire [13:0] _GEN_11650 = 14'h2d82 == index ? 14'h1681 : _GEN_11649;
  wire [13:0] _GEN_11651 = 14'h2d83 == index ? 14'hf01 : _GEN_11650;
  wire [13:0] _GEN_11652 = 14'h2d84 == index ? 14'hb03 : _GEN_11651;
  wire [13:0] _GEN_11653 = 14'h2d85 == index ? 14'h901 : _GEN_11652;
  wire [13:0] _GEN_11654 = 14'h2d86 == index ? 14'h781 : _GEN_11653;
  wire [13:0] _GEN_11655 = 14'h2d87 == index ? 14'h680 : _GEN_11654;
  wire [13:0] _GEN_11656 = 14'h2d88 == index ? 14'h583 : _GEN_11655;
  wire [13:0] _GEN_11657 = 14'h2d89 == index ? 14'h501 : _GEN_11656;
  wire [13:0] _GEN_11658 = 14'h2d8a == index ? 14'h481 : _GEN_11657;
  wire [13:0] _GEN_11659 = 14'h2d8b == index ? 14'h403 : _GEN_11658;
  wire [13:0] _GEN_11660 = 14'h2d8c == index ? 14'h387 : _GEN_11659;
  wire [13:0] _GEN_11661 = 14'h2d8d == index ? 14'h380 : _GEN_11660;
  wire [13:0] _GEN_11662 = 14'h2d8e == index ? 14'h307 : _GEN_11661;
  wire [13:0] _GEN_11663 = 14'h2d8f == index ? 14'h301 : _GEN_11662;
  wire [13:0] _GEN_11664 = 14'h2d90 == index ? 14'h28b : _GEN_11663;
  wire [13:0] _GEN_11665 = 14'h2d91 == index ? 14'h286 : _GEN_11664;
  wire [13:0] _GEN_11666 = 14'h2d92 == index ? 14'h281 : _GEN_11665;
  wire [13:0] _GEN_11667 = 14'h2d93 == index ? 14'h20f : _GEN_11666;
  wire [13:0] _GEN_11668 = 14'h2d94 == index ? 14'h20b : _GEN_11667;
  wire [13:0] _GEN_11669 = 14'h2d95 == index ? 14'h207 : _GEN_11668;
  wire [13:0] _GEN_11670 = 14'h2d96 == index ? 14'h203 : _GEN_11669;
  wire [13:0] _GEN_11671 = 14'h2d97 == index ? 14'h196 : _GEN_11670;
  wire [13:0] _GEN_11672 = 14'h2d98 == index ? 14'h193 : _GEN_11671;
  wire [13:0] _GEN_11673 = 14'h2d99 == index ? 14'h190 : _GEN_11672;
  wire [13:0] _GEN_11674 = 14'h2d9a == index ? 14'h18d : _GEN_11673;
  wire [13:0] _GEN_11675 = 14'h2d9b == index ? 14'h18a : _GEN_11674;
  wire [13:0] _GEN_11676 = 14'h2d9c == index ? 14'h187 : _GEN_11675;
  wire [13:0] _GEN_11677 = 14'h2d9d == index ? 14'h184 : _GEN_11676;
  wire [13:0] _GEN_11678 = 14'h2d9e == index ? 14'h181 : _GEN_11677;
  wire [13:0] _GEN_11679 = 14'h2d9f == index ? 14'h11d : _GEN_11678;
  wire [13:0] _GEN_11680 = 14'h2da0 == index ? 14'h11b : _GEN_11679;
  wire [13:0] _GEN_11681 = 14'h2da1 == index ? 14'h119 : _GEN_11680;
  wire [13:0] _GEN_11682 = 14'h2da2 == index ? 14'h117 : _GEN_11681;
  wire [13:0] _GEN_11683 = 14'h2da3 == index ? 14'h115 : _GEN_11682;
  wire [13:0] _GEN_11684 = 14'h2da4 == index ? 14'h113 : _GEN_11683;
  wire [13:0] _GEN_11685 = 14'h2da5 == index ? 14'h111 : _GEN_11684;
  wire [13:0] _GEN_11686 = 14'h2da6 == index ? 14'h10f : _GEN_11685;
  wire [13:0] _GEN_11687 = 14'h2da7 == index ? 14'h10d : _GEN_11686;
  wire [13:0] _GEN_11688 = 14'h2da8 == index ? 14'h10b : _GEN_11687;
  wire [13:0] _GEN_11689 = 14'h2da9 == index ? 14'h109 : _GEN_11688;
  wire [13:0] _GEN_11690 = 14'h2daa == index ? 14'h107 : _GEN_11689;
  wire [13:0] _GEN_11691 = 14'h2dab == index ? 14'h105 : _GEN_11690;
  wire [13:0] _GEN_11692 = 14'h2dac == index ? 14'h103 : _GEN_11691;
  wire [13:0] _GEN_11693 = 14'h2dad == index ? 14'h101 : _GEN_11692;
  wire [13:0] _GEN_11694 = 14'h2dae == index ? 14'had : _GEN_11693;
  wire [13:0] _GEN_11695 = 14'h2daf == index ? 14'hac : _GEN_11694;
  wire [13:0] _GEN_11696 = 14'h2db0 == index ? 14'hab : _GEN_11695;
  wire [13:0] _GEN_11697 = 14'h2db1 == index ? 14'haa : _GEN_11696;
  wire [13:0] _GEN_11698 = 14'h2db2 == index ? 14'ha9 : _GEN_11697;
  wire [13:0] _GEN_11699 = 14'h2db3 == index ? 14'ha8 : _GEN_11698;
  wire [13:0] _GEN_11700 = 14'h2db4 == index ? 14'ha7 : _GEN_11699;
  wire [13:0] _GEN_11701 = 14'h2db5 == index ? 14'ha6 : _GEN_11700;
  wire [13:0] _GEN_11702 = 14'h2db6 == index ? 14'ha5 : _GEN_11701;
  wire [13:0] _GEN_11703 = 14'h2db7 == index ? 14'ha4 : _GEN_11702;
  wire [13:0] _GEN_11704 = 14'h2db8 == index ? 14'ha3 : _GEN_11703;
  wire [13:0] _GEN_11705 = 14'h2db9 == index ? 14'ha2 : _GEN_11704;
  wire [13:0] _GEN_11706 = 14'h2dba == index ? 14'ha1 : _GEN_11705;
  wire [13:0] _GEN_11707 = 14'h2dbb == index ? 14'ha0 : _GEN_11706;
  wire [13:0] _GEN_11708 = 14'h2dbc == index ? 14'h9f : _GEN_11707;
  wire [13:0] _GEN_11709 = 14'h2dbd == index ? 14'h9e : _GEN_11708;
  wire [13:0] _GEN_11710 = 14'h2dbe == index ? 14'h9d : _GEN_11709;
  wire [13:0] _GEN_11711 = 14'h2dbf == index ? 14'h9c : _GEN_11710;
  wire [13:0] _GEN_11712 = 14'h2dc0 == index ? 14'h9b : _GEN_11711;
  wire [13:0] _GEN_11713 = 14'h2dc1 == index ? 14'h9a : _GEN_11712;
  wire [13:0] _GEN_11714 = 14'h2dc2 == index ? 14'h99 : _GEN_11713;
  wire [13:0] _GEN_11715 = 14'h2dc3 == index ? 14'h98 : _GEN_11714;
  wire [13:0] _GEN_11716 = 14'h2dc4 == index ? 14'h97 : _GEN_11715;
  wire [13:0] _GEN_11717 = 14'h2dc5 == index ? 14'h96 : _GEN_11716;
  wire [13:0] _GEN_11718 = 14'h2dc6 == index ? 14'h95 : _GEN_11717;
  wire [13:0] _GEN_11719 = 14'h2dc7 == index ? 14'h94 : _GEN_11718;
  wire [13:0] _GEN_11720 = 14'h2dc8 == index ? 14'h93 : _GEN_11719;
  wire [13:0] _GEN_11721 = 14'h2dc9 == index ? 14'h92 : _GEN_11720;
  wire [13:0] _GEN_11722 = 14'h2dca == index ? 14'h91 : _GEN_11721;
  wire [13:0] _GEN_11723 = 14'h2dcb == index ? 14'h90 : _GEN_11722;
  wire [13:0] _GEN_11724 = 14'h2dcc == index ? 14'h8f : _GEN_11723;
  wire [13:0] _GEN_11725 = 14'h2dcd == index ? 14'h8e : _GEN_11724;
  wire [13:0] _GEN_11726 = 14'h2dce == index ? 14'h8d : _GEN_11725;
  wire [13:0] _GEN_11727 = 14'h2dcf == index ? 14'h8c : _GEN_11726;
  wire [13:0] _GEN_11728 = 14'h2dd0 == index ? 14'h8b : _GEN_11727;
  wire [13:0] _GEN_11729 = 14'h2dd1 == index ? 14'h8a : _GEN_11728;
  wire [13:0] _GEN_11730 = 14'h2dd2 == index ? 14'h89 : _GEN_11729;
  wire [13:0] _GEN_11731 = 14'h2dd3 == index ? 14'h88 : _GEN_11730;
  wire [13:0] _GEN_11732 = 14'h2dd4 == index ? 14'h87 : _GEN_11731;
  wire [13:0] _GEN_11733 = 14'h2dd5 == index ? 14'h86 : _GEN_11732;
  wire [13:0] _GEN_11734 = 14'h2dd6 == index ? 14'h85 : _GEN_11733;
  wire [13:0] _GEN_11735 = 14'h2dd7 == index ? 14'h84 : _GEN_11734;
  wire [13:0] _GEN_11736 = 14'h2dd8 == index ? 14'h83 : _GEN_11735;
  wire [13:0] _GEN_11737 = 14'h2dd9 == index ? 14'h82 : _GEN_11736;
  wire [13:0] _GEN_11738 = 14'h2dda == index ? 14'h81 : _GEN_11737;
  wire [13:0] _GEN_11739 = 14'h2ddb == index ? 14'h80 : _GEN_11738;
  wire [13:0] _GEN_11740 = 14'h2ddc == index ? 14'h5b : _GEN_11739;
  wire [13:0] _GEN_11741 = 14'h2ddd == index ? 14'h5b : _GEN_11740;
  wire [13:0] _GEN_11742 = 14'h2dde == index ? 14'h5b : _GEN_11741;
  wire [13:0] _GEN_11743 = 14'h2ddf == index ? 14'h5b : _GEN_11742;
  wire [13:0] _GEN_11744 = 14'h2de0 == index ? 14'h5b : _GEN_11743;
  wire [13:0] _GEN_11745 = 14'h2de1 == index ? 14'h5b : _GEN_11744;
  wire [13:0] _GEN_11746 = 14'h2de2 == index ? 14'h5b : _GEN_11745;
  wire [13:0] _GEN_11747 = 14'h2de3 == index ? 14'h5b : _GEN_11746;
  wire [13:0] _GEN_11748 = 14'h2de4 == index ? 14'h5b : _GEN_11747;
  wire [13:0] _GEN_11749 = 14'h2de5 == index ? 14'h5b : _GEN_11748;
  wire [13:0] _GEN_11750 = 14'h2de6 == index ? 14'h5b : _GEN_11749;
  wire [13:0] _GEN_11751 = 14'h2de7 == index ? 14'h5b : _GEN_11750;
  wire [13:0] _GEN_11752 = 14'h2de8 == index ? 14'h5b : _GEN_11751;
  wire [13:0] _GEN_11753 = 14'h2de9 == index ? 14'h5b : _GEN_11752;
  wire [13:0] _GEN_11754 = 14'h2dea == index ? 14'h5b : _GEN_11753;
  wire [13:0] _GEN_11755 = 14'h2deb == index ? 14'h5b : _GEN_11754;
  wire [13:0] _GEN_11756 = 14'h2dec == index ? 14'h5b : _GEN_11755;
  wire [13:0] _GEN_11757 = 14'h2ded == index ? 14'h5b : _GEN_11756;
  wire [13:0] _GEN_11758 = 14'h2dee == index ? 14'h5b : _GEN_11757;
  wire [13:0] _GEN_11759 = 14'h2def == index ? 14'h5b : _GEN_11758;
  wire [13:0] _GEN_11760 = 14'h2df0 == index ? 14'h5b : _GEN_11759;
  wire [13:0] _GEN_11761 = 14'h2df1 == index ? 14'h5b : _GEN_11760;
  wire [13:0] _GEN_11762 = 14'h2df2 == index ? 14'h5b : _GEN_11761;
  wire [13:0] _GEN_11763 = 14'h2df3 == index ? 14'h5b : _GEN_11762;
  wire [13:0] _GEN_11764 = 14'h2df4 == index ? 14'h5b : _GEN_11763;
  wire [13:0] _GEN_11765 = 14'h2df5 == index ? 14'h5b : _GEN_11764;
  wire [13:0] _GEN_11766 = 14'h2df6 == index ? 14'h5b : _GEN_11765;
  wire [13:0] _GEN_11767 = 14'h2df7 == index ? 14'h5b : _GEN_11766;
  wire [13:0] _GEN_11768 = 14'h2df8 == index ? 14'h5b : _GEN_11767;
  wire [13:0] _GEN_11769 = 14'h2df9 == index ? 14'h5b : _GEN_11768;
  wire [13:0] _GEN_11770 = 14'h2dfa == index ? 14'h5b : _GEN_11769;
  wire [13:0] _GEN_11771 = 14'h2dfb == index ? 14'h5b : _GEN_11770;
  wire [13:0] _GEN_11772 = 14'h2dfc == index ? 14'h5b : _GEN_11771;
  wire [13:0] _GEN_11773 = 14'h2dfd == index ? 14'h5b : _GEN_11772;
  wire [13:0] _GEN_11774 = 14'h2dfe == index ? 14'h5b : _GEN_11773;
  wire [13:0] _GEN_11775 = 14'h2dff == index ? 14'h5b : _GEN_11774;
  wire [13:0] _GEN_11776 = 14'h2e00 == index ? 14'h0 : _GEN_11775;
  wire [13:0] _GEN_11777 = 14'h2e01 == index ? 14'h2e00 : _GEN_11776;
  wire [13:0] _GEN_11778 = 14'h2e02 == index ? 14'h1700 : _GEN_11777;
  wire [13:0] _GEN_11779 = 14'h2e03 == index ? 14'hf02 : _GEN_11778;
  wire [13:0] _GEN_11780 = 14'h2e04 == index ? 14'hb80 : _GEN_11779;
  wire [13:0] _GEN_11781 = 14'h2e05 == index ? 14'h902 : _GEN_11780;
  wire [13:0] _GEN_11782 = 14'h2e06 == index ? 14'h782 : _GEN_11781;
  wire [13:0] _GEN_11783 = 14'h2e07 == index ? 14'h681 : _GEN_11782;
  wire [13:0] _GEN_11784 = 14'h2e08 == index ? 14'h584 : _GEN_11783;
  wire [13:0] _GEN_11785 = 14'h2e09 == index ? 14'h502 : _GEN_11784;
  wire [13:0] _GEN_11786 = 14'h2e0a == index ? 14'h482 : _GEN_11785;
  wire [13:0] _GEN_11787 = 14'h2e0b == index ? 14'h404 : _GEN_11786;
  wire [13:0] _GEN_11788 = 14'h2e0c == index ? 14'h388 : _GEN_11787;
  wire [13:0] _GEN_11789 = 14'h2e0d == index ? 14'h381 : _GEN_11788;
  wire [13:0] _GEN_11790 = 14'h2e0e == index ? 14'h308 : _GEN_11789;
  wire [13:0] _GEN_11791 = 14'h2e0f == index ? 14'h302 : _GEN_11790;
  wire [13:0] _GEN_11792 = 14'h2e10 == index ? 14'h28c : _GEN_11791;
  wire [13:0] _GEN_11793 = 14'h2e11 == index ? 14'h287 : _GEN_11792;
  wire [13:0] _GEN_11794 = 14'h2e12 == index ? 14'h282 : _GEN_11793;
  wire [13:0] _GEN_11795 = 14'h2e13 == index ? 14'h210 : _GEN_11794;
  wire [13:0] _GEN_11796 = 14'h2e14 == index ? 14'h20c : _GEN_11795;
  wire [13:0] _GEN_11797 = 14'h2e15 == index ? 14'h208 : _GEN_11796;
  wire [13:0] _GEN_11798 = 14'h2e16 == index ? 14'h204 : _GEN_11797;
  wire [13:0] _GEN_11799 = 14'h2e17 == index ? 14'h200 : _GEN_11798;
  wire [13:0] _GEN_11800 = 14'h2e18 == index ? 14'h194 : _GEN_11799;
  wire [13:0] _GEN_11801 = 14'h2e19 == index ? 14'h191 : _GEN_11800;
  wire [13:0] _GEN_11802 = 14'h2e1a == index ? 14'h18e : _GEN_11801;
  wire [13:0] _GEN_11803 = 14'h2e1b == index ? 14'h18b : _GEN_11802;
  wire [13:0] _GEN_11804 = 14'h2e1c == index ? 14'h188 : _GEN_11803;
  wire [13:0] _GEN_11805 = 14'h2e1d == index ? 14'h185 : _GEN_11804;
  wire [13:0] _GEN_11806 = 14'h2e1e == index ? 14'h182 : _GEN_11805;
  wire [13:0] _GEN_11807 = 14'h2e1f == index ? 14'h11e : _GEN_11806;
  wire [13:0] _GEN_11808 = 14'h2e20 == index ? 14'h11c : _GEN_11807;
  wire [13:0] _GEN_11809 = 14'h2e21 == index ? 14'h11a : _GEN_11808;
  wire [13:0] _GEN_11810 = 14'h2e22 == index ? 14'h118 : _GEN_11809;
  wire [13:0] _GEN_11811 = 14'h2e23 == index ? 14'h116 : _GEN_11810;
  wire [13:0] _GEN_11812 = 14'h2e24 == index ? 14'h114 : _GEN_11811;
  wire [13:0] _GEN_11813 = 14'h2e25 == index ? 14'h112 : _GEN_11812;
  wire [13:0] _GEN_11814 = 14'h2e26 == index ? 14'h110 : _GEN_11813;
  wire [13:0] _GEN_11815 = 14'h2e27 == index ? 14'h10e : _GEN_11814;
  wire [13:0] _GEN_11816 = 14'h2e28 == index ? 14'h10c : _GEN_11815;
  wire [13:0] _GEN_11817 = 14'h2e29 == index ? 14'h10a : _GEN_11816;
  wire [13:0] _GEN_11818 = 14'h2e2a == index ? 14'h108 : _GEN_11817;
  wire [13:0] _GEN_11819 = 14'h2e2b == index ? 14'h106 : _GEN_11818;
  wire [13:0] _GEN_11820 = 14'h2e2c == index ? 14'h104 : _GEN_11819;
  wire [13:0] _GEN_11821 = 14'h2e2d == index ? 14'h102 : _GEN_11820;
  wire [13:0] _GEN_11822 = 14'h2e2e == index ? 14'h100 : _GEN_11821;
  wire [13:0] _GEN_11823 = 14'h2e2f == index ? 14'had : _GEN_11822;
  wire [13:0] _GEN_11824 = 14'h2e30 == index ? 14'hac : _GEN_11823;
  wire [13:0] _GEN_11825 = 14'h2e31 == index ? 14'hab : _GEN_11824;
  wire [13:0] _GEN_11826 = 14'h2e32 == index ? 14'haa : _GEN_11825;
  wire [13:0] _GEN_11827 = 14'h2e33 == index ? 14'ha9 : _GEN_11826;
  wire [13:0] _GEN_11828 = 14'h2e34 == index ? 14'ha8 : _GEN_11827;
  wire [13:0] _GEN_11829 = 14'h2e35 == index ? 14'ha7 : _GEN_11828;
  wire [13:0] _GEN_11830 = 14'h2e36 == index ? 14'ha6 : _GEN_11829;
  wire [13:0] _GEN_11831 = 14'h2e37 == index ? 14'ha5 : _GEN_11830;
  wire [13:0] _GEN_11832 = 14'h2e38 == index ? 14'ha4 : _GEN_11831;
  wire [13:0] _GEN_11833 = 14'h2e39 == index ? 14'ha3 : _GEN_11832;
  wire [13:0] _GEN_11834 = 14'h2e3a == index ? 14'ha2 : _GEN_11833;
  wire [13:0] _GEN_11835 = 14'h2e3b == index ? 14'ha1 : _GEN_11834;
  wire [13:0] _GEN_11836 = 14'h2e3c == index ? 14'ha0 : _GEN_11835;
  wire [13:0] _GEN_11837 = 14'h2e3d == index ? 14'h9f : _GEN_11836;
  wire [13:0] _GEN_11838 = 14'h2e3e == index ? 14'h9e : _GEN_11837;
  wire [13:0] _GEN_11839 = 14'h2e3f == index ? 14'h9d : _GEN_11838;
  wire [13:0] _GEN_11840 = 14'h2e40 == index ? 14'h9c : _GEN_11839;
  wire [13:0] _GEN_11841 = 14'h2e41 == index ? 14'h9b : _GEN_11840;
  wire [13:0] _GEN_11842 = 14'h2e42 == index ? 14'h9a : _GEN_11841;
  wire [13:0] _GEN_11843 = 14'h2e43 == index ? 14'h99 : _GEN_11842;
  wire [13:0] _GEN_11844 = 14'h2e44 == index ? 14'h98 : _GEN_11843;
  wire [13:0] _GEN_11845 = 14'h2e45 == index ? 14'h97 : _GEN_11844;
  wire [13:0] _GEN_11846 = 14'h2e46 == index ? 14'h96 : _GEN_11845;
  wire [13:0] _GEN_11847 = 14'h2e47 == index ? 14'h95 : _GEN_11846;
  wire [13:0] _GEN_11848 = 14'h2e48 == index ? 14'h94 : _GEN_11847;
  wire [13:0] _GEN_11849 = 14'h2e49 == index ? 14'h93 : _GEN_11848;
  wire [13:0] _GEN_11850 = 14'h2e4a == index ? 14'h92 : _GEN_11849;
  wire [13:0] _GEN_11851 = 14'h2e4b == index ? 14'h91 : _GEN_11850;
  wire [13:0] _GEN_11852 = 14'h2e4c == index ? 14'h90 : _GEN_11851;
  wire [13:0] _GEN_11853 = 14'h2e4d == index ? 14'h8f : _GEN_11852;
  wire [13:0] _GEN_11854 = 14'h2e4e == index ? 14'h8e : _GEN_11853;
  wire [13:0] _GEN_11855 = 14'h2e4f == index ? 14'h8d : _GEN_11854;
  wire [13:0] _GEN_11856 = 14'h2e50 == index ? 14'h8c : _GEN_11855;
  wire [13:0] _GEN_11857 = 14'h2e51 == index ? 14'h8b : _GEN_11856;
  wire [13:0] _GEN_11858 = 14'h2e52 == index ? 14'h8a : _GEN_11857;
  wire [13:0] _GEN_11859 = 14'h2e53 == index ? 14'h89 : _GEN_11858;
  wire [13:0] _GEN_11860 = 14'h2e54 == index ? 14'h88 : _GEN_11859;
  wire [13:0] _GEN_11861 = 14'h2e55 == index ? 14'h87 : _GEN_11860;
  wire [13:0] _GEN_11862 = 14'h2e56 == index ? 14'h86 : _GEN_11861;
  wire [13:0] _GEN_11863 = 14'h2e57 == index ? 14'h85 : _GEN_11862;
  wire [13:0] _GEN_11864 = 14'h2e58 == index ? 14'h84 : _GEN_11863;
  wire [13:0] _GEN_11865 = 14'h2e59 == index ? 14'h83 : _GEN_11864;
  wire [13:0] _GEN_11866 = 14'h2e5a == index ? 14'h82 : _GEN_11865;
  wire [13:0] _GEN_11867 = 14'h2e5b == index ? 14'h81 : _GEN_11866;
  wire [13:0] _GEN_11868 = 14'h2e5c == index ? 14'h80 : _GEN_11867;
  wire [13:0] _GEN_11869 = 14'h2e5d == index ? 14'h5c : _GEN_11868;
  wire [13:0] _GEN_11870 = 14'h2e5e == index ? 14'h5c : _GEN_11869;
  wire [13:0] _GEN_11871 = 14'h2e5f == index ? 14'h5c : _GEN_11870;
  wire [13:0] _GEN_11872 = 14'h2e60 == index ? 14'h5c : _GEN_11871;
  wire [13:0] _GEN_11873 = 14'h2e61 == index ? 14'h5c : _GEN_11872;
  wire [13:0] _GEN_11874 = 14'h2e62 == index ? 14'h5c : _GEN_11873;
  wire [13:0] _GEN_11875 = 14'h2e63 == index ? 14'h5c : _GEN_11874;
  wire [13:0] _GEN_11876 = 14'h2e64 == index ? 14'h5c : _GEN_11875;
  wire [13:0] _GEN_11877 = 14'h2e65 == index ? 14'h5c : _GEN_11876;
  wire [13:0] _GEN_11878 = 14'h2e66 == index ? 14'h5c : _GEN_11877;
  wire [13:0] _GEN_11879 = 14'h2e67 == index ? 14'h5c : _GEN_11878;
  wire [13:0] _GEN_11880 = 14'h2e68 == index ? 14'h5c : _GEN_11879;
  wire [13:0] _GEN_11881 = 14'h2e69 == index ? 14'h5c : _GEN_11880;
  wire [13:0] _GEN_11882 = 14'h2e6a == index ? 14'h5c : _GEN_11881;
  wire [13:0] _GEN_11883 = 14'h2e6b == index ? 14'h5c : _GEN_11882;
  wire [13:0] _GEN_11884 = 14'h2e6c == index ? 14'h5c : _GEN_11883;
  wire [13:0] _GEN_11885 = 14'h2e6d == index ? 14'h5c : _GEN_11884;
  wire [13:0] _GEN_11886 = 14'h2e6e == index ? 14'h5c : _GEN_11885;
  wire [13:0] _GEN_11887 = 14'h2e6f == index ? 14'h5c : _GEN_11886;
  wire [13:0] _GEN_11888 = 14'h2e70 == index ? 14'h5c : _GEN_11887;
  wire [13:0] _GEN_11889 = 14'h2e71 == index ? 14'h5c : _GEN_11888;
  wire [13:0] _GEN_11890 = 14'h2e72 == index ? 14'h5c : _GEN_11889;
  wire [13:0] _GEN_11891 = 14'h2e73 == index ? 14'h5c : _GEN_11890;
  wire [13:0] _GEN_11892 = 14'h2e74 == index ? 14'h5c : _GEN_11891;
  wire [13:0] _GEN_11893 = 14'h2e75 == index ? 14'h5c : _GEN_11892;
  wire [13:0] _GEN_11894 = 14'h2e76 == index ? 14'h5c : _GEN_11893;
  wire [13:0] _GEN_11895 = 14'h2e77 == index ? 14'h5c : _GEN_11894;
  wire [13:0] _GEN_11896 = 14'h2e78 == index ? 14'h5c : _GEN_11895;
  wire [13:0] _GEN_11897 = 14'h2e79 == index ? 14'h5c : _GEN_11896;
  wire [13:0] _GEN_11898 = 14'h2e7a == index ? 14'h5c : _GEN_11897;
  wire [13:0] _GEN_11899 = 14'h2e7b == index ? 14'h5c : _GEN_11898;
  wire [13:0] _GEN_11900 = 14'h2e7c == index ? 14'h5c : _GEN_11899;
  wire [13:0] _GEN_11901 = 14'h2e7d == index ? 14'h5c : _GEN_11900;
  wire [13:0] _GEN_11902 = 14'h2e7e == index ? 14'h5c : _GEN_11901;
  wire [13:0] _GEN_11903 = 14'h2e7f == index ? 14'h5c : _GEN_11902;
  wire [13:0] _GEN_11904 = 14'h2e80 == index ? 14'h0 : _GEN_11903;
  wire [13:0] _GEN_11905 = 14'h2e81 == index ? 14'h2e80 : _GEN_11904;
  wire [13:0] _GEN_11906 = 14'h2e82 == index ? 14'h1701 : _GEN_11905;
  wire [13:0] _GEN_11907 = 14'h2e83 == index ? 14'hf80 : _GEN_11906;
  wire [13:0] _GEN_11908 = 14'h2e84 == index ? 14'hb81 : _GEN_11907;
  wire [13:0] _GEN_11909 = 14'h2e85 == index ? 14'h903 : _GEN_11908;
  wire [13:0] _GEN_11910 = 14'h2e86 == index ? 14'h783 : _GEN_11909;
  wire [13:0] _GEN_11911 = 14'h2e87 == index ? 14'h682 : _GEN_11910;
  wire [13:0] _GEN_11912 = 14'h2e88 == index ? 14'h585 : _GEN_11911;
  wire [13:0] _GEN_11913 = 14'h2e89 == index ? 14'h503 : _GEN_11912;
  wire [13:0] _GEN_11914 = 14'h2e8a == index ? 14'h483 : _GEN_11913;
  wire [13:0] _GEN_11915 = 14'h2e8b == index ? 14'h405 : _GEN_11914;
  wire [13:0] _GEN_11916 = 14'h2e8c == index ? 14'h389 : _GEN_11915;
  wire [13:0] _GEN_11917 = 14'h2e8d == index ? 14'h382 : _GEN_11916;
  wire [13:0] _GEN_11918 = 14'h2e8e == index ? 14'h309 : _GEN_11917;
  wire [13:0] _GEN_11919 = 14'h2e8f == index ? 14'h303 : _GEN_11918;
  wire [13:0] _GEN_11920 = 14'h2e90 == index ? 14'h28d : _GEN_11919;
  wire [13:0] _GEN_11921 = 14'h2e91 == index ? 14'h288 : _GEN_11920;
  wire [13:0] _GEN_11922 = 14'h2e92 == index ? 14'h283 : _GEN_11921;
  wire [13:0] _GEN_11923 = 14'h2e93 == index ? 14'h211 : _GEN_11922;
  wire [13:0] _GEN_11924 = 14'h2e94 == index ? 14'h20d : _GEN_11923;
  wire [13:0] _GEN_11925 = 14'h2e95 == index ? 14'h209 : _GEN_11924;
  wire [13:0] _GEN_11926 = 14'h2e96 == index ? 14'h205 : _GEN_11925;
  wire [13:0] _GEN_11927 = 14'h2e97 == index ? 14'h201 : _GEN_11926;
  wire [13:0] _GEN_11928 = 14'h2e98 == index ? 14'h195 : _GEN_11927;
  wire [13:0] _GEN_11929 = 14'h2e99 == index ? 14'h192 : _GEN_11928;
  wire [13:0] _GEN_11930 = 14'h2e9a == index ? 14'h18f : _GEN_11929;
  wire [13:0] _GEN_11931 = 14'h2e9b == index ? 14'h18c : _GEN_11930;
  wire [13:0] _GEN_11932 = 14'h2e9c == index ? 14'h189 : _GEN_11931;
  wire [13:0] _GEN_11933 = 14'h2e9d == index ? 14'h186 : _GEN_11932;
  wire [13:0] _GEN_11934 = 14'h2e9e == index ? 14'h183 : _GEN_11933;
  wire [13:0] _GEN_11935 = 14'h2e9f == index ? 14'h180 : _GEN_11934;
  wire [13:0] _GEN_11936 = 14'h2ea0 == index ? 14'h11d : _GEN_11935;
  wire [13:0] _GEN_11937 = 14'h2ea1 == index ? 14'h11b : _GEN_11936;
  wire [13:0] _GEN_11938 = 14'h2ea2 == index ? 14'h119 : _GEN_11937;
  wire [13:0] _GEN_11939 = 14'h2ea3 == index ? 14'h117 : _GEN_11938;
  wire [13:0] _GEN_11940 = 14'h2ea4 == index ? 14'h115 : _GEN_11939;
  wire [13:0] _GEN_11941 = 14'h2ea5 == index ? 14'h113 : _GEN_11940;
  wire [13:0] _GEN_11942 = 14'h2ea6 == index ? 14'h111 : _GEN_11941;
  wire [13:0] _GEN_11943 = 14'h2ea7 == index ? 14'h10f : _GEN_11942;
  wire [13:0] _GEN_11944 = 14'h2ea8 == index ? 14'h10d : _GEN_11943;
  wire [13:0] _GEN_11945 = 14'h2ea9 == index ? 14'h10b : _GEN_11944;
  wire [13:0] _GEN_11946 = 14'h2eaa == index ? 14'h109 : _GEN_11945;
  wire [13:0] _GEN_11947 = 14'h2eab == index ? 14'h107 : _GEN_11946;
  wire [13:0] _GEN_11948 = 14'h2eac == index ? 14'h105 : _GEN_11947;
  wire [13:0] _GEN_11949 = 14'h2ead == index ? 14'h103 : _GEN_11948;
  wire [13:0] _GEN_11950 = 14'h2eae == index ? 14'h101 : _GEN_11949;
  wire [13:0] _GEN_11951 = 14'h2eaf == index ? 14'hae : _GEN_11950;
  wire [13:0] _GEN_11952 = 14'h2eb0 == index ? 14'had : _GEN_11951;
  wire [13:0] _GEN_11953 = 14'h2eb1 == index ? 14'hac : _GEN_11952;
  wire [13:0] _GEN_11954 = 14'h2eb2 == index ? 14'hab : _GEN_11953;
  wire [13:0] _GEN_11955 = 14'h2eb3 == index ? 14'haa : _GEN_11954;
  wire [13:0] _GEN_11956 = 14'h2eb4 == index ? 14'ha9 : _GEN_11955;
  wire [13:0] _GEN_11957 = 14'h2eb5 == index ? 14'ha8 : _GEN_11956;
  wire [13:0] _GEN_11958 = 14'h2eb6 == index ? 14'ha7 : _GEN_11957;
  wire [13:0] _GEN_11959 = 14'h2eb7 == index ? 14'ha6 : _GEN_11958;
  wire [13:0] _GEN_11960 = 14'h2eb8 == index ? 14'ha5 : _GEN_11959;
  wire [13:0] _GEN_11961 = 14'h2eb9 == index ? 14'ha4 : _GEN_11960;
  wire [13:0] _GEN_11962 = 14'h2eba == index ? 14'ha3 : _GEN_11961;
  wire [13:0] _GEN_11963 = 14'h2ebb == index ? 14'ha2 : _GEN_11962;
  wire [13:0] _GEN_11964 = 14'h2ebc == index ? 14'ha1 : _GEN_11963;
  wire [13:0] _GEN_11965 = 14'h2ebd == index ? 14'ha0 : _GEN_11964;
  wire [13:0] _GEN_11966 = 14'h2ebe == index ? 14'h9f : _GEN_11965;
  wire [13:0] _GEN_11967 = 14'h2ebf == index ? 14'h9e : _GEN_11966;
  wire [13:0] _GEN_11968 = 14'h2ec0 == index ? 14'h9d : _GEN_11967;
  wire [13:0] _GEN_11969 = 14'h2ec1 == index ? 14'h9c : _GEN_11968;
  wire [13:0] _GEN_11970 = 14'h2ec2 == index ? 14'h9b : _GEN_11969;
  wire [13:0] _GEN_11971 = 14'h2ec3 == index ? 14'h9a : _GEN_11970;
  wire [13:0] _GEN_11972 = 14'h2ec4 == index ? 14'h99 : _GEN_11971;
  wire [13:0] _GEN_11973 = 14'h2ec5 == index ? 14'h98 : _GEN_11972;
  wire [13:0] _GEN_11974 = 14'h2ec6 == index ? 14'h97 : _GEN_11973;
  wire [13:0] _GEN_11975 = 14'h2ec7 == index ? 14'h96 : _GEN_11974;
  wire [13:0] _GEN_11976 = 14'h2ec8 == index ? 14'h95 : _GEN_11975;
  wire [13:0] _GEN_11977 = 14'h2ec9 == index ? 14'h94 : _GEN_11976;
  wire [13:0] _GEN_11978 = 14'h2eca == index ? 14'h93 : _GEN_11977;
  wire [13:0] _GEN_11979 = 14'h2ecb == index ? 14'h92 : _GEN_11978;
  wire [13:0] _GEN_11980 = 14'h2ecc == index ? 14'h91 : _GEN_11979;
  wire [13:0] _GEN_11981 = 14'h2ecd == index ? 14'h90 : _GEN_11980;
  wire [13:0] _GEN_11982 = 14'h2ece == index ? 14'h8f : _GEN_11981;
  wire [13:0] _GEN_11983 = 14'h2ecf == index ? 14'h8e : _GEN_11982;
  wire [13:0] _GEN_11984 = 14'h2ed0 == index ? 14'h8d : _GEN_11983;
  wire [13:0] _GEN_11985 = 14'h2ed1 == index ? 14'h8c : _GEN_11984;
  wire [13:0] _GEN_11986 = 14'h2ed2 == index ? 14'h8b : _GEN_11985;
  wire [13:0] _GEN_11987 = 14'h2ed3 == index ? 14'h8a : _GEN_11986;
  wire [13:0] _GEN_11988 = 14'h2ed4 == index ? 14'h89 : _GEN_11987;
  wire [13:0] _GEN_11989 = 14'h2ed5 == index ? 14'h88 : _GEN_11988;
  wire [13:0] _GEN_11990 = 14'h2ed6 == index ? 14'h87 : _GEN_11989;
  wire [13:0] _GEN_11991 = 14'h2ed7 == index ? 14'h86 : _GEN_11990;
  wire [13:0] _GEN_11992 = 14'h2ed8 == index ? 14'h85 : _GEN_11991;
  wire [13:0] _GEN_11993 = 14'h2ed9 == index ? 14'h84 : _GEN_11992;
  wire [13:0] _GEN_11994 = 14'h2eda == index ? 14'h83 : _GEN_11993;
  wire [13:0] _GEN_11995 = 14'h2edb == index ? 14'h82 : _GEN_11994;
  wire [13:0] _GEN_11996 = 14'h2edc == index ? 14'h81 : _GEN_11995;
  wire [13:0] _GEN_11997 = 14'h2edd == index ? 14'h80 : _GEN_11996;
  wire [13:0] _GEN_11998 = 14'h2ede == index ? 14'h5d : _GEN_11997;
  wire [13:0] _GEN_11999 = 14'h2edf == index ? 14'h5d : _GEN_11998;
  wire [13:0] _GEN_12000 = 14'h2ee0 == index ? 14'h5d : _GEN_11999;
  wire [13:0] _GEN_12001 = 14'h2ee1 == index ? 14'h5d : _GEN_12000;
  wire [13:0] _GEN_12002 = 14'h2ee2 == index ? 14'h5d : _GEN_12001;
  wire [13:0] _GEN_12003 = 14'h2ee3 == index ? 14'h5d : _GEN_12002;
  wire [13:0] _GEN_12004 = 14'h2ee4 == index ? 14'h5d : _GEN_12003;
  wire [13:0] _GEN_12005 = 14'h2ee5 == index ? 14'h5d : _GEN_12004;
  wire [13:0] _GEN_12006 = 14'h2ee6 == index ? 14'h5d : _GEN_12005;
  wire [13:0] _GEN_12007 = 14'h2ee7 == index ? 14'h5d : _GEN_12006;
  wire [13:0] _GEN_12008 = 14'h2ee8 == index ? 14'h5d : _GEN_12007;
  wire [13:0] _GEN_12009 = 14'h2ee9 == index ? 14'h5d : _GEN_12008;
  wire [13:0] _GEN_12010 = 14'h2eea == index ? 14'h5d : _GEN_12009;
  wire [13:0] _GEN_12011 = 14'h2eeb == index ? 14'h5d : _GEN_12010;
  wire [13:0] _GEN_12012 = 14'h2eec == index ? 14'h5d : _GEN_12011;
  wire [13:0] _GEN_12013 = 14'h2eed == index ? 14'h5d : _GEN_12012;
  wire [13:0] _GEN_12014 = 14'h2eee == index ? 14'h5d : _GEN_12013;
  wire [13:0] _GEN_12015 = 14'h2eef == index ? 14'h5d : _GEN_12014;
  wire [13:0] _GEN_12016 = 14'h2ef0 == index ? 14'h5d : _GEN_12015;
  wire [13:0] _GEN_12017 = 14'h2ef1 == index ? 14'h5d : _GEN_12016;
  wire [13:0] _GEN_12018 = 14'h2ef2 == index ? 14'h5d : _GEN_12017;
  wire [13:0] _GEN_12019 = 14'h2ef3 == index ? 14'h5d : _GEN_12018;
  wire [13:0] _GEN_12020 = 14'h2ef4 == index ? 14'h5d : _GEN_12019;
  wire [13:0] _GEN_12021 = 14'h2ef5 == index ? 14'h5d : _GEN_12020;
  wire [13:0] _GEN_12022 = 14'h2ef6 == index ? 14'h5d : _GEN_12021;
  wire [13:0] _GEN_12023 = 14'h2ef7 == index ? 14'h5d : _GEN_12022;
  wire [13:0] _GEN_12024 = 14'h2ef8 == index ? 14'h5d : _GEN_12023;
  wire [13:0] _GEN_12025 = 14'h2ef9 == index ? 14'h5d : _GEN_12024;
  wire [13:0] _GEN_12026 = 14'h2efa == index ? 14'h5d : _GEN_12025;
  wire [13:0] _GEN_12027 = 14'h2efb == index ? 14'h5d : _GEN_12026;
  wire [13:0] _GEN_12028 = 14'h2efc == index ? 14'h5d : _GEN_12027;
  wire [13:0] _GEN_12029 = 14'h2efd == index ? 14'h5d : _GEN_12028;
  wire [13:0] _GEN_12030 = 14'h2efe == index ? 14'h5d : _GEN_12029;
  wire [13:0] _GEN_12031 = 14'h2eff == index ? 14'h5d : _GEN_12030;
  wire [13:0] _GEN_12032 = 14'h2f00 == index ? 14'h0 : _GEN_12031;
  wire [13:0] _GEN_12033 = 14'h2f01 == index ? 14'h2f00 : _GEN_12032;
  wire [13:0] _GEN_12034 = 14'h2f02 == index ? 14'h1780 : _GEN_12033;
  wire [13:0] _GEN_12035 = 14'h2f03 == index ? 14'hf81 : _GEN_12034;
  wire [13:0] _GEN_12036 = 14'h2f04 == index ? 14'hb82 : _GEN_12035;
  wire [13:0] _GEN_12037 = 14'h2f05 == index ? 14'h904 : _GEN_12036;
  wire [13:0] _GEN_12038 = 14'h2f06 == index ? 14'h784 : _GEN_12037;
  wire [13:0] _GEN_12039 = 14'h2f07 == index ? 14'h683 : _GEN_12038;
  wire [13:0] _GEN_12040 = 14'h2f08 == index ? 14'h586 : _GEN_12039;
  wire [13:0] _GEN_12041 = 14'h2f09 == index ? 14'h504 : _GEN_12040;
  wire [13:0] _GEN_12042 = 14'h2f0a == index ? 14'h484 : _GEN_12041;
  wire [13:0] _GEN_12043 = 14'h2f0b == index ? 14'h406 : _GEN_12042;
  wire [13:0] _GEN_12044 = 14'h2f0c == index ? 14'h38a : _GEN_12043;
  wire [13:0] _GEN_12045 = 14'h2f0d == index ? 14'h383 : _GEN_12044;
  wire [13:0] _GEN_12046 = 14'h2f0e == index ? 14'h30a : _GEN_12045;
  wire [13:0] _GEN_12047 = 14'h2f0f == index ? 14'h304 : _GEN_12046;
  wire [13:0] _GEN_12048 = 14'h2f10 == index ? 14'h28e : _GEN_12047;
  wire [13:0] _GEN_12049 = 14'h2f11 == index ? 14'h289 : _GEN_12048;
  wire [13:0] _GEN_12050 = 14'h2f12 == index ? 14'h284 : _GEN_12049;
  wire [13:0] _GEN_12051 = 14'h2f13 == index ? 14'h212 : _GEN_12050;
  wire [13:0] _GEN_12052 = 14'h2f14 == index ? 14'h20e : _GEN_12051;
  wire [13:0] _GEN_12053 = 14'h2f15 == index ? 14'h20a : _GEN_12052;
  wire [13:0] _GEN_12054 = 14'h2f16 == index ? 14'h206 : _GEN_12053;
  wire [13:0] _GEN_12055 = 14'h2f17 == index ? 14'h202 : _GEN_12054;
  wire [13:0] _GEN_12056 = 14'h2f18 == index ? 14'h196 : _GEN_12055;
  wire [13:0] _GEN_12057 = 14'h2f19 == index ? 14'h193 : _GEN_12056;
  wire [13:0] _GEN_12058 = 14'h2f1a == index ? 14'h190 : _GEN_12057;
  wire [13:0] _GEN_12059 = 14'h2f1b == index ? 14'h18d : _GEN_12058;
  wire [13:0] _GEN_12060 = 14'h2f1c == index ? 14'h18a : _GEN_12059;
  wire [13:0] _GEN_12061 = 14'h2f1d == index ? 14'h187 : _GEN_12060;
  wire [13:0] _GEN_12062 = 14'h2f1e == index ? 14'h184 : _GEN_12061;
  wire [13:0] _GEN_12063 = 14'h2f1f == index ? 14'h181 : _GEN_12062;
  wire [13:0] _GEN_12064 = 14'h2f20 == index ? 14'h11e : _GEN_12063;
  wire [13:0] _GEN_12065 = 14'h2f21 == index ? 14'h11c : _GEN_12064;
  wire [13:0] _GEN_12066 = 14'h2f22 == index ? 14'h11a : _GEN_12065;
  wire [13:0] _GEN_12067 = 14'h2f23 == index ? 14'h118 : _GEN_12066;
  wire [13:0] _GEN_12068 = 14'h2f24 == index ? 14'h116 : _GEN_12067;
  wire [13:0] _GEN_12069 = 14'h2f25 == index ? 14'h114 : _GEN_12068;
  wire [13:0] _GEN_12070 = 14'h2f26 == index ? 14'h112 : _GEN_12069;
  wire [13:0] _GEN_12071 = 14'h2f27 == index ? 14'h110 : _GEN_12070;
  wire [13:0] _GEN_12072 = 14'h2f28 == index ? 14'h10e : _GEN_12071;
  wire [13:0] _GEN_12073 = 14'h2f29 == index ? 14'h10c : _GEN_12072;
  wire [13:0] _GEN_12074 = 14'h2f2a == index ? 14'h10a : _GEN_12073;
  wire [13:0] _GEN_12075 = 14'h2f2b == index ? 14'h108 : _GEN_12074;
  wire [13:0] _GEN_12076 = 14'h2f2c == index ? 14'h106 : _GEN_12075;
  wire [13:0] _GEN_12077 = 14'h2f2d == index ? 14'h104 : _GEN_12076;
  wire [13:0] _GEN_12078 = 14'h2f2e == index ? 14'h102 : _GEN_12077;
  wire [13:0] _GEN_12079 = 14'h2f2f == index ? 14'h100 : _GEN_12078;
  wire [13:0] _GEN_12080 = 14'h2f30 == index ? 14'hae : _GEN_12079;
  wire [13:0] _GEN_12081 = 14'h2f31 == index ? 14'had : _GEN_12080;
  wire [13:0] _GEN_12082 = 14'h2f32 == index ? 14'hac : _GEN_12081;
  wire [13:0] _GEN_12083 = 14'h2f33 == index ? 14'hab : _GEN_12082;
  wire [13:0] _GEN_12084 = 14'h2f34 == index ? 14'haa : _GEN_12083;
  wire [13:0] _GEN_12085 = 14'h2f35 == index ? 14'ha9 : _GEN_12084;
  wire [13:0] _GEN_12086 = 14'h2f36 == index ? 14'ha8 : _GEN_12085;
  wire [13:0] _GEN_12087 = 14'h2f37 == index ? 14'ha7 : _GEN_12086;
  wire [13:0] _GEN_12088 = 14'h2f38 == index ? 14'ha6 : _GEN_12087;
  wire [13:0] _GEN_12089 = 14'h2f39 == index ? 14'ha5 : _GEN_12088;
  wire [13:0] _GEN_12090 = 14'h2f3a == index ? 14'ha4 : _GEN_12089;
  wire [13:0] _GEN_12091 = 14'h2f3b == index ? 14'ha3 : _GEN_12090;
  wire [13:0] _GEN_12092 = 14'h2f3c == index ? 14'ha2 : _GEN_12091;
  wire [13:0] _GEN_12093 = 14'h2f3d == index ? 14'ha1 : _GEN_12092;
  wire [13:0] _GEN_12094 = 14'h2f3e == index ? 14'ha0 : _GEN_12093;
  wire [13:0] _GEN_12095 = 14'h2f3f == index ? 14'h9f : _GEN_12094;
  wire [13:0] _GEN_12096 = 14'h2f40 == index ? 14'h9e : _GEN_12095;
  wire [13:0] _GEN_12097 = 14'h2f41 == index ? 14'h9d : _GEN_12096;
  wire [13:0] _GEN_12098 = 14'h2f42 == index ? 14'h9c : _GEN_12097;
  wire [13:0] _GEN_12099 = 14'h2f43 == index ? 14'h9b : _GEN_12098;
  wire [13:0] _GEN_12100 = 14'h2f44 == index ? 14'h9a : _GEN_12099;
  wire [13:0] _GEN_12101 = 14'h2f45 == index ? 14'h99 : _GEN_12100;
  wire [13:0] _GEN_12102 = 14'h2f46 == index ? 14'h98 : _GEN_12101;
  wire [13:0] _GEN_12103 = 14'h2f47 == index ? 14'h97 : _GEN_12102;
  wire [13:0] _GEN_12104 = 14'h2f48 == index ? 14'h96 : _GEN_12103;
  wire [13:0] _GEN_12105 = 14'h2f49 == index ? 14'h95 : _GEN_12104;
  wire [13:0] _GEN_12106 = 14'h2f4a == index ? 14'h94 : _GEN_12105;
  wire [13:0] _GEN_12107 = 14'h2f4b == index ? 14'h93 : _GEN_12106;
  wire [13:0] _GEN_12108 = 14'h2f4c == index ? 14'h92 : _GEN_12107;
  wire [13:0] _GEN_12109 = 14'h2f4d == index ? 14'h91 : _GEN_12108;
  wire [13:0] _GEN_12110 = 14'h2f4e == index ? 14'h90 : _GEN_12109;
  wire [13:0] _GEN_12111 = 14'h2f4f == index ? 14'h8f : _GEN_12110;
  wire [13:0] _GEN_12112 = 14'h2f50 == index ? 14'h8e : _GEN_12111;
  wire [13:0] _GEN_12113 = 14'h2f51 == index ? 14'h8d : _GEN_12112;
  wire [13:0] _GEN_12114 = 14'h2f52 == index ? 14'h8c : _GEN_12113;
  wire [13:0] _GEN_12115 = 14'h2f53 == index ? 14'h8b : _GEN_12114;
  wire [13:0] _GEN_12116 = 14'h2f54 == index ? 14'h8a : _GEN_12115;
  wire [13:0] _GEN_12117 = 14'h2f55 == index ? 14'h89 : _GEN_12116;
  wire [13:0] _GEN_12118 = 14'h2f56 == index ? 14'h88 : _GEN_12117;
  wire [13:0] _GEN_12119 = 14'h2f57 == index ? 14'h87 : _GEN_12118;
  wire [13:0] _GEN_12120 = 14'h2f58 == index ? 14'h86 : _GEN_12119;
  wire [13:0] _GEN_12121 = 14'h2f59 == index ? 14'h85 : _GEN_12120;
  wire [13:0] _GEN_12122 = 14'h2f5a == index ? 14'h84 : _GEN_12121;
  wire [13:0] _GEN_12123 = 14'h2f5b == index ? 14'h83 : _GEN_12122;
  wire [13:0] _GEN_12124 = 14'h2f5c == index ? 14'h82 : _GEN_12123;
  wire [13:0] _GEN_12125 = 14'h2f5d == index ? 14'h81 : _GEN_12124;
  wire [13:0] _GEN_12126 = 14'h2f5e == index ? 14'h80 : _GEN_12125;
  wire [13:0] _GEN_12127 = 14'h2f5f == index ? 14'h5e : _GEN_12126;
  wire [13:0] _GEN_12128 = 14'h2f60 == index ? 14'h5e : _GEN_12127;
  wire [13:0] _GEN_12129 = 14'h2f61 == index ? 14'h5e : _GEN_12128;
  wire [13:0] _GEN_12130 = 14'h2f62 == index ? 14'h5e : _GEN_12129;
  wire [13:0] _GEN_12131 = 14'h2f63 == index ? 14'h5e : _GEN_12130;
  wire [13:0] _GEN_12132 = 14'h2f64 == index ? 14'h5e : _GEN_12131;
  wire [13:0] _GEN_12133 = 14'h2f65 == index ? 14'h5e : _GEN_12132;
  wire [13:0] _GEN_12134 = 14'h2f66 == index ? 14'h5e : _GEN_12133;
  wire [13:0] _GEN_12135 = 14'h2f67 == index ? 14'h5e : _GEN_12134;
  wire [13:0] _GEN_12136 = 14'h2f68 == index ? 14'h5e : _GEN_12135;
  wire [13:0] _GEN_12137 = 14'h2f69 == index ? 14'h5e : _GEN_12136;
  wire [13:0] _GEN_12138 = 14'h2f6a == index ? 14'h5e : _GEN_12137;
  wire [13:0] _GEN_12139 = 14'h2f6b == index ? 14'h5e : _GEN_12138;
  wire [13:0] _GEN_12140 = 14'h2f6c == index ? 14'h5e : _GEN_12139;
  wire [13:0] _GEN_12141 = 14'h2f6d == index ? 14'h5e : _GEN_12140;
  wire [13:0] _GEN_12142 = 14'h2f6e == index ? 14'h5e : _GEN_12141;
  wire [13:0] _GEN_12143 = 14'h2f6f == index ? 14'h5e : _GEN_12142;
  wire [13:0] _GEN_12144 = 14'h2f70 == index ? 14'h5e : _GEN_12143;
  wire [13:0] _GEN_12145 = 14'h2f71 == index ? 14'h5e : _GEN_12144;
  wire [13:0] _GEN_12146 = 14'h2f72 == index ? 14'h5e : _GEN_12145;
  wire [13:0] _GEN_12147 = 14'h2f73 == index ? 14'h5e : _GEN_12146;
  wire [13:0] _GEN_12148 = 14'h2f74 == index ? 14'h5e : _GEN_12147;
  wire [13:0] _GEN_12149 = 14'h2f75 == index ? 14'h5e : _GEN_12148;
  wire [13:0] _GEN_12150 = 14'h2f76 == index ? 14'h5e : _GEN_12149;
  wire [13:0] _GEN_12151 = 14'h2f77 == index ? 14'h5e : _GEN_12150;
  wire [13:0] _GEN_12152 = 14'h2f78 == index ? 14'h5e : _GEN_12151;
  wire [13:0] _GEN_12153 = 14'h2f79 == index ? 14'h5e : _GEN_12152;
  wire [13:0] _GEN_12154 = 14'h2f7a == index ? 14'h5e : _GEN_12153;
  wire [13:0] _GEN_12155 = 14'h2f7b == index ? 14'h5e : _GEN_12154;
  wire [13:0] _GEN_12156 = 14'h2f7c == index ? 14'h5e : _GEN_12155;
  wire [13:0] _GEN_12157 = 14'h2f7d == index ? 14'h5e : _GEN_12156;
  wire [13:0] _GEN_12158 = 14'h2f7e == index ? 14'h5e : _GEN_12157;
  wire [13:0] _GEN_12159 = 14'h2f7f == index ? 14'h5e : _GEN_12158;
  wire [13:0] _GEN_12160 = 14'h2f80 == index ? 14'h0 : _GEN_12159;
  wire [13:0] _GEN_12161 = 14'h2f81 == index ? 14'h2f80 : _GEN_12160;
  wire [13:0] _GEN_12162 = 14'h2f82 == index ? 14'h1781 : _GEN_12161;
  wire [13:0] _GEN_12163 = 14'h2f83 == index ? 14'hf82 : _GEN_12162;
  wire [13:0] _GEN_12164 = 14'h2f84 == index ? 14'hb83 : _GEN_12163;
  wire [13:0] _GEN_12165 = 14'h2f85 == index ? 14'h980 : _GEN_12164;
  wire [13:0] _GEN_12166 = 14'h2f86 == index ? 14'h785 : _GEN_12165;
  wire [13:0] _GEN_12167 = 14'h2f87 == index ? 14'h684 : _GEN_12166;
  wire [13:0] _GEN_12168 = 14'h2f88 == index ? 14'h587 : _GEN_12167;
  wire [13:0] _GEN_12169 = 14'h2f89 == index ? 14'h505 : _GEN_12168;
  wire [13:0] _GEN_12170 = 14'h2f8a == index ? 14'h485 : _GEN_12169;
  wire [13:0] _GEN_12171 = 14'h2f8b == index ? 14'h407 : _GEN_12170;
  wire [13:0] _GEN_12172 = 14'h2f8c == index ? 14'h38b : _GEN_12171;
  wire [13:0] _GEN_12173 = 14'h2f8d == index ? 14'h384 : _GEN_12172;
  wire [13:0] _GEN_12174 = 14'h2f8e == index ? 14'h30b : _GEN_12173;
  wire [13:0] _GEN_12175 = 14'h2f8f == index ? 14'h305 : _GEN_12174;
  wire [13:0] _GEN_12176 = 14'h2f90 == index ? 14'h28f : _GEN_12175;
  wire [13:0] _GEN_12177 = 14'h2f91 == index ? 14'h28a : _GEN_12176;
  wire [13:0] _GEN_12178 = 14'h2f92 == index ? 14'h285 : _GEN_12177;
  wire [13:0] _GEN_12179 = 14'h2f93 == index ? 14'h280 : _GEN_12178;
  wire [13:0] _GEN_12180 = 14'h2f94 == index ? 14'h20f : _GEN_12179;
  wire [13:0] _GEN_12181 = 14'h2f95 == index ? 14'h20b : _GEN_12180;
  wire [13:0] _GEN_12182 = 14'h2f96 == index ? 14'h207 : _GEN_12181;
  wire [13:0] _GEN_12183 = 14'h2f97 == index ? 14'h203 : _GEN_12182;
  wire [13:0] _GEN_12184 = 14'h2f98 == index ? 14'h197 : _GEN_12183;
  wire [13:0] _GEN_12185 = 14'h2f99 == index ? 14'h194 : _GEN_12184;
  wire [13:0] _GEN_12186 = 14'h2f9a == index ? 14'h191 : _GEN_12185;
  wire [13:0] _GEN_12187 = 14'h2f9b == index ? 14'h18e : _GEN_12186;
  wire [13:0] _GEN_12188 = 14'h2f9c == index ? 14'h18b : _GEN_12187;
  wire [13:0] _GEN_12189 = 14'h2f9d == index ? 14'h188 : _GEN_12188;
  wire [13:0] _GEN_12190 = 14'h2f9e == index ? 14'h185 : _GEN_12189;
  wire [13:0] _GEN_12191 = 14'h2f9f == index ? 14'h182 : _GEN_12190;
  wire [13:0] _GEN_12192 = 14'h2fa0 == index ? 14'h11f : _GEN_12191;
  wire [13:0] _GEN_12193 = 14'h2fa1 == index ? 14'h11d : _GEN_12192;
  wire [13:0] _GEN_12194 = 14'h2fa2 == index ? 14'h11b : _GEN_12193;
  wire [13:0] _GEN_12195 = 14'h2fa3 == index ? 14'h119 : _GEN_12194;
  wire [13:0] _GEN_12196 = 14'h2fa4 == index ? 14'h117 : _GEN_12195;
  wire [13:0] _GEN_12197 = 14'h2fa5 == index ? 14'h115 : _GEN_12196;
  wire [13:0] _GEN_12198 = 14'h2fa6 == index ? 14'h113 : _GEN_12197;
  wire [13:0] _GEN_12199 = 14'h2fa7 == index ? 14'h111 : _GEN_12198;
  wire [13:0] _GEN_12200 = 14'h2fa8 == index ? 14'h10f : _GEN_12199;
  wire [13:0] _GEN_12201 = 14'h2fa9 == index ? 14'h10d : _GEN_12200;
  wire [13:0] _GEN_12202 = 14'h2faa == index ? 14'h10b : _GEN_12201;
  wire [13:0] _GEN_12203 = 14'h2fab == index ? 14'h109 : _GEN_12202;
  wire [13:0] _GEN_12204 = 14'h2fac == index ? 14'h107 : _GEN_12203;
  wire [13:0] _GEN_12205 = 14'h2fad == index ? 14'h105 : _GEN_12204;
  wire [13:0] _GEN_12206 = 14'h2fae == index ? 14'h103 : _GEN_12205;
  wire [13:0] _GEN_12207 = 14'h2faf == index ? 14'h101 : _GEN_12206;
  wire [13:0] _GEN_12208 = 14'h2fb0 == index ? 14'haf : _GEN_12207;
  wire [13:0] _GEN_12209 = 14'h2fb1 == index ? 14'hae : _GEN_12208;
  wire [13:0] _GEN_12210 = 14'h2fb2 == index ? 14'had : _GEN_12209;
  wire [13:0] _GEN_12211 = 14'h2fb3 == index ? 14'hac : _GEN_12210;
  wire [13:0] _GEN_12212 = 14'h2fb4 == index ? 14'hab : _GEN_12211;
  wire [13:0] _GEN_12213 = 14'h2fb5 == index ? 14'haa : _GEN_12212;
  wire [13:0] _GEN_12214 = 14'h2fb6 == index ? 14'ha9 : _GEN_12213;
  wire [13:0] _GEN_12215 = 14'h2fb7 == index ? 14'ha8 : _GEN_12214;
  wire [13:0] _GEN_12216 = 14'h2fb8 == index ? 14'ha7 : _GEN_12215;
  wire [13:0] _GEN_12217 = 14'h2fb9 == index ? 14'ha6 : _GEN_12216;
  wire [13:0] _GEN_12218 = 14'h2fba == index ? 14'ha5 : _GEN_12217;
  wire [13:0] _GEN_12219 = 14'h2fbb == index ? 14'ha4 : _GEN_12218;
  wire [13:0] _GEN_12220 = 14'h2fbc == index ? 14'ha3 : _GEN_12219;
  wire [13:0] _GEN_12221 = 14'h2fbd == index ? 14'ha2 : _GEN_12220;
  wire [13:0] _GEN_12222 = 14'h2fbe == index ? 14'ha1 : _GEN_12221;
  wire [13:0] _GEN_12223 = 14'h2fbf == index ? 14'ha0 : _GEN_12222;
  wire [13:0] _GEN_12224 = 14'h2fc0 == index ? 14'h9f : _GEN_12223;
  wire [13:0] _GEN_12225 = 14'h2fc1 == index ? 14'h9e : _GEN_12224;
  wire [13:0] _GEN_12226 = 14'h2fc2 == index ? 14'h9d : _GEN_12225;
  wire [13:0] _GEN_12227 = 14'h2fc3 == index ? 14'h9c : _GEN_12226;
  wire [13:0] _GEN_12228 = 14'h2fc4 == index ? 14'h9b : _GEN_12227;
  wire [13:0] _GEN_12229 = 14'h2fc5 == index ? 14'h9a : _GEN_12228;
  wire [13:0] _GEN_12230 = 14'h2fc6 == index ? 14'h99 : _GEN_12229;
  wire [13:0] _GEN_12231 = 14'h2fc7 == index ? 14'h98 : _GEN_12230;
  wire [13:0] _GEN_12232 = 14'h2fc8 == index ? 14'h97 : _GEN_12231;
  wire [13:0] _GEN_12233 = 14'h2fc9 == index ? 14'h96 : _GEN_12232;
  wire [13:0] _GEN_12234 = 14'h2fca == index ? 14'h95 : _GEN_12233;
  wire [13:0] _GEN_12235 = 14'h2fcb == index ? 14'h94 : _GEN_12234;
  wire [13:0] _GEN_12236 = 14'h2fcc == index ? 14'h93 : _GEN_12235;
  wire [13:0] _GEN_12237 = 14'h2fcd == index ? 14'h92 : _GEN_12236;
  wire [13:0] _GEN_12238 = 14'h2fce == index ? 14'h91 : _GEN_12237;
  wire [13:0] _GEN_12239 = 14'h2fcf == index ? 14'h90 : _GEN_12238;
  wire [13:0] _GEN_12240 = 14'h2fd0 == index ? 14'h8f : _GEN_12239;
  wire [13:0] _GEN_12241 = 14'h2fd1 == index ? 14'h8e : _GEN_12240;
  wire [13:0] _GEN_12242 = 14'h2fd2 == index ? 14'h8d : _GEN_12241;
  wire [13:0] _GEN_12243 = 14'h2fd3 == index ? 14'h8c : _GEN_12242;
  wire [13:0] _GEN_12244 = 14'h2fd4 == index ? 14'h8b : _GEN_12243;
  wire [13:0] _GEN_12245 = 14'h2fd5 == index ? 14'h8a : _GEN_12244;
  wire [13:0] _GEN_12246 = 14'h2fd6 == index ? 14'h89 : _GEN_12245;
  wire [13:0] _GEN_12247 = 14'h2fd7 == index ? 14'h88 : _GEN_12246;
  wire [13:0] _GEN_12248 = 14'h2fd8 == index ? 14'h87 : _GEN_12247;
  wire [13:0] _GEN_12249 = 14'h2fd9 == index ? 14'h86 : _GEN_12248;
  wire [13:0] _GEN_12250 = 14'h2fda == index ? 14'h85 : _GEN_12249;
  wire [13:0] _GEN_12251 = 14'h2fdb == index ? 14'h84 : _GEN_12250;
  wire [13:0] _GEN_12252 = 14'h2fdc == index ? 14'h83 : _GEN_12251;
  wire [13:0] _GEN_12253 = 14'h2fdd == index ? 14'h82 : _GEN_12252;
  wire [13:0] _GEN_12254 = 14'h2fde == index ? 14'h81 : _GEN_12253;
  wire [13:0] _GEN_12255 = 14'h2fdf == index ? 14'h80 : _GEN_12254;
  wire [13:0] _GEN_12256 = 14'h2fe0 == index ? 14'h5f : _GEN_12255;
  wire [13:0] _GEN_12257 = 14'h2fe1 == index ? 14'h5f : _GEN_12256;
  wire [13:0] _GEN_12258 = 14'h2fe2 == index ? 14'h5f : _GEN_12257;
  wire [13:0] _GEN_12259 = 14'h2fe3 == index ? 14'h5f : _GEN_12258;
  wire [13:0] _GEN_12260 = 14'h2fe4 == index ? 14'h5f : _GEN_12259;
  wire [13:0] _GEN_12261 = 14'h2fe5 == index ? 14'h5f : _GEN_12260;
  wire [13:0] _GEN_12262 = 14'h2fe6 == index ? 14'h5f : _GEN_12261;
  wire [13:0] _GEN_12263 = 14'h2fe7 == index ? 14'h5f : _GEN_12262;
  wire [13:0] _GEN_12264 = 14'h2fe8 == index ? 14'h5f : _GEN_12263;
  wire [13:0] _GEN_12265 = 14'h2fe9 == index ? 14'h5f : _GEN_12264;
  wire [13:0] _GEN_12266 = 14'h2fea == index ? 14'h5f : _GEN_12265;
  wire [13:0] _GEN_12267 = 14'h2feb == index ? 14'h5f : _GEN_12266;
  wire [13:0] _GEN_12268 = 14'h2fec == index ? 14'h5f : _GEN_12267;
  wire [13:0] _GEN_12269 = 14'h2fed == index ? 14'h5f : _GEN_12268;
  wire [13:0] _GEN_12270 = 14'h2fee == index ? 14'h5f : _GEN_12269;
  wire [13:0] _GEN_12271 = 14'h2fef == index ? 14'h5f : _GEN_12270;
  wire [13:0] _GEN_12272 = 14'h2ff0 == index ? 14'h5f : _GEN_12271;
  wire [13:0] _GEN_12273 = 14'h2ff1 == index ? 14'h5f : _GEN_12272;
  wire [13:0] _GEN_12274 = 14'h2ff2 == index ? 14'h5f : _GEN_12273;
  wire [13:0] _GEN_12275 = 14'h2ff3 == index ? 14'h5f : _GEN_12274;
  wire [13:0] _GEN_12276 = 14'h2ff4 == index ? 14'h5f : _GEN_12275;
  wire [13:0] _GEN_12277 = 14'h2ff5 == index ? 14'h5f : _GEN_12276;
  wire [13:0] _GEN_12278 = 14'h2ff6 == index ? 14'h5f : _GEN_12277;
  wire [13:0] _GEN_12279 = 14'h2ff7 == index ? 14'h5f : _GEN_12278;
  wire [13:0] _GEN_12280 = 14'h2ff8 == index ? 14'h5f : _GEN_12279;
  wire [13:0] _GEN_12281 = 14'h2ff9 == index ? 14'h5f : _GEN_12280;
  wire [13:0] _GEN_12282 = 14'h2ffa == index ? 14'h5f : _GEN_12281;
  wire [13:0] _GEN_12283 = 14'h2ffb == index ? 14'h5f : _GEN_12282;
  wire [13:0] _GEN_12284 = 14'h2ffc == index ? 14'h5f : _GEN_12283;
  wire [13:0] _GEN_12285 = 14'h2ffd == index ? 14'h5f : _GEN_12284;
  wire [13:0] _GEN_12286 = 14'h2ffe == index ? 14'h5f : _GEN_12285;
  wire [13:0] _GEN_12287 = 14'h2fff == index ? 14'h5f : _GEN_12286;
  wire [13:0] _GEN_12288 = 14'h3000 == index ? 14'h0 : _GEN_12287;
  wire [13:0] _GEN_12289 = 14'h3001 == index ? 14'h3000 : _GEN_12288;
  wire [13:0] _GEN_12290 = 14'h3002 == index ? 14'h1800 : _GEN_12289;
  wire [13:0] _GEN_12291 = 14'h3003 == index ? 14'h1000 : _GEN_12290;
  wire [13:0] _GEN_12292 = 14'h3004 == index ? 14'hc00 : _GEN_12291;
  wire [13:0] _GEN_12293 = 14'h3005 == index ? 14'h981 : _GEN_12292;
  wire [13:0] _GEN_12294 = 14'h3006 == index ? 14'h800 : _GEN_12293;
  wire [13:0] _GEN_12295 = 14'h3007 == index ? 14'h685 : _GEN_12294;
  wire [13:0] _GEN_12296 = 14'h3008 == index ? 14'h600 : _GEN_12295;
  wire [13:0] _GEN_12297 = 14'h3009 == index ? 14'h506 : _GEN_12296;
  wire [13:0] _GEN_12298 = 14'h300a == index ? 14'h486 : _GEN_12297;
  wire [13:0] _GEN_12299 = 14'h300b == index ? 14'h408 : _GEN_12298;
  wire [13:0] _GEN_12300 = 14'h300c == index ? 14'h400 : _GEN_12299;
  wire [13:0] _GEN_12301 = 14'h300d == index ? 14'h385 : _GEN_12300;
  wire [13:0] _GEN_12302 = 14'h300e == index ? 14'h30c : _GEN_12301;
  wire [13:0] _GEN_12303 = 14'h300f == index ? 14'h306 : _GEN_12302;
  wire [13:0] _GEN_12304 = 14'h3010 == index ? 14'h300 : _GEN_12303;
  wire [13:0] _GEN_12305 = 14'h3011 == index ? 14'h28b : _GEN_12304;
  wire [13:0] _GEN_12306 = 14'h3012 == index ? 14'h286 : _GEN_12305;
  wire [13:0] _GEN_12307 = 14'h3013 == index ? 14'h281 : _GEN_12306;
  wire [13:0] _GEN_12308 = 14'h3014 == index ? 14'h210 : _GEN_12307;
  wire [13:0] _GEN_12309 = 14'h3015 == index ? 14'h20c : _GEN_12308;
  wire [13:0] _GEN_12310 = 14'h3016 == index ? 14'h208 : _GEN_12309;
  wire [13:0] _GEN_12311 = 14'h3017 == index ? 14'h204 : _GEN_12310;
  wire [13:0] _GEN_12312 = 14'h3018 == index ? 14'h200 : _GEN_12311;
  wire [13:0] _GEN_12313 = 14'h3019 == index ? 14'h195 : _GEN_12312;
  wire [13:0] _GEN_12314 = 14'h301a == index ? 14'h192 : _GEN_12313;
  wire [13:0] _GEN_12315 = 14'h301b == index ? 14'h18f : _GEN_12314;
  wire [13:0] _GEN_12316 = 14'h301c == index ? 14'h18c : _GEN_12315;
  wire [13:0] _GEN_12317 = 14'h301d == index ? 14'h189 : _GEN_12316;
  wire [13:0] _GEN_12318 = 14'h301e == index ? 14'h186 : _GEN_12317;
  wire [13:0] _GEN_12319 = 14'h301f == index ? 14'h183 : _GEN_12318;
  wire [13:0] _GEN_12320 = 14'h3020 == index ? 14'h180 : _GEN_12319;
  wire [13:0] _GEN_12321 = 14'h3021 == index ? 14'h11e : _GEN_12320;
  wire [13:0] _GEN_12322 = 14'h3022 == index ? 14'h11c : _GEN_12321;
  wire [13:0] _GEN_12323 = 14'h3023 == index ? 14'h11a : _GEN_12322;
  wire [13:0] _GEN_12324 = 14'h3024 == index ? 14'h118 : _GEN_12323;
  wire [13:0] _GEN_12325 = 14'h3025 == index ? 14'h116 : _GEN_12324;
  wire [13:0] _GEN_12326 = 14'h3026 == index ? 14'h114 : _GEN_12325;
  wire [13:0] _GEN_12327 = 14'h3027 == index ? 14'h112 : _GEN_12326;
  wire [13:0] _GEN_12328 = 14'h3028 == index ? 14'h110 : _GEN_12327;
  wire [13:0] _GEN_12329 = 14'h3029 == index ? 14'h10e : _GEN_12328;
  wire [13:0] _GEN_12330 = 14'h302a == index ? 14'h10c : _GEN_12329;
  wire [13:0] _GEN_12331 = 14'h302b == index ? 14'h10a : _GEN_12330;
  wire [13:0] _GEN_12332 = 14'h302c == index ? 14'h108 : _GEN_12331;
  wire [13:0] _GEN_12333 = 14'h302d == index ? 14'h106 : _GEN_12332;
  wire [13:0] _GEN_12334 = 14'h302e == index ? 14'h104 : _GEN_12333;
  wire [13:0] _GEN_12335 = 14'h302f == index ? 14'h102 : _GEN_12334;
  wire [13:0] _GEN_12336 = 14'h3030 == index ? 14'h100 : _GEN_12335;
  wire [13:0] _GEN_12337 = 14'h3031 == index ? 14'haf : _GEN_12336;
  wire [13:0] _GEN_12338 = 14'h3032 == index ? 14'hae : _GEN_12337;
  wire [13:0] _GEN_12339 = 14'h3033 == index ? 14'had : _GEN_12338;
  wire [13:0] _GEN_12340 = 14'h3034 == index ? 14'hac : _GEN_12339;
  wire [13:0] _GEN_12341 = 14'h3035 == index ? 14'hab : _GEN_12340;
  wire [13:0] _GEN_12342 = 14'h3036 == index ? 14'haa : _GEN_12341;
  wire [13:0] _GEN_12343 = 14'h3037 == index ? 14'ha9 : _GEN_12342;
  wire [13:0] _GEN_12344 = 14'h3038 == index ? 14'ha8 : _GEN_12343;
  wire [13:0] _GEN_12345 = 14'h3039 == index ? 14'ha7 : _GEN_12344;
  wire [13:0] _GEN_12346 = 14'h303a == index ? 14'ha6 : _GEN_12345;
  wire [13:0] _GEN_12347 = 14'h303b == index ? 14'ha5 : _GEN_12346;
  wire [13:0] _GEN_12348 = 14'h303c == index ? 14'ha4 : _GEN_12347;
  wire [13:0] _GEN_12349 = 14'h303d == index ? 14'ha3 : _GEN_12348;
  wire [13:0] _GEN_12350 = 14'h303e == index ? 14'ha2 : _GEN_12349;
  wire [13:0] _GEN_12351 = 14'h303f == index ? 14'ha1 : _GEN_12350;
  wire [13:0] _GEN_12352 = 14'h3040 == index ? 14'ha0 : _GEN_12351;
  wire [13:0] _GEN_12353 = 14'h3041 == index ? 14'h9f : _GEN_12352;
  wire [13:0] _GEN_12354 = 14'h3042 == index ? 14'h9e : _GEN_12353;
  wire [13:0] _GEN_12355 = 14'h3043 == index ? 14'h9d : _GEN_12354;
  wire [13:0] _GEN_12356 = 14'h3044 == index ? 14'h9c : _GEN_12355;
  wire [13:0] _GEN_12357 = 14'h3045 == index ? 14'h9b : _GEN_12356;
  wire [13:0] _GEN_12358 = 14'h3046 == index ? 14'h9a : _GEN_12357;
  wire [13:0] _GEN_12359 = 14'h3047 == index ? 14'h99 : _GEN_12358;
  wire [13:0] _GEN_12360 = 14'h3048 == index ? 14'h98 : _GEN_12359;
  wire [13:0] _GEN_12361 = 14'h3049 == index ? 14'h97 : _GEN_12360;
  wire [13:0] _GEN_12362 = 14'h304a == index ? 14'h96 : _GEN_12361;
  wire [13:0] _GEN_12363 = 14'h304b == index ? 14'h95 : _GEN_12362;
  wire [13:0] _GEN_12364 = 14'h304c == index ? 14'h94 : _GEN_12363;
  wire [13:0] _GEN_12365 = 14'h304d == index ? 14'h93 : _GEN_12364;
  wire [13:0] _GEN_12366 = 14'h304e == index ? 14'h92 : _GEN_12365;
  wire [13:0] _GEN_12367 = 14'h304f == index ? 14'h91 : _GEN_12366;
  wire [13:0] _GEN_12368 = 14'h3050 == index ? 14'h90 : _GEN_12367;
  wire [13:0] _GEN_12369 = 14'h3051 == index ? 14'h8f : _GEN_12368;
  wire [13:0] _GEN_12370 = 14'h3052 == index ? 14'h8e : _GEN_12369;
  wire [13:0] _GEN_12371 = 14'h3053 == index ? 14'h8d : _GEN_12370;
  wire [13:0] _GEN_12372 = 14'h3054 == index ? 14'h8c : _GEN_12371;
  wire [13:0] _GEN_12373 = 14'h3055 == index ? 14'h8b : _GEN_12372;
  wire [13:0] _GEN_12374 = 14'h3056 == index ? 14'h8a : _GEN_12373;
  wire [13:0] _GEN_12375 = 14'h3057 == index ? 14'h89 : _GEN_12374;
  wire [13:0] _GEN_12376 = 14'h3058 == index ? 14'h88 : _GEN_12375;
  wire [13:0] _GEN_12377 = 14'h3059 == index ? 14'h87 : _GEN_12376;
  wire [13:0] _GEN_12378 = 14'h305a == index ? 14'h86 : _GEN_12377;
  wire [13:0] _GEN_12379 = 14'h305b == index ? 14'h85 : _GEN_12378;
  wire [13:0] _GEN_12380 = 14'h305c == index ? 14'h84 : _GEN_12379;
  wire [13:0] _GEN_12381 = 14'h305d == index ? 14'h83 : _GEN_12380;
  wire [13:0] _GEN_12382 = 14'h305e == index ? 14'h82 : _GEN_12381;
  wire [13:0] _GEN_12383 = 14'h305f == index ? 14'h81 : _GEN_12382;
  wire [13:0] _GEN_12384 = 14'h3060 == index ? 14'h80 : _GEN_12383;
  wire [13:0] _GEN_12385 = 14'h3061 == index ? 14'h60 : _GEN_12384;
  wire [13:0] _GEN_12386 = 14'h3062 == index ? 14'h60 : _GEN_12385;
  wire [13:0] _GEN_12387 = 14'h3063 == index ? 14'h60 : _GEN_12386;
  wire [13:0] _GEN_12388 = 14'h3064 == index ? 14'h60 : _GEN_12387;
  wire [13:0] _GEN_12389 = 14'h3065 == index ? 14'h60 : _GEN_12388;
  wire [13:0] _GEN_12390 = 14'h3066 == index ? 14'h60 : _GEN_12389;
  wire [13:0] _GEN_12391 = 14'h3067 == index ? 14'h60 : _GEN_12390;
  wire [13:0] _GEN_12392 = 14'h3068 == index ? 14'h60 : _GEN_12391;
  wire [13:0] _GEN_12393 = 14'h3069 == index ? 14'h60 : _GEN_12392;
  wire [13:0] _GEN_12394 = 14'h306a == index ? 14'h60 : _GEN_12393;
  wire [13:0] _GEN_12395 = 14'h306b == index ? 14'h60 : _GEN_12394;
  wire [13:0] _GEN_12396 = 14'h306c == index ? 14'h60 : _GEN_12395;
  wire [13:0] _GEN_12397 = 14'h306d == index ? 14'h60 : _GEN_12396;
  wire [13:0] _GEN_12398 = 14'h306e == index ? 14'h60 : _GEN_12397;
  wire [13:0] _GEN_12399 = 14'h306f == index ? 14'h60 : _GEN_12398;
  wire [13:0] _GEN_12400 = 14'h3070 == index ? 14'h60 : _GEN_12399;
  wire [13:0] _GEN_12401 = 14'h3071 == index ? 14'h60 : _GEN_12400;
  wire [13:0] _GEN_12402 = 14'h3072 == index ? 14'h60 : _GEN_12401;
  wire [13:0] _GEN_12403 = 14'h3073 == index ? 14'h60 : _GEN_12402;
  wire [13:0] _GEN_12404 = 14'h3074 == index ? 14'h60 : _GEN_12403;
  wire [13:0] _GEN_12405 = 14'h3075 == index ? 14'h60 : _GEN_12404;
  wire [13:0] _GEN_12406 = 14'h3076 == index ? 14'h60 : _GEN_12405;
  wire [13:0] _GEN_12407 = 14'h3077 == index ? 14'h60 : _GEN_12406;
  wire [13:0] _GEN_12408 = 14'h3078 == index ? 14'h60 : _GEN_12407;
  wire [13:0] _GEN_12409 = 14'h3079 == index ? 14'h60 : _GEN_12408;
  wire [13:0] _GEN_12410 = 14'h307a == index ? 14'h60 : _GEN_12409;
  wire [13:0] _GEN_12411 = 14'h307b == index ? 14'h60 : _GEN_12410;
  wire [13:0] _GEN_12412 = 14'h307c == index ? 14'h60 : _GEN_12411;
  wire [13:0] _GEN_12413 = 14'h307d == index ? 14'h60 : _GEN_12412;
  wire [13:0] _GEN_12414 = 14'h307e == index ? 14'h60 : _GEN_12413;
  wire [13:0] _GEN_12415 = 14'h307f == index ? 14'h60 : _GEN_12414;
  wire [13:0] _GEN_12416 = 14'h3080 == index ? 14'h0 : _GEN_12415;
  wire [13:0] _GEN_12417 = 14'h3081 == index ? 14'h3080 : _GEN_12416;
  wire [13:0] _GEN_12418 = 14'h3082 == index ? 14'h1801 : _GEN_12417;
  wire [13:0] _GEN_12419 = 14'h3083 == index ? 14'h1001 : _GEN_12418;
  wire [13:0] _GEN_12420 = 14'h3084 == index ? 14'hc01 : _GEN_12419;
  wire [13:0] _GEN_12421 = 14'h3085 == index ? 14'h982 : _GEN_12420;
  wire [13:0] _GEN_12422 = 14'h3086 == index ? 14'h801 : _GEN_12421;
  wire [13:0] _GEN_12423 = 14'h3087 == index ? 14'h686 : _GEN_12422;
  wire [13:0] _GEN_12424 = 14'h3088 == index ? 14'h601 : _GEN_12423;
  wire [13:0] _GEN_12425 = 14'h3089 == index ? 14'h507 : _GEN_12424;
  wire [13:0] _GEN_12426 = 14'h308a == index ? 14'h487 : _GEN_12425;
  wire [13:0] _GEN_12427 = 14'h308b == index ? 14'h409 : _GEN_12426;
  wire [13:0] _GEN_12428 = 14'h308c == index ? 14'h401 : _GEN_12427;
  wire [13:0] _GEN_12429 = 14'h308d == index ? 14'h386 : _GEN_12428;
  wire [13:0] _GEN_12430 = 14'h308e == index ? 14'h30d : _GEN_12429;
  wire [13:0] _GEN_12431 = 14'h308f == index ? 14'h307 : _GEN_12430;
  wire [13:0] _GEN_12432 = 14'h3090 == index ? 14'h301 : _GEN_12431;
  wire [13:0] _GEN_12433 = 14'h3091 == index ? 14'h28c : _GEN_12432;
  wire [13:0] _GEN_12434 = 14'h3092 == index ? 14'h287 : _GEN_12433;
  wire [13:0] _GEN_12435 = 14'h3093 == index ? 14'h282 : _GEN_12434;
  wire [13:0] _GEN_12436 = 14'h3094 == index ? 14'h211 : _GEN_12435;
  wire [13:0] _GEN_12437 = 14'h3095 == index ? 14'h20d : _GEN_12436;
  wire [13:0] _GEN_12438 = 14'h3096 == index ? 14'h209 : _GEN_12437;
  wire [13:0] _GEN_12439 = 14'h3097 == index ? 14'h205 : _GEN_12438;
  wire [13:0] _GEN_12440 = 14'h3098 == index ? 14'h201 : _GEN_12439;
  wire [13:0] _GEN_12441 = 14'h3099 == index ? 14'h196 : _GEN_12440;
  wire [13:0] _GEN_12442 = 14'h309a == index ? 14'h193 : _GEN_12441;
  wire [13:0] _GEN_12443 = 14'h309b == index ? 14'h190 : _GEN_12442;
  wire [13:0] _GEN_12444 = 14'h309c == index ? 14'h18d : _GEN_12443;
  wire [13:0] _GEN_12445 = 14'h309d == index ? 14'h18a : _GEN_12444;
  wire [13:0] _GEN_12446 = 14'h309e == index ? 14'h187 : _GEN_12445;
  wire [13:0] _GEN_12447 = 14'h309f == index ? 14'h184 : _GEN_12446;
  wire [13:0] _GEN_12448 = 14'h30a0 == index ? 14'h181 : _GEN_12447;
  wire [13:0] _GEN_12449 = 14'h30a1 == index ? 14'h11f : _GEN_12448;
  wire [13:0] _GEN_12450 = 14'h30a2 == index ? 14'h11d : _GEN_12449;
  wire [13:0] _GEN_12451 = 14'h30a3 == index ? 14'h11b : _GEN_12450;
  wire [13:0] _GEN_12452 = 14'h30a4 == index ? 14'h119 : _GEN_12451;
  wire [13:0] _GEN_12453 = 14'h30a5 == index ? 14'h117 : _GEN_12452;
  wire [13:0] _GEN_12454 = 14'h30a6 == index ? 14'h115 : _GEN_12453;
  wire [13:0] _GEN_12455 = 14'h30a7 == index ? 14'h113 : _GEN_12454;
  wire [13:0] _GEN_12456 = 14'h30a8 == index ? 14'h111 : _GEN_12455;
  wire [13:0] _GEN_12457 = 14'h30a9 == index ? 14'h10f : _GEN_12456;
  wire [13:0] _GEN_12458 = 14'h30aa == index ? 14'h10d : _GEN_12457;
  wire [13:0] _GEN_12459 = 14'h30ab == index ? 14'h10b : _GEN_12458;
  wire [13:0] _GEN_12460 = 14'h30ac == index ? 14'h109 : _GEN_12459;
  wire [13:0] _GEN_12461 = 14'h30ad == index ? 14'h107 : _GEN_12460;
  wire [13:0] _GEN_12462 = 14'h30ae == index ? 14'h105 : _GEN_12461;
  wire [13:0] _GEN_12463 = 14'h30af == index ? 14'h103 : _GEN_12462;
  wire [13:0] _GEN_12464 = 14'h30b0 == index ? 14'h101 : _GEN_12463;
  wire [13:0] _GEN_12465 = 14'h30b1 == index ? 14'hb0 : _GEN_12464;
  wire [13:0] _GEN_12466 = 14'h30b2 == index ? 14'haf : _GEN_12465;
  wire [13:0] _GEN_12467 = 14'h30b3 == index ? 14'hae : _GEN_12466;
  wire [13:0] _GEN_12468 = 14'h30b4 == index ? 14'had : _GEN_12467;
  wire [13:0] _GEN_12469 = 14'h30b5 == index ? 14'hac : _GEN_12468;
  wire [13:0] _GEN_12470 = 14'h30b6 == index ? 14'hab : _GEN_12469;
  wire [13:0] _GEN_12471 = 14'h30b7 == index ? 14'haa : _GEN_12470;
  wire [13:0] _GEN_12472 = 14'h30b8 == index ? 14'ha9 : _GEN_12471;
  wire [13:0] _GEN_12473 = 14'h30b9 == index ? 14'ha8 : _GEN_12472;
  wire [13:0] _GEN_12474 = 14'h30ba == index ? 14'ha7 : _GEN_12473;
  wire [13:0] _GEN_12475 = 14'h30bb == index ? 14'ha6 : _GEN_12474;
  wire [13:0] _GEN_12476 = 14'h30bc == index ? 14'ha5 : _GEN_12475;
  wire [13:0] _GEN_12477 = 14'h30bd == index ? 14'ha4 : _GEN_12476;
  wire [13:0] _GEN_12478 = 14'h30be == index ? 14'ha3 : _GEN_12477;
  wire [13:0] _GEN_12479 = 14'h30bf == index ? 14'ha2 : _GEN_12478;
  wire [13:0] _GEN_12480 = 14'h30c0 == index ? 14'ha1 : _GEN_12479;
  wire [13:0] _GEN_12481 = 14'h30c1 == index ? 14'ha0 : _GEN_12480;
  wire [13:0] _GEN_12482 = 14'h30c2 == index ? 14'h9f : _GEN_12481;
  wire [13:0] _GEN_12483 = 14'h30c3 == index ? 14'h9e : _GEN_12482;
  wire [13:0] _GEN_12484 = 14'h30c4 == index ? 14'h9d : _GEN_12483;
  wire [13:0] _GEN_12485 = 14'h30c5 == index ? 14'h9c : _GEN_12484;
  wire [13:0] _GEN_12486 = 14'h30c6 == index ? 14'h9b : _GEN_12485;
  wire [13:0] _GEN_12487 = 14'h30c7 == index ? 14'h9a : _GEN_12486;
  wire [13:0] _GEN_12488 = 14'h30c8 == index ? 14'h99 : _GEN_12487;
  wire [13:0] _GEN_12489 = 14'h30c9 == index ? 14'h98 : _GEN_12488;
  wire [13:0] _GEN_12490 = 14'h30ca == index ? 14'h97 : _GEN_12489;
  wire [13:0] _GEN_12491 = 14'h30cb == index ? 14'h96 : _GEN_12490;
  wire [13:0] _GEN_12492 = 14'h30cc == index ? 14'h95 : _GEN_12491;
  wire [13:0] _GEN_12493 = 14'h30cd == index ? 14'h94 : _GEN_12492;
  wire [13:0] _GEN_12494 = 14'h30ce == index ? 14'h93 : _GEN_12493;
  wire [13:0] _GEN_12495 = 14'h30cf == index ? 14'h92 : _GEN_12494;
  wire [13:0] _GEN_12496 = 14'h30d0 == index ? 14'h91 : _GEN_12495;
  wire [13:0] _GEN_12497 = 14'h30d1 == index ? 14'h90 : _GEN_12496;
  wire [13:0] _GEN_12498 = 14'h30d2 == index ? 14'h8f : _GEN_12497;
  wire [13:0] _GEN_12499 = 14'h30d3 == index ? 14'h8e : _GEN_12498;
  wire [13:0] _GEN_12500 = 14'h30d4 == index ? 14'h8d : _GEN_12499;
  wire [13:0] _GEN_12501 = 14'h30d5 == index ? 14'h8c : _GEN_12500;
  wire [13:0] _GEN_12502 = 14'h30d6 == index ? 14'h8b : _GEN_12501;
  wire [13:0] _GEN_12503 = 14'h30d7 == index ? 14'h8a : _GEN_12502;
  wire [13:0] _GEN_12504 = 14'h30d8 == index ? 14'h89 : _GEN_12503;
  wire [13:0] _GEN_12505 = 14'h30d9 == index ? 14'h88 : _GEN_12504;
  wire [13:0] _GEN_12506 = 14'h30da == index ? 14'h87 : _GEN_12505;
  wire [13:0] _GEN_12507 = 14'h30db == index ? 14'h86 : _GEN_12506;
  wire [13:0] _GEN_12508 = 14'h30dc == index ? 14'h85 : _GEN_12507;
  wire [13:0] _GEN_12509 = 14'h30dd == index ? 14'h84 : _GEN_12508;
  wire [13:0] _GEN_12510 = 14'h30de == index ? 14'h83 : _GEN_12509;
  wire [13:0] _GEN_12511 = 14'h30df == index ? 14'h82 : _GEN_12510;
  wire [13:0] _GEN_12512 = 14'h30e0 == index ? 14'h81 : _GEN_12511;
  wire [13:0] _GEN_12513 = 14'h30e1 == index ? 14'h80 : _GEN_12512;
  wire [13:0] _GEN_12514 = 14'h30e2 == index ? 14'h61 : _GEN_12513;
  wire [13:0] _GEN_12515 = 14'h30e3 == index ? 14'h61 : _GEN_12514;
  wire [13:0] _GEN_12516 = 14'h30e4 == index ? 14'h61 : _GEN_12515;
  wire [13:0] _GEN_12517 = 14'h30e5 == index ? 14'h61 : _GEN_12516;
  wire [13:0] _GEN_12518 = 14'h30e6 == index ? 14'h61 : _GEN_12517;
  wire [13:0] _GEN_12519 = 14'h30e7 == index ? 14'h61 : _GEN_12518;
  wire [13:0] _GEN_12520 = 14'h30e8 == index ? 14'h61 : _GEN_12519;
  wire [13:0] _GEN_12521 = 14'h30e9 == index ? 14'h61 : _GEN_12520;
  wire [13:0] _GEN_12522 = 14'h30ea == index ? 14'h61 : _GEN_12521;
  wire [13:0] _GEN_12523 = 14'h30eb == index ? 14'h61 : _GEN_12522;
  wire [13:0] _GEN_12524 = 14'h30ec == index ? 14'h61 : _GEN_12523;
  wire [13:0] _GEN_12525 = 14'h30ed == index ? 14'h61 : _GEN_12524;
  wire [13:0] _GEN_12526 = 14'h30ee == index ? 14'h61 : _GEN_12525;
  wire [13:0] _GEN_12527 = 14'h30ef == index ? 14'h61 : _GEN_12526;
  wire [13:0] _GEN_12528 = 14'h30f0 == index ? 14'h61 : _GEN_12527;
  wire [13:0] _GEN_12529 = 14'h30f1 == index ? 14'h61 : _GEN_12528;
  wire [13:0] _GEN_12530 = 14'h30f2 == index ? 14'h61 : _GEN_12529;
  wire [13:0] _GEN_12531 = 14'h30f3 == index ? 14'h61 : _GEN_12530;
  wire [13:0] _GEN_12532 = 14'h30f4 == index ? 14'h61 : _GEN_12531;
  wire [13:0] _GEN_12533 = 14'h30f5 == index ? 14'h61 : _GEN_12532;
  wire [13:0] _GEN_12534 = 14'h30f6 == index ? 14'h61 : _GEN_12533;
  wire [13:0] _GEN_12535 = 14'h30f7 == index ? 14'h61 : _GEN_12534;
  wire [13:0] _GEN_12536 = 14'h30f8 == index ? 14'h61 : _GEN_12535;
  wire [13:0] _GEN_12537 = 14'h30f9 == index ? 14'h61 : _GEN_12536;
  wire [13:0] _GEN_12538 = 14'h30fa == index ? 14'h61 : _GEN_12537;
  wire [13:0] _GEN_12539 = 14'h30fb == index ? 14'h61 : _GEN_12538;
  wire [13:0] _GEN_12540 = 14'h30fc == index ? 14'h61 : _GEN_12539;
  wire [13:0] _GEN_12541 = 14'h30fd == index ? 14'h61 : _GEN_12540;
  wire [13:0] _GEN_12542 = 14'h30fe == index ? 14'h61 : _GEN_12541;
  wire [13:0] _GEN_12543 = 14'h30ff == index ? 14'h61 : _GEN_12542;
  wire [13:0] _GEN_12544 = 14'h3100 == index ? 14'h0 : _GEN_12543;
  wire [13:0] _GEN_12545 = 14'h3101 == index ? 14'h3100 : _GEN_12544;
  wire [13:0] _GEN_12546 = 14'h3102 == index ? 14'h1880 : _GEN_12545;
  wire [13:0] _GEN_12547 = 14'h3103 == index ? 14'h1002 : _GEN_12546;
  wire [13:0] _GEN_12548 = 14'h3104 == index ? 14'hc02 : _GEN_12547;
  wire [13:0] _GEN_12549 = 14'h3105 == index ? 14'h983 : _GEN_12548;
  wire [13:0] _GEN_12550 = 14'h3106 == index ? 14'h802 : _GEN_12549;
  wire [13:0] _GEN_12551 = 14'h3107 == index ? 14'h700 : _GEN_12550;
  wire [13:0] _GEN_12552 = 14'h3108 == index ? 14'h602 : _GEN_12551;
  wire [13:0] _GEN_12553 = 14'h3109 == index ? 14'h508 : _GEN_12552;
  wire [13:0] _GEN_12554 = 14'h310a == index ? 14'h488 : _GEN_12553;
  wire [13:0] _GEN_12555 = 14'h310b == index ? 14'h40a : _GEN_12554;
  wire [13:0] _GEN_12556 = 14'h310c == index ? 14'h402 : _GEN_12555;
  wire [13:0] _GEN_12557 = 14'h310d == index ? 14'h387 : _GEN_12556;
  wire [13:0] _GEN_12558 = 14'h310e == index ? 14'h380 : _GEN_12557;
  wire [13:0] _GEN_12559 = 14'h310f == index ? 14'h308 : _GEN_12558;
  wire [13:0] _GEN_12560 = 14'h3110 == index ? 14'h302 : _GEN_12559;
  wire [13:0] _GEN_12561 = 14'h3111 == index ? 14'h28d : _GEN_12560;
  wire [13:0] _GEN_12562 = 14'h3112 == index ? 14'h288 : _GEN_12561;
  wire [13:0] _GEN_12563 = 14'h3113 == index ? 14'h283 : _GEN_12562;
  wire [13:0] _GEN_12564 = 14'h3114 == index ? 14'h212 : _GEN_12563;
  wire [13:0] _GEN_12565 = 14'h3115 == index ? 14'h20e : _GEN_12564;
  wire [13:0] _GEN_12566 = 14'h3116 == index ? 14'h20a : _GEN_12565;
  wire [13:0] _GEN_12567 = 14'h3117 == index ? 14'h206 : _GEN_12566;
  wire [13:0] _GEN_12568 = 14'h3118 == index ? 14'h202 : _GEN_12567;
  wire [13:0] _GEN_12569 = 14'h3119 == index ? 14'h197 : _GEN_12568;
  wire [13:0] _GEN_12570 = 14'h311a == index ? 14'h194 : _GEN_12569;
  wire [13:0] _GEN_12571 = 14'h311b == index ? 14'h191 : _GEN_12570;
  wire [13:0] _GEN_12572 = 14'h311c == index ? 14'h18e : _GEN_12571;
  wire [13:0] _GEN_12573 = 14'h311d == index ? 14'h18b : _GEN_12572;
  wire [13:0] _GEN_12574 = 14'h311e == index ? 14'h188 : _GEN_12573;
  wire [13:0] _GEN_12575 = 14'h311f == index ? 14'h185 : _GEN_12574;
  wire [13:0] _GEN_12576 = 14'h3120 == index ? 14'h182 : _GEN_12575;
  wire [13:0] _GEN_12577 = 14'h3121 == index ? 14'h120 : _GEN_12576;
  wire [13:0] _GEN_12578 = 14'h3122 == index ? 14'h11e : _GEN_12577;
  wire [13:0] _GEN_12579 = 14'h3123 == index ? 14'h11c : _GEN_12578;
  wire [13:0] _GEN_12580 = 14'h3124 == index ? 14'h11a : _GEN_12579;
  wire [13:0] _GEN_12581 = 14'h3125 == index ? 14'h118 : _GEN_12580;
  wire [13:0] _GEN_12582 = 14'h3126 == index ? 14'h116 : _GEN_12581;
  wire [13:0] _GEN_12583 = 14'h3127 == index ? 14'h114 : _GEN_12582;
  wire [13:0] _GEN_12584 = 14'h3128 == index ? 14'h112 : _GEN_12583;
  wire [13:0] _GEN_12585 = 14'h3129 == index ? 14'h110 : _GEN_12584;
  wire [13:0] _GEN_12586 = 14'h312a == index ? 14'h10e : _GEN_12585;
  wire [13:0] _GEN_12587 = 14'h312b == index ? 14'h10c : _GEN_12586;
  wire [13:0] _GEN_12588 = 14'h312c == index ? 14'h10a : _GEN_12587;
  wire [13:0] _GEN_12589 = 14'h312d == index ? 14'h108 : _GEN_12588;
  wire [13:0] _GEN_12590 = 14'h312e == index ? 14'h106 : _GEN_12589;
  wire [13:0] _GEN_12591 = 14'h312f == index ? 14'h104 : _GEN_12590;
  wire [13:0] _GEN_12592 = 14'h3130 == index ? 14'h102 : _GEN_12591;
  wire [13:0] _GEN_12593 = 14'h3131 == index ? 14'h100 : _GEN_12592;
  wire [13:0] _GEN_12594 = 14'h3132 == index ? 14'hb0 : _GEN_12593;
  wire [13:0] _GEN_12595 = 14'h3133 == index ? 14'haf : _GEN_12594;
  wire [13:0] _GEN_12596 = 14'h3134 == index ? 14'hae : _GEN_12595;
  wire [13:0] _GEN_12597 = 14'h3135 == index ? 14'had : _GEN_12596;
  wire [13:0] _GEN_12598 = 14'h3136 == index ? 14'hac : _GEN_12597;
  wire [13:0] _GEN_12599 = 14'h3137 == index ? 14'hab : _GEN_12598;
  wire [13:0] _GEN_12600 = 14'h3138 == index ? 14'haa : _GEN_12599;
  wire [13:0] _GEN_12601 = 14'h3139 == index ? 14'ha9 : _GEN_12600;
  wire [13:0] _GEN_12602 = 14'h313a == index ? 14'ha8 : _GEN_12601;
  wire [13:0] _GEN_12603 = 14'h313b == index ? 14'ha7 : _GEN_12602;
  wire [13:0] _GEN_12604 = 14'h313c == index ? 14'ha6 : _GEN_12603;
  wire [13:0] _GEN_12605 = 14'h313d == index ? 14'ha5 : _GEN_12604;
  wire [13:0] _GEN_12606 = 14'h313e == index ? 14'ha4 : _GEN_12605;
  wire [13:0] _GEN_12607 = 14'h313f == index ? 14'ha3 : _GEN_12606;
  wire [13:0] _GEN_12608 = 14'h3140 == index ? 14'ha2 : _GEN_12607;
  wire [13:0] _GEN_12609 = 14'h3141 == index ? 14'ha1 : _GEN_12608;
  wire [13:0] _GEN_12610 = 14'h3142 == index ? 14'ha0 : _GEN_12609;
  wire [13:0] _GEN_12611 = 14'h3143 == index ? 14'h9f : _GEN_12610;
  wire [13:0] _GEN_12612 = 14'h3144 == index ? 14'h9e : _GEN_12611;
  wire [13:0] _GEN_12613 = 14'h3145 == index ? 14'h9d : _GEN_12612;
  wire [13:0] _GEN_12614 = 14'h3146 == index ? 14'h9c : _GEN_12613;
  wire [13:0] _GEN_12615 = 14'h3147 == index ? 14'h9b : _GEN_12614;
  wire [13:0] _GEN_12616 = 14'h3148 == index ? 14'h9a : _GEN_12615;
  wire [13:0] _GEN_12617 = 14'h3149 == index ? 14'h99 : _GEN_12616;
  wire [13:0] _GEN_12618 = 14'h314a == index ? 14'h98 : _GEN_12617;
  wire [13:0] _GEN_12619 = 14'h314b == index ? 14'h97 : _GEN_12618;
  wire [13:0] _GEN_12620 = 14'h314c == index ? 14'h96 : _GEN_12619;
  wire [13:0] _GEN_12621 = 14'h314d == index ? 14'h95 : _GEN_12620;
  wire [13:0] _GEN_12622 = 14'h314e == index ? 14'h94 : _GEN_12621;
  wire [13:0] _GEN_12623 = 14'h314f == index ? 14'h93 : _GEN_12622;
  wire [13:0] _GEN_12624 = 14'h3150 == index ? 14'h92 : _GEN_12623;
  wire [13:0] _GEN_12625 = 14'h3151 == index ? 14'h91 : _GEN_12624;
  wire [13:0] _GEN_12626 = 14'h3152 == index ? 14'h90 : _GEN_12625;
  wire [13:0] _GEN_12627 = 14'h3153 == index ? 14'h8f : _GEN_12626;
  wire [13:0] _GEN_12628 = 14'h3154 == index ? 14'h8e : _GEN_12627;
  wire [13:0] _GEN_12629 = 14'h3155 == index ? 14'h8d : _GEN_12628;
  wire [13:0] _GEN_12630 = 14'h3156 == index ? 14'h8c : _GEN_12629;
  wire [13:0] _GEN_12631 = 14'h3157 == index ? 14'h8b : _GEN_12630;
  wire [13:0] _GEN_12632 = 14'h3158 == index ? 14'h8a : _GEN_12631;
  wire [13:0] _GEN_12633 = 14'h3159 == index ? 14'h89 : _GEN_12632;
  wire [13:0] _GEN_12634 = 14'h315a == index ? 14'h88 : _GEN_12633;
  wire [13:0] _GEN_12635 = 14'h315b == index ? 14'h87 : _GEN_12634;
  wire [13:0] _GEN_12636 = 14'h315c == index ? 14'h86 : _GEN_12635;
  wire [13:0] _GEN_12637 = 14'h315d == index ? 14'h85 : _GEN_12636;
  wire [13:0] _GEN_12638 = 14'h315e == index ? 14'h84 : _GEN_12637;
  wire [13:0] _GEN_12639 = 14'h315f == index ? 14'h83 : _GEN_12638;
  wire [13:0] _GEN_12640 = 14'h3160 == index ? 14'h82 : _GEN_12639;
  wire [13:0] _GEN_12641 = 14'h3161 == index ? 14'h81 : _GEN_12640;
  wire [13:0] _GEN_12642 = 14'h3162 == index ? 14'h80 : _GEN_12641;
  wire [13:0] _GEN_12643 = 14'h3163 == index ? 14'h62 : _GEN_12642;
  wire [13:0] _GEN_12644 = 14'h3164 == index ? 14'h62 : _GEN_12643;
  wire [13:0] _GEN_12645 = 14'h3165 == index ? 14'h62 : _GEN_12644;
  wire [13:0] _GEN_12646 = 14'h3166 == index ? 14'h62 : _GEN_12645;
  wire [13:0] _GEN_12647 = 14'h3167 == index ? 14'h62 : _GEN_12646;
  wire [13:0] _GEN_12648 = 14'h3168 == index ? 14'h62 : _GEN_12647;
  wire [13:0] _GEN_12649 = 14'h3169 == index ? 14'h62 : _GEN_12648;
  wire [13:0] _GEN_12650 = 14'h316a == index ? 14'h62 : _GEN_12649;
  wire [13:0] _GEN_12651 = 14'h316b == index ? 14'h62 : _GEN_12650;
  wire [13:0] _GEN_12652 = 14'h316c == index ? 14'h62 : _GEN_12651;
  wire [13:0] _GEN_12653 = 14'h316d == index ? 14'h62 : _GEN_12652;
  wire [13:0] _GEN_12654 = 14'h316e == index ? 14'h62 : _GEN_12653;
  wire [13:0] _GEN_12655 = 14'h316f == index ? 14'h62 : _GEN_12654;
  wire [13:0] _GEN_12656 = 14'h3170 == index ? 14'h62 : _GEN_12655;
  wire [13:0] _GEN_12657 = 14'h3171 == index ? 14'h62 : _GEN_12656;
  wire [13:0] _GEN_12658 = 14'h3172 == index ? 14'h62 : _GEN_12657;
  wire [13:0] _GEN_12659 = 14'h3173 == index ? 14'h62 : _GEN_12658;
  wire [13:0] _GEN_12660 = 14'h3174 == index ? 14'h62 : _GEN_12659;
  wire [13:0] _GEN_12661 = 14'h3175 == index ? 14'h62 : _GEN_12660;
  wire [13:0] _GEN_12662 = 14'h3176 == index ? 14'h62 : _GEN_12661;
  wire [13:0] _GEN_12663 = 14'h3177 == index ? 14'h62 : _GEN_12662;
  wire [13:0] _GEN_12664 = 14'h3178 == index ? 14'h62 : _GEN_12663;
  wire [13:0] _GEN_12665 = 14'h3179 == index ? 14'h62 : _GEN_12664;
  wire [13:0] _GEN_12666 = 14'h317a == index ? 14'h62 : _GEN_12665;
  wire [13:0] _GEN_12667 = 14'h317b == index ? 14'h62 : _GEN_12666;
  wire [13:0] _GEN_12668 = 14'h317c == index ? 14'h62 : _GEN_12667;
  wire [13:0] _GEN_12669 = 14'h317d == index ? 14'h62 : _GEN_12668;
  wire [13:0] _GEN_12670 = 14'h317e == index ? 14'h62 : _GEN_12669;
  wire [13:0] _GEN_12671 = 14'h317f == index ? 14'h62 : _GEN_12670;
  wire [13:0] _GEN_12672 = 14'h3180 == index ? 14'h0 : _GEN_12671;
  wire [13:0] _GEN_12673 = 14'h3181 == index ? 14'h3180 : _GEN_12672;
  wire [13:0] _GEN_12674 = 14'h3182 == index ? 14'h1881 : _GEN_12673;
  wire [13:0] _GEN_12675 = 14'h3183 == index ? 14'h1080 : _GEN_12674;
  wire [13:0] _GEN_12676 = 14'h3184 == index ? 14'hc03 : _GEN_12675;
  wire [13:0] _GEN_12677 = 14'h3185 == index ? 14'h984 : _GEN_12676;
  wire [13:0] _GEN_12678 = 14'h3186 == index ? 14'h803 : _GEN_12677;
  wire [13:0] _GEN_12679 = 14'h3187 == index ? 14'h701 : _GEN_12678;
  wire [13:0] _GEN_12680 = 14'h3188 == index ? 14'h603 : _GEN_12679;
  wire [13:0] _GEN_12681 = 14'h3189 == index ? 14'h580 : _GEN_12680;
  wire [13:0] _GEN_12682 = 14'h318a == index ? 14'h489 : _GEN_12681;
  wire [13:0] _GEN_12683 = 14'h318b == index ? 14'h480 : _GEN_12682;
  wire [13:0] _GEN_12684 = 14'h318c == index ? 14'h403 : _GEN_12683;
  wire [13:0] _GEN_12685 = 14'h318d == index ? 14'h388 : _GEN_12684;
  wire [13:0] _GEN_12686 = 14'h318e == index ? 14'h381 : _GEN_12685;
  wire [13:0] _GEN_12687 = 14'h318f == index ? 14'h309 : _GEN_12686;
  wire [13:0] _GEN_12688 = 14'h3190 == index ? 14'h303 : _GEN_12687;
  wire [13:0] _GEN_12689 = 14'h3191 == index ? 14'h28e : _GEN_12688;
  wire [13:0] _GEN_12690 = 14'h3192 == index ? 14'h289 : _GEN_12689;
  wire [13:0] _GEN_12691 = 14'h3193 == index ? 14'h284 : _GEN_12690;
  wire [13:0] _GEN_12692 = 14'h3194 == index ? 14'h213 : _GEN_12691;
  wire [13:0] _GEN_12693 = 14'h3195 == index ? 14'h20f : _GEN_12692;
  wire [13:0] _GEN_12694 = 14'h3196 == index ? 14'h20b : _GEN_12693;
  wire [13:0] _GEN_12695 = 14'h3197 == index ? 14'h207 : _GEN_12694;
  wire [13:0] _GEN_12696 = 14'h3198 == index ? 14'h203 : _GEN_12695;
  wire [13:0] _GEN_12697 = 14'h3199 == index ? 14'h198 : _GEN_12696;
  wire [13:0] _GEN_12698 = 14'h319a == index ? 14'h195 : _GEN_12697;
  wire [13:0] _GEN_12699 = 14'h319b == index ? 14'h192 : _GEN_12698;
  wire [13:0] _GEN_12700 = 14'h319c == index ? 14'h18f : _GEN_12699;
  wire [13:0] _GEN_12701 = 14'h319d == index ? 14'h18c : _GEN_12700;
  wire [13:0] _GEN_12702 = 14'h319e == index ? 14'h189 : _GEN_12701;
  wire [13:0] _GEN_12703 = 14'h319f == index ? 14'h186 : _GEN_12702;
  wire [13:0] _GEN_12704 = 14'h31a0 == index ? 14'h183 : _GEN_12703;
  wire [13:0] _GEN_12705 = 14'h31a1 == index ? 14'h180 : _GEN_12704;
  wire [13:0] _GEN_12706 = 14'h31a2 == index ? 14'h11f : _GEN_12705;
  wire [13:0] _GEN_12707 = 14'h31a3 == index ? 14'h11d : _GEN_12706;
  wire [13:0] _GEN_12708 = 14'h31a4 == index ? 14'h11b : _GEN_12707;
  wire [13:0] _GEN_12709 = 14'h31a5 == index ? 14'h119 : _GEN_12708;
  wire [13:0] _GEN_12710 = 14'h31a6 == index ? 14'h117 : _GEN_12709;
  wire [13:0] _GEN_12711 = 14'h31a7 == index ? 14'h115 : _GEN_12710;
  wire [13:0] _GEN_12712 = 14'h31a8 == index ? 14'h113 : _GEN_12711;
  wire [13:0] _GEN_12713 = 14'h31a9 == index ? 14'h111 : _GEN_12712;
  wire [13:0] _GEN_12714 = 14'h31aa == index ? 14'h10f : _GEN_12713;
  wire [13:0] _GEN_12715 = 14'h31ab == index ? 14'h10d : _GEN_12714;
  wire [13:0] _GEN_12716 = 14'h31ac == index ? 14'h10b : _GEN_12715;
  wire [13:0] _GEN_12717 = 14'h31ad == index ? 14'h109 : _GEN_12716;
  wire [13:0] _GEN_12718 = 14'h31ae == index ? 14'h107 : _GEN_12717;
  wire [13:0] _GEN_12719 = 14'h31af == index ? 14'h105 : _GEN_12718;
  wire [13:0] _GEN_12720 = 14'h31b0 == index ? 14'h103 : _GEN_12719;
  wire [13:0] _GEN_12721 = 14'h31b1 == index ? 14'h101 : _GEN_12720;
  wire [13:0] _GEN_12722 = 14'h31b2 == index ? 14'hb1 : _GEN_12721;
  wire [13:0] _GEN_12723 = 14'h31b3 == index ? 14'hb0 : _GEN_12722;
  wire [13:0] _GEN_12724 = 14'h31b4 == index ? 14'haf : _GEN_12723;
  wire [13:0] _GEN_12725 = 14'h31b5 == index ? 14'hae : _GEN_12724;
  wire [13:0] _GEN_12726 = 14'h31b6 == index ? 14'had : _GEN_12725;
  wire [13:0] _GEN_12727 = 14'h31b7 == index ? 14'hac : _GEN_12726;
  wire [13:0] _GEN_12728 = 14'h31b8 == index ? 14'hab : _GEN_12727;
  wire [13:0] _GEN_12729 = 14'h31b9 == index ? 14'haa : _GEN_12728;
  wire [13:0] _GEN_12730 = 14'h31ba == index ? 14'ha9 : _GEN_12729;
  wire [13:0] _GEN_12731 = 14'h31bb == index ? 14'ha8 : _GEN_12730;
  wire [13:0] _GEN_12732 = 14'h31bc == index ? 14'ha7 : _GEN_12731;
  wire [13:0] _GEN_12733 = 14'h31bd == index ? 14'ha6 : _GEN_12732;
  wire [13:0] _GEN_12734 = 14'h31be == index ? 14'ha5 : _GEN_12733;
  wire [13:0] _GEN_12735 = 14'h31bf == index ? 14'ha4 : _GEN_12734;
  wire [13:0] _GEN_12736 = 14'h31c0 == index ? 14'ha3 : _GEN_12735;
  wire [13:0] _GEN_12737 = 14'h31c1 == index ? 14'ha2 : _GEN_12736;
  wire [13:0] _GEN_12738 = 14'h31c2 == index ? 14'ha1 : _GEN_12737;
  wire [13:0] _GEN_12739 = 14'h31c3 == index ? 14'ha0 : _GEN_12738;
  wire [13:0] _GEN_12740 = 14'h31c4 == index ? 14'h9f : _GEN_12739;
  wire [13:0] _GEN_12741 = 14'h31c5 == index ? 14'h9e : _GEN_12740;
  wire [13:0] _GEN_12742 = 14'h31c6 == index ? 14'h9d : _GEN_12741;
  wire [13:0] _GEN_12743 = 14'h31c7 == index ? 14'h9c : _GEN_12742;
  wire [13:0] _GEN_12744 = 14'h31c8 == index ? 14'h9b : _GEN_12743;
  wire [13:0] _GEN_12745 = 14'h31c9 == index ? 14'h9a : _GEN_12744;
  wire [13:0] _GEN_12746 = 14'h31ca == index ? 14'h99 : _GEN_12745;
  wire [13:0] _GEN_12747 = 14'h31cb == index ? 14'h98 : _GEN_12746;
  wire [13:0] _GEN_12748 = 14'h31cc == index ? 14'h97 : _GEN_12747;
  wire [13:0] _GEN_12749 = 14'h31cd == index ? 14'h96 : _GEN_12748;
  wire [13:0] _GEN_12750 = 14'h31ce == index ? 14'h95 : _GEN_12749;
  wire [13:0] _GEN_12751 = 14'h31cf == index ? 14'h94 : _GEN_12750;
  wire [13:0] _GEN_12752 = 14'h31d0 == index ? 14'h93 : _GEN_12751;
  wire [13:0] _GEN_12753 = 14'h31d1 == index ? 14'h92 : _GEN_12752;
  wire [13:0] _GEN_12754 = 14'h31d2 == index ? 14'h91 : _GEN_12753;
  wire [13:0] _GEN_12755 = 14'h31d3 == index ? 14'h90 : _GEN_12754;
  wire [13:0] _GEN_12756 = 14'h31d4 == index ? 14'h8f : _GEN_12755;
  wire [13:0] _GEN_12757 = 14'h31d5 == index ? 14'h8e : _GEN_12756;
  wire [13:0] _GEN_12758 = 14'h31d6 == index ? 14'h8d : _GEN_12757;
  wire [13:0] _GEN_12759 = 14'h31d7 == index ? 14'h8c : _GEN_12758;
  wire [13:0] _GEN_12760 = 14'h31d8 == index ? 14'h8b : _GEN_12759;
  wire [13:0] _GEN_12761 = 14'h31d9 == index ? 14'h8a : _GEN_12760;
  wire [13:0] _GEN_12762 = 14'h31da == index ? 14'h89 : _GEN_12761;
  wire [13:0] _GEN_12763 = 14'h31db == index ? 14'h88 : _GEN_12762;
  wire [13:0] _GEN_12764 = 14'h31dc == index ? 14'h87 : _GEN_12763;
  wire [13:0] _GEN_12765 = 14'h31dd == index ? 14'h86 : _GEN_12764;
  wire [13:0] _GEN_12766 = 14'h31de == index ? 14'h85 : _GEN_12765;
  wire [13:0] _GEN_12767 = 14'h31df == index ? 14'h84 : _GEN_12766;
  wire [13:0] _GEN_12768 = 14'h31e0 == index ? 14'h83 : _GEN_12767;
  wire [13:0] _GEN_12769 = 14'h31e1 == index ? 14'h82 : _GEN_12768;
  wire [13:0] _GEN_12770 = 14'h31e2 == index ? 14'h81 : _GEN_12769;
  wire [13:0] _GEN_12771 = 14'h31e3 == index ? 14'h80 : _GEN_12770;
  wire [13:0] _GEN_12772 = 14'h31e4 == index ? 14'h63 : _GEN_12771;
  wire [13:0] _GEN_12773 = 14'h31e5 == index ? 14'h63 : _GEN_12772;
  wire [13:0] _GEN_12774 = 14'h31e6 == index ? 14'h63 : _GEN_12773;
  wire [13:0] _GEN_12775 = 14'h31e7 == index ? 14'h63 : _GEN_12774;
  wire [13:0] _GEN_12776 = 14'h31e8 == index ? 14'h63 : _GEN_12775;
  wire [13:0] _GEN_12777 = 14'h31e9 == index ? 14'h63 : _GEN_12776;
  wire [13:0] _GEN_12778 = 14'h31ea == index ? 14'h63 : _GEN_12777;
  wire [13:0] _GEN_12779 = 14'h31eb == index ? 14'h63 : _GEN_12778;
  wire [13:0] _GEN_12780 = 14'h31ec == index ? 14'h63 : _GEN_12779;
  wire [13:0] _GEN_12781 = 14'h31ed == index ? 14'h63 : _GEN_12780;
  wire [13:0] _GEN_12782 = 14'h31ee == index ? 14'h63 : _GEN_12781;
  wire [13:0] _GEN_12783 = 14'h31ef == index ? 14'h63 : _GEN_12782;
  wire [13:0] _GEN_12784 = 14'h31f0 == index ? 14'h63 : _GEN_12783;
  wire [13:0] _GEN_12785 = 14'h31f1 == index ? 14'h63 : _GEN_12784;
  wire [13:0] _GEN_12786 = 14'h31f2 == index ? 14'h63 : _GEN_12785;
  wire [13:0] _GEN_12787 = 14'h31f3 == index ? 14'h63 : _GEN_12786;
  wire [13:0] _GEN_12788 = 14'h31f4 == index ? 14'h63 : _GEN_12787;
  wire [13:0] _GEN_12789 = 14'h31f5 == index ? 14'h63 : _GEN_12788;
  wire [13:0] _GEN_12790 = 14'h31f6 == index ? 14'h63 : _GEN_12789;
  wire [13:0] _GEN_12791 = 14'h31f7 == index ? 14'h63 : _GEN_12790;
  wire [13:0] _GEN_12792 = 14'h31f8 == index ? 14'h63 : _GEN_12791;
  wire [13:0] _GEN_12793 = 14'h31f9 == index ? 14'h63 : _GEN_12792;
  wire [13:0] _GEN_12794 = 14'h31fa == index ? 14'h63 : _GEN_12793;
  wire [13:0] _GEN_12795 = 14'h31fb == index ? 14'h63 : _GEN_12794;
  wire [13:0] _GEN_12796 = 14'h31fc == index ? 14'h63 : _GEN_12795;
  wire [13:0] _GEN_12797 = 14'h31fd == index ? 14'h63 : _GEN_12796;
  wire [13:0] _GEN_12798 = 14'h31fe == index ? 14'h63 : _GEN_12797;
  wire [13:0] _GEN_12799 = 14'h31ff == index ? 14'h63 : _GEN_12798;
  wire [13:0] _GEN_12800 = 14'h3200 == index ? 14'h0 : _GEN_12799;
  wire [13:0] _GEN_12801 = 14'h3201 == index ? 14'h3200 : _GEN_12800;
  wire [13:0] _GEN_12802 = 14'h3202 == index ? 14'h1900 : _GEN_12801;
  wire [13:0] _GEN_12803 = 14'h3203 == index ? 14'h1081 : _GEN_12802;
  wire [13:0] _GEN_12804 = 14'h3204 == index ? 14'hc80 : _GEN_12803;
  wire [13:0] _GEN_12805 = 14'h3205 == index ? 14'ha00 : _GEN_12804;
  wire [13:0] _GEN_12806 = 14'h3206 == index ? 14'h804 : _GEN_12805;
  wire [13:0] _GEN_12807 = 14'h3207 == index ? 14'h702 : _GEN_12806;
  wire [13:0] _GEN_12808 = 14'h3208 == index ? 14'h604 : _GEN_12807;
  wire [13:0] _GEN_12809 = 14'h3209 == index ? 14'h581 : _GEN_12808;
  wire [13:0] _GEN_12810 = 14'h320a == index ? 14'h500 : _GEN_12809;
  wire [13:0] _GEN_12811 = 14'h320b == index ? 14'h481 : _GEN_12810;
  wire [13:0] _GEN_12812 = 14'h320c == index ? 14'h404 : _GEN_12811;
  wire [13:0] _GEN_12813 = 14'h320d == index ? 14'h389 : _GEN_12812;
  wire [13:0] _GEN_12814 = 14'h320e == index ? 14'h382 : _GEN_12813;
  wire [13:0] _GEN_12815 = 14'h320f == index ? 14'h30a : _GEN_12814;
  wire [13:0] _GEN_12816 = 14'h3210 == index ? 14'h304 : _GEN_12815;
  wire [13:0] _GEN_12817 = 14'h3211 == index ? 14'h28f : _GEN_12816;
  wire [13:0] _GEN_12818 = 14'h3212 == index ? 14'h28a : _GEN_12817;
  wire [13:0] _GEN_12819 = 14'h3213 == index ? 14'h285 : _GEN_12818;
  wire [13:0] _GEN_12820 = 14'h3214 == index ? 14'h280 : _GEN_12819;
  wire [13:0] _GEN_12821 = 14'h3215 == index ? 14'h210 : _GEN_12820;
  wire [13:0] _GEN_12822 = 14'h3216 == index ? 14'h20c : _GEN_12821;
  wire [13:0] _GEN_12823 = 14'h3217 == index ? 14'h208 : _GEN_12822;
  wire [13:0] _GEN_12824 = 14'h3218 == index ? 14'h204 : _GEN_12823;
  wire [13:0] _GEN_12825 = 14'h3219 == index ? 14'h200 : _GEN_12824;
  wire [13:0] _GEN_12826 = 14'h321a == index ? 14'h196 : _GEN_12825;
  wire [13:0] _GEN_12827 = 14'h321b == index ? 14'h193 : _GEN_12826;
  wire [13:0] _GEN_12828 = 14'h321c == index ? 14'h190 : _GEN_12827;
  wire [13:0] _GEN_12829 = 14'h321d == index ? 14'h18d : _GEN_12828;
  wire [13:0] _GEN_12830 = 14'h321e == index ? 14'h18a : _GEN_12829;
  wire [13:0] _GEN_12831 = 14'h321f == index ? 14'h187 : _GEN_12830;
  wire [13:0] _GEN_12832 = 14'h3220 == index ? 14'h184 : _GEN_12831;
  wire [13:0] _GEN_12833 = 14'h3221 == index ? 14'h181 : _GEN_12832;
  wire [13:0] _GEN_12834 = 14'h3222 == index ? 14'h120 : _GEN_12833;
  wire [13:0] _GEN_12835 = 14'h3223 == index ? 14'h11e : _GEN_12834;
  wire [13:0] _GEN_12836 = 14'h3224 == index ? 14'h11c : _GEN_12835;
  wire [13:0] _GEN_12837 = 14'h3225 == index ? 14'h11a : _GEN_12836;
  wire [13:0] _GEN_12838 = 14'h3226 == index ? 14'h118 : _GEN_12837;
  wire [13:0] _GEN_12839 = 14'h3227 == index ? 14'h116 : _GEN_12838;
  wire [13:0] _GEN_12840 = 14'h3228 == index ? 14'h114 : _GEN_12839;
  wire [13:0] _GEN_12841 = 14'h3229 == index ? 14'h112 : _GEN_12840;
  wire [13:0] _GEN_12842 = 14'h322a == index ? 14'h110 : _GEN_12841;
  wire [13:0] _GEN_12843 = 14'h322b == index ? 14'h10e : _GEN_12842;
  wire [13:0] _GEN_12844 = 14'h322c == index ? 14'h10c : _GEN_12843;
  wire [13:0] _GEN_12845 = 14'h322d == index ? 14'h10a : _GEN_12844;
  wire [13:0] _GEN_12846 = 14'h322e == index ? 14'h108 : _GEN_12845;
  wire [13:0] _GEN_12847 = 14'h322f == index ? 14'h106 : _GEN_12846;
  wire [13:0] _GEN_12848 = 14'h3230 == index ? 14'h104 : _GEN_12847;
  wire [13:0] _GEN_12849 = 14'h3231 == index ? 14'h102 : _GEN_12848;
  wire [13:0] _GEN_12850 = 14'h3232 == index ? 14'h100 : _GEN_12849;
  wire [13:0] _GEN_12851 = 14'h3233 == index ? 14'hb1 : _GEN_12850;
  wire [13:0] _GEN_12852 = 14'h3234 == index ? 14'hb0 : _GEN_12851;
  wire [13:0] _GEN_12853 = 14'h3235 == index ? 14'haf : _GEN_12852;
  wire [13:0] _GEN_12854 = 14'h3236 == index ? 14'hae : _GEN_12853;
  wire [13:0] _GEN_12855 = 14'h3237 == index ? 14'had : _GEN_12854;
  wire [13:0] _GEN_12856 = 14'h3238 == index ? 14'hac : _GEN_12855;
  wire [13:0] _GEN_12857 = 14'h3239 == index ? 14'hab : _GEN_12856;
  wire [13:0] _GEN_12858 = 14'h323a == index ? 14'haa : _GEN_12857;
  wire [13:0] _GEN_12859 = 14'h323b == index ? 14'ha9 : _GEN_12858;
  wire [13:0] _GEN_12860 = 14'h323c == index ? 14'ha8 : _GEN_12859;
  wire [13:0] _GEN_12861 = 14'h323d == index ? 14'ha7 : _GEN_12860;
  wire [13:0] _GEN_12862 = 14'h323e == index ? 14'ha6 : _GEN_12861;
  wire [13:0] _GEN_12863 = 14'h323f == index ? 14'ha5 : _GEN_12862;
  wire [13:0] _GEN_12864 = 14'h3240 == index ? 14'ha4 : _GEN_12863;
  wire [13:0] _GEN_12865 = 14'h3241 == index ? 14'ha3 : _GEN_12864;
  wire [13:0] _GEN_12866 = 14'h3242 == index ? 14'ha2 : _GEN_12865;
  wire [13:0] _GEN_12867 = 14'h3243 == index ? 14'ha1 : _GEN_12866;
  wire [13:0] _GEN_12868 = 14'h3244 == index ? 14'ha0 : _GEN_12867;
  wire [13:0] _GEN_12869 = 14'h3245 == index ? 14'h9f : _GEN_12868;
  wire [13:0] _GEN_12870 = 14'h3246 == index ? 14'h9e : _GEN_12869;
  wire [13:0] _GEN_12871 = 14'h3247 == index ? 14'h9d : _GEN_12870;
  wire [13:0] _GEN_12872 = 14'h3248 == index ? 14'h9c : _GEN_12871;
  wire [13:0] _GEN_12873 = 14'h3249 == index ? 14'h9b : _GEN_12872;
  wire [13:0] _GEN_12874 = 14'h324a == index ? 14'h9a : _GEN_12873;
  wire [13:0] _GEN_12875 = 14'h324b == index ? 14'h99 : _GEN_12874;
  wire [13:0] _GEN_12876 = 14'h324c == index ? 14'h98 : _GEN_12875;
  wire [13:0] _GEN_12877 = 14'h324d == index ? 14'h97 : _GEN_12876;
  wire [13:0] _GEN_12878 = 14'h324e == index ? 14'h96 : _GEN_12877;
  wire [13:0] _GEN_12879 = 14'h324f == index ? 14'h95 : _GEN_12878;
  wire [13:0] _GEN_12880 = 14'h3250 == index ? 14'h94 : _GEN_12879;
  wire [13:0] _GEN_12881 = 14'h3251 == index ? 14'h93 : _GEN_12880;
  wire [13:0] _GEN_12882 = 14'h3252 == index ? 14'h92 : _GEN_12881;
  wire [13:0] _GEN_12883 = 14'h3253 == index ? 14'h91 : _GEN_12882;
  wire [13:0] _GEN_12884 = 14'h3254 == index ? 14'h90 : _GEN_12883;
  wire [13:0] _GEN_12885 = 14'h3255 == index ? 14'h8f : _GEN_12884;
  wire [13:0] _GEN_12886 = 14'h3256 == index ? 14'h8e : _GEN_12885;
  wire [13:0] _GEN_12887 = 14'h3257 == index ? 14'h8d : _GEN_12886;
  wire [13:0] _GEN_12888 = 14'h3258 == index ? 14'h8c : _GEN_12887;
  wire [13:0] _GEN_12889 = 14'h3259 == index ? 14'h8b : _GEN_12888;
  wire [13:0] _GEN_12890 = 14'h325a == index ? 14'h8a : _GEN_12889;
  wire [13:0] _GEN_12891 = 14'h325b == index ? 14'h89 : _GEN_12890;
  wire [13:0] _GEN_12892 = 14'h325c == index ? 14'h88 : _GEN_12891;
  wire [13:0] _GEN_12893 = 14'h325d == index ? 14'h87 : _GEN_12892;
  wire [13:0] _GEN_12894 = 14'h325e == index ? 14'h86 : _GEN_12893;
  wire [13:0] _GEN_12895 = 14'h325f == index ? 14'h85 : _GEN_12894;
  wire [13:0] _GEN_12896 = 14'h3260 == index ? 14'h84 : _GEN_12895;
  wire [13:0] _GEN_12897 = 14'h3261 == index ? 14'h83 : _GEN_12896;
  wire [13:0] _GEN_12898 = 14'h3262 == index ? 14'h82 : _GEN_12897;
  wire [13:0] _GEN_12899 = 14'h3263 == index ? 14'h81 : _GEN_12898;
  wire [13:0] _GEN_12900 = 14'h3264 == index ? 14'h80 : _GEN_12899;
  wire [13:0] _GEN_12901 = 14'h3265 == index ? 14'h64 : _GEN_12900;
  wire [13:0] _GEN_12902 = 14'h3266 == index ? 14'h64 : _GEN_12901;
  wire [13:0] _GEN_12903 = 14'h3267 == index ? 14'h64 : _GEN_12902;
  wire [13:0] _GEN_12904 = 14'h3268 == index ? 14'h64 : _GEN_12903;
  wire [13:0] _GEN_12905 = 14'h3269 == index ? 14'h64 : _GEN_12904;
  wire [13:0] _GEN_12906 = 14'h326a == index ? 14'h64 : _GEN_12905;
  wire [13:0] _GEN_12907 = 14'h326b == index ? 14'h64 : _GEN_12906;
  wire [13:0] _GEN_12908 = 14'h326c == index ? 14'h64 : _GEN_12907;
  wire [13:0] _GEN_12909 = 14'h326d == index ? 14'h64 : _GEN_12908;
  wire [13:0] _GEN_12910 = 14'h326e == index ? 14'h64 : _GEN_12909;
  wire [13:0] _GEN_12911 = 14'h326f == index ? 14'h64 : _GEN_12910;
  wire [13:0] _GEN_12912 = 14'h3270 == index ? 14'h64 : _GEN_12911;
  wire [13:0] _GEN_12913 = 14'h3271 == index ? 14'h64 : _GEN_12912;
  wire [13:0] _GEN_12914 = 14'h3272 == index ? 14'h64 : _GEN_12913;
  wire [13:0] _GEN_12915 = 14'h3273 == index ? 14'h64 : _GEN_12914;
  wire [13:0] _GEN_12916 = 14'h3274 == index ? 14'h64 : _GEN_12915;
  wire [13:0] _GEN_12917 = 14'h3275 == index ? 14'h64 : _GEN_12916;
  wire [13:0] _GEN_12918 = 14'h3276 == index ? 14'h64 : _GEN_12917;
  wire [13:0] _GEN_12919 = 14'h3277 == index ? 14'h64 : _GEN_12918;
  wire [13:0] _GEN_12920 = 14'h3278 == index ? 14'h64 : _GEN_12919;
  wire [13:0] _GEN_12921 = 14'h3279 == index ? 14'h64 : _GEN_12920;
  wire [13:0] _GEN_12922 = 14'h327a == index ? 14'h64 : _GEN_12921;
  wire [13:0] _GEN_12923 = 14'h327b == index ? 14'h64 : _GEN_12922;
  wire [13:0] _GEN_12924 = 14'h327c == index ? 14'h64 : _GEN_12923;
  wire [13:0] _GEN_12925 = 14'h327d == index ? 14'h64 : _GEN_12924;
  wire [13:0] _GEN_12926 = 14'h327e == index ? 14'h64 : _GEN_12925;
  wire [13:0] _GEN_12927 = 14'h327f == index ? 14'h64 : _GEN_12926;
  wire [13:0] _GEN_12928 = 14'h3280 == index ? 14'h0 : _GEN_12927;
  wire [13:0] _GEN_12929 = 14'h3281 == index ? 14'h3280 : _GEN_12928;
  wire [13:0] _GEN_12930 = 14'h3282 == index ? 14'h1901 : _GEN_12929;
  wire [13:0] _GEN_12931 = 14'h3283 == index ? 14'h1082 : _GEN_12930;
  wire [13:0] _GEN_12932 = 14'h3284 == index ? 14'hc81 : _GEN_12931;
  wire [13:0] _GEN_12933 = 14'h3285 == index ? 14'ha01 : _GEN_12932;
  wire [13:0] _GEN_12934 = 14'h3286 == index ? 14'h805 : _GEN_12933;
  wire [13:0] _GEN_12935 = 14'h3287 == index ? 14'h703 : _GEN_12934;
  wire [13:0] _GEN_12936 = 14'h3288 == index ? 14'h605 : _GEN_12935;
  wire [13:0] _GEN_12937 = 14'h3289 == index ? 14'h582 : _GEN_12936;
  wire [13:0] _GEN_12938 = 14'h328a == index ? 14'h501 : _GEN_12937;
  wire [13:0] _GEN_12939 = 14'h328b == index ? 14'h482 : _GEN_12938;
  wire [13:0] _GEN_12940 = 14'h328c == index ? 14'h405 : _GEN_12939;
  wire [13:0] _GEN_12941 = 14'h328d == index ? 14'h38a : _GEN_12940;
  wire [13:0] _GEN_12942 = 14'h328e == index ? 14'h383 : _GEN_12941;
  wire [13:0] _GEN_12943 = 14'h328f == index ? 14'h30b : _GEN_12942;
  wire [13:0] _GEN_12944 = 14'h3290 == index ? 14'h305 : _GEN_12943;
  wire [13:0] _GEN_12945 = 14'h3291 == index ? 14'h290 : _GEN_12944;
  wire [13:0] _GEN_12946 = 14'h3292 == index ? 14'h28b : _GEN_12945;
  wire [13:0] _GEN_12947 = 14'h3293 == index ? 14'h286 : _GEN_12946;
  wire [13:0] _GEN_12948 = 14'h3294 == index ? 14'h281 : _GEN_12947;
  wire [13:0] _GEN_12949 = 14'h3295 == index ? 14'h211 : _GEN_12948;
  wire [13:0] _GEN_12950 = 14'h3296 == index ? 14'h20d : _GEN_12949;
  wire [13:0] _GEN_12951 = 14'h3297 == index ? 14'h209 : _GEN_12950;
  wire [13:0] _GEN_12952 = 14'h3298 == index ? 14'h205 : _GEN_12951;
  wire [13:0] _GEN_12953 = 14'h3299 == index ? 14'h201 : _GEN_12952;
  wire [13:0] _GEN_12954 = 14'h329a == index ? 14'h197 : _GEN_12953;
  wire [13:0] _GEN_12955 = 14'h329b == index ? 14'h194 : _GEN_12954;
  wire [13:0] _GEN_12956 = 14'h329c == index ? 14'h191 : _GEN_12955;
  wire [13:0] _GEN_12957 = 14'h329d == index ? 14'h18e : _GEN_12956;
  wire [13:0] _GEN_12958 = 14'h329e == index ? 14'h18b : _GEN_12957;
  wire [13:0] _GEN_12959 = 14'h329f == index ? 14'h188 : _GEN_12958;
  wire [13:0] _GEN_12960 = 14'h32a0 == index ? 14'h185 : _GEN_12959;
  wire [13:0] _GEN_12961 = 14'h32a1 == index ? 14'h182 : _GEN_12960;
  wire [13:0] _GEN_12962 = 14'h32a2 == index ? 14'h121 : _GEN_12961;
  wire [13:0] _GEN_12963 = 14'h32a3 == index ? 14'h11f : _GEN_12962;
  wire [13:0] _GEN_12964 = 14'h32a4 == index ? 14'h11d : _GEN_12963;
  wire [13:0] _GEN_12965 = 14'h32a5 == index ? 14'h11b : _GEN_12964;
  wire [13:0] _GEN_12966 = 14'h32a6 == index ? 14'h119 : _GEN_12965;
  wire [13:0] _GEN_12967 = 14'h32a7 == index ? 14'h117 : _GEN_12966;
  wire [13:0] _GEN_12968 = 14'h32a8 == index ? 14'h115 : _GEN_12967;
  wire [13:0] _GEN_12969 = 14'h32a9 == index ? 14'h113 : _GEN_12968;
  wire [13:0] _GEN_12970 = 14'h32aa == index ? 14'h111 : _GEN_12969;
  wire [13:0] _GEN_12971 = 14'h32ab == index ? 14'h10f : _GEN_12970;
  wire [13:0] _GEN_12972 = 14'h32ac == index ? 14'h10d : _GEN_12971;
  wire [13:0] _GEN_12973 = 14'h32ad == index ? 14'h10b : _GEN_12972;
  wire [13:0] _GEN_12974 = 14'h32ae == index ? 14'h109 : _GEN_12973;
  wire [13:0] _GEN_12975 = 14'h32af == index ? 14'h107 : _GEN_12974;
  wire [13:0] _GEN_12976 = 14'h32b0 == index ? 14'h105 : _GEN_12975;
  wire [13:0] _GEN_12977 = 14'h32b1 == index ? 14'h103 : _GEN_12976;
  wire [13:0] _GEN_12978 = 14'h32b2 == index ? 14'h101 : _GEN_12977;
  wire [13:0] _GEN_12979 = 14'h32b3 == index ? 14'hb2 : _GEN_12978;
  wire [13:0] _GEN_12980 = 14'h32b4 == index ? 14'hb1 : _GEN_12979;
  wire [13:0] _GEN_12981 = 14'h32b5 == index ? 14'hb0 : _GEN_12980;
  wire [13:0] _GEN_12982 = 14'h32b6 == index ? 14'haf : _GEN_12981;
  wire [13:0] _GEN_12983 = 14'h32b7 == index ? 14'hae : _GEN_12982;
  wire [13:0] _GEN_12984 = 14'h32b8 == index ? 14'had : _GEN_12983;
  wire [13:0] _GEN_12985 = 14'h32b9 == index ? 14'hac : _GEN_12984;
  wire [13:0] _GEN_12986 = 14'h32ba == index ? 14'hab : _GEN_12985;
  wire [13:0] _GEN_12987 = 14'h32bb == index ? 14'haa : _GEN_12986;
  wire [13:0] _GEN_12988 = 14'h32bc == index ? 14'ha9 : _GEN_12987;
  wire [13:0] _GEN_12989 = 14'h32bd == index ? 14'ha8 : _GEN_12988;
  wire [13:0] _GEN_12990 = 14'h32be == index ? 14'ha7 : _GEN_12989;
  wire [13:0] _GEN_12991 = 14'h32bf == index ? 14'ha6 : _GEN_12990;
  wire [13:0] _GEN_12992 = 14'h32c0 == index ? 14'ha5 : _GEN_12991;
  wire [13:0] _GEN_12993 = 14'h32c1 == index ? 14'ha4 : _GEN_12992;
  wire [13:0] _GEN_12994 = 14'h32c2 == index ? 14'ha3 : _GEN_12993;
  wire [13:0] _GEN_12995 = 14'h32c3 == index ? 14'ha2 : _GEN_12994;
  wire [13:0] _GEN_12996 = 14'h32c4 == index ? 14'ha1 : _GEN_12995;
  wire [13:0] _GEN_12997 = 14'h32c5 == index ? 14'ha0 : _GEN_12996;
  wire [13:0] _GEN_12998 = 14'h32c6 == index ? 14'h9f : _GEN_12997;
  wire [13:0] _GEN_12999 = 14'h32c7 == index ? 14'h9e : _GEN_12998;
  wire [13:0] _GEN_13000 = 14'h32c8 == index ? 14'h9d : _GEN_12999;
  wire [13:0] _GEN_13001 = 14'h32c9 == index ? 14'h9c : _GEN_13000;
  wire [13:0] _GEN_13002 = 14'h32ca == index ? 14'h9b : _GEN_13001;
  wire [13:0] _GEN_13003 = 14'h32cb == index ? 14'h9a : _GEN_13002;
  wire [13:0] _GEN_13004 = 14'h32cc == index ? 14'h99 : _GEN_13003;
  wire [13:0] _GEN_13005 = 14'h32cd == index ? 14'h98 : _GEN_13004;
  wire [13:0] _GEN_13006 = 14'h32ce == index ? 14'h97 : _GEN_13005;
  wire [13:0] _GEN_13007 = 14'h32cf == index ? 14'h96 : _GEN_13006;
  wire [13:0] _GEN_13008 = 14'h32d0 == index ? 14'h95 : _GEN_13007;
  wire [13:0] _GEN_13009 = 14'h32d1 == index ? 14'h94 : _GEN_13008;
  wire [13:0] _GEN_13010 = 14'h32d2 == index ? 14'h93 : _GEN_13009;
  wire [13:0] _GEN_13011 = 14'h32d3 == index ? 14'h92 : _GEN_13010;
  wire [13:0] _GEN_13012 = 14'h32d4 == index ? 14'h91 : _GEN_13011;
  wire [13:0] _GEN_13013 = 14'h32d5 == index ? 14'h90 : _GEN_13012;
  wire [13:0] _GEN_13014 = 14'h32d6 == index ? 14'h8f : _GEN_13013;
  wire [13:0] _GEN_13015 = 14'h32d7 == index ? 14'h8e : _GEN_13014;
  wire [13:0] _GEN_13016 = 14'h32d8 == index ? 14'h8d : _GEN_13015;
  wire [13:0] _GEN_13017 = 14'h32d9 == index ? 14'h8c : _GEN_13016;
  wire [13:0] _GEN_13018 = 14'h32da == index ? 14'h8b : _GEN_13017;
  wire [13:0] _GEN_13019 = 14'h32db == index ? 14'h8a : _GEN_13018;
  wire [13:0] _GEN_13020 = 14'h32dc == index ? 14'h89 : _GEN_13019;
  wire [13:0] _GEN_13021 = 14'h32dd == index ? 14'h88 : _GEN_13020;
  wire [13:0] _GEN_13022 = 14'h32de == index ? 14'h87 : _GEN_13021;
  wire [13:0] _GEN_13023 = 14'h32df == index ? 14'h86 : _GEN_13022;
  wire [13:0] _GEN_13024 = 14'h32e0 == index ? 14'h85 : _GEN_13023;
  wire [13:0] _GEN_13025 = 14'h32e1 == index ? 14'h84 : _GEN_13024;
  wire [13:0] _GEN_13026 = 14'h32e2 == index ? 14'h83 : _GEN_13025;
  wire [13:0] _GEN_13027 = 14'h32e3 == index ? 14'h82 : _GEN_13026;
  wire [13:0] _GEN_13028 = 14'h32e4 == index ? 14'h81 : _GEN_13027;
  wire [13:0] _GEN_13029 = 14'h32e5 == index ? 14'h80 : _GEN_13028;
  wire [13:0] _GEN_13030 = 14'h32e6 == index ? 14'h65 : _GEN_13029;
  wire [13:0] _GEN_13031 = 14'h32e7 == index ? 14'h65 : _GEN_13030;
  wire [13:0] _GEN_13032 = 14'h32e8 == index ? 14'h65 : _GEN_13031;
  wire [13:0] _GEN_13033 = 14'h32e9 == index ? 14'h65 : _GEN_13032;
  wire [13:0] _GEN_13034 = 14'h32ea == index ? 14'h65 : _GEN_13033;
  wire [13:0] _GEN_13035 = 14'h32eb == index ? 14'h65 : _GEN_13034;
  wire [13:0] _GEN_13036 = 14'h32ec == index ? 14'h65 : _GEN_13035;
  wire [13:0] _GEN_13037 = 14'h32ed == index ? 14'h65 : _GEN_13036;
  wire [13:0] _GEN_13038 = 14'h32ee == index ? 14'h65 : _GEN_13037;
  wire [13:0] _GEN_13039 = 14'h32ef == index ? 14'h65 : _GEN_13038;
  wire [13:0] _GEN_13040 = 14'h32f0 == index ? 14'h65 : _GEN_13039;
  wire [13:0] _GEN_13041 = 14'h32f1 == index ? 14'h65 : _GEN_13040;
  wire [13:0] _GEN_13042 = 14'h32f2 == index ? 14'h65 : _GEN_13041;
  wire [13:0] _GEN_13043 = 14'h32f3 == index ? 14'h65 : _GEN_13042;
  wire [13:0] _GEN_13044 = 14'h32f4 == index ? 14'h65 : _GEN_13043;
  wire [13:0] _GEN_13045 = 14'h32f5 == index ? 14'h65 : _GEN_13044;
  wire [13:0] _GEN_13046 = 14'h32f6 == index ? 14'h65 : _GEN_13045;
  wire [13:0] _GEN_13047 = 14'h32f7 == index ? 14'h65 : _GEN_13046;
  wire [13:0] _GEN_13048 = 14'h32f8 == index ? 14'h65 : _GEN_13047;
  wire [13:0] _GEN_13049 = 14'h32f9 == index ? 14'h65 : _GEN_13048;
  wire [13:0] _GEN_13050 = 14'h32fa == index ? 14'h65 : _GEN_13049;
  wire [13:0] _GEN_13051 = 14'h32fb == index ? 14'h65 : _GEN_13050;
  wire [13:0] _GEN_13052 = 14'h32fc == index ? 14'h65 : _GEN_13051;
  wire [13:0] _GEN_13053 = 14'h32fd == index ? 14'h65 : _GEN_13052;
  wire [13:0] _GEN_13054 = 14'h32fe == index ? 14'h65 : _GEN_13053;
  wire [13:0] _GEN_13055 = 14'h32ff == index ? 14'h65 : _GEN_13054;
  wire [13:0] _GEN_13056 = 14'h3300 == index ? 14'h0 : _GEN_13055;
  wire [13:0] _GEN_13057 = 14'h3301 == index ? 14'h3300 : _GEN_13056;
  wire [13:0] _GEN_13058 = 14'h3302 == index ? 14'h1980 : _GEN_13057;
  wire [13:0] _GEN_13059 = 14'h3303 == index ? 14'h1100 : _GEN_13058;
  wire [13:0] _GEN_13060 = 14'h3304 == index ? 14'hc82 : _GEN_13059;
  wire [13:0] _GEN_13061 = 14'h3305 == index ? 14'ha02 : _GEN_13060;
  wire [13:0] _GEN_13062 = 14'h3306 == index ? 14'h880 : _GEN_13061;
  wire [13:0] _GEN_13063 = 14'h3307 == index ? 14'h704 : _GEN_13062;
  wire [13:0] _GEN_13064 = 14'h3308 == index ? 14'h606 : _GEN_13063;
  wire [13:0] _GEN_13065 = 14'h3309 == index ? 14'h583 : _GEN_13064;
  wire [13:0] _GEN_13066 = 14'h330a == index ? 14'h502 : _GEN_13065;
  wire [13:0] _GEN_13067 = 14'h330b == index ? 14'h483 : _GEN_13066;
  wire [13:0] _GEN_13068 = 14'h330c == index ? 14'h406 : _GEN_13067;
  wire [13:0] _GEN_13069 = 14'h330d == index ? 14'h38b : _GEN_13068;
  wire [13:0] _GEN_13070 = 14'h330e == index ? 14'h384 : _GEN_13069;
  wire [13:0] _GEN_13071 = 14'h330f == index ? 14'h30c : _GEN_13070;
  wire [13:0] _GEN_13072 = 14'h3310 == index ? 14'h306 : _GEN_13071;
  wire [13:0] _GEN_13073 = 14'h3311 == index ? 14'h300 : _GEN_13072;
  wire [13:0] _GEN_13074 = 14'h3312 == index ? 14'h28c : _GEN_13073;
  wire [13:0] _GEN_13075 = 14'h3313 == index ? 14'h287 : _GEN_13074;
  wire [13:0] _GEN_13076 = 14'h3314 == index ? 14'h282 : _GEN_13075;
  wire [13:0] _GEN_13077 = 14'h3315 == index ? 14'h212 : _GEN_13076;
  wire [13:0] _GEN_13078 = 14'h3316 == index ? 14'h20e : _GEN_13077;
  wire [13:0] _GEN_13079 = 14'h3317 == index ? 14'h20a : _GEN_13078;
  wire [13:0] _GEN_13080 = 14'h3318 == index ? 14'h206 : _GEN_13079;
  wire [13:0] _GEN_13081 = 14'h3319 == index ? 14'h202 : _GEN_13080;
  wire [13:0] _GEN_13082 = 14'h331a == index ? 14'h198 : _GEN_13081;
  wire [13:0] _GEN_13083 = 14'h331b == index ? 14'h195 : _GEN_13082;
  wire [13:0] _GEN_13084 = 14'h331c == index ? 14'h192 : _GEN_13083;
  wire [13:0] _GEN_13085 = 14'h331d == index ? 14'h18f : _GEN_13084;
  wire [13:0] _GEN_13086 = 14'h331e == index ? 14'h18c : _GEN_13085;
  wire [13:0] _GEN_13087 = 14'h331f == index ? 14'h189 : _GEN_13086;
  wire [13:0] _GEN_13088 = 14'h3320 == index ? 14'h186 : _GEN_13087;
  wire [13:0] _GEN_13089 = 14'h3321 == index ? 14'h183 : _GEN_13088;
  wire [13:0] _GEN_13090 = 14'h3322 == index ? 14'h180 : _GEN_13089;
  wire [13:0] _GEN_13091 = 14'h3323 == index ? 14'h120 : _GEN_13090;
  wire [13:0] _GEN_13092 = 14'h3324 == index ? 14'h11e : _GEN_13091;
  wire [13:0] _GEN_13093 = 14'h3325 == index ? 14'h11c : _GEN_13092;
  wire [13:0] _GEN_13094 = 14'h3326 == index ? 14'h11a : _GEN_13093;
  wire [13:0] _GEN_13095 = 14'h3327 == index ? 14'h118 : _GEN_13094;
  wire [13:0] _GEN_13096 = 14'h3328 == index ? 14'h116 : _GEN_13095;
  wire [13:0] _GEN_13097 = 14'h3329 == index ? 14'h114 : _GEN_13096;
  wire [13:0] _GEN_13098 = 14'h332a == index ? 14'h112 : _GEN_13097;
  wire [13:0] _GEN_13099 = 14'h332b == index ? 14'h110 : _GEN_13098;
  wire [13:0] _GEN_13100 = 14'h332c == index ? 14'h10e : _GEN_13099;
  wire [13:0] _GEN_13101 = 14'h332d == index ? 14'h10c : _GEN_13100;
  wire [13:0] _GEN_13102 = 14'h332e == index ? 14'h10a : _GEN_13101;
  wire [13:0] _GEN_13103 = 14'h332f == index ? 14'h108 : _GEN_13102;
  wire [13:0] _GEN_13104 = 14'h3330 == index ? 14'h106 : _GEN_13103;
  wire [13:0] _GEN_13105 = 14'h3331 == index ? 14'h104 : _GEN_13104;
  wire [13:0] _GEN_13106 = 14'h3332 == index ? 14'h102 : _GEN_13105;
  wire [13:0] _GEN_13107 = 14'h3333 == index ? 14'h100 : _GEN_13106;
  wire [13:0] _GEN_13108 = 14'h3334 == index ? 14'hb2 : _GEN_13107;
  wire [13:0] _GEN_13109 = 14'h3335 == index ? 14'hb1 : _GEN_13108;
  wire [13:0] _GEN_13110 = 14'h3336 == index ? 14'hb0 : _GEN_13109;
  wire [13:0] _GEN_13111 = 14'h3337 == index ? 14'haf : _GEN_13110;
  wire [13:0] _GEN_13112 = 14'h3338 == index ? 14'hae : _GEN_13111;
  wire [13:0] _GEN_13113 = 14'h3339 == index ? 14'had : _GEN_13112;
  wire [13:0] _GEN_13114 = 14'h333a == index ? 14'hac : _GEN_13113;
  wire [13:0] _GEN_13115 = 14'h333b == index ? 14'hab : _GEN_13114;
  wire [13:0] _GEN_13116 = 14'h333c == index ? 14'haa : _GEN_13115;
  wire [13:0] _GEN_13117 = 14'h333d == index ? 14'ha9 : _GEN_13116;
  wire [13:0] _GEN_13118 = 14'h333e == index ? 14'ha8 : _GEN_13117;
  wire [13:0] _GEN_13119 = 14'h333f == index ? 14'ha7 : _GEN_13118;
  wire [13:0] _GEN_13120 = 14'h3340 == index ? 14'ha6 : _GEN_13119;
  wire [13:0] _GEN_13121 = 14'h3341 == index ? 14'ha5 : _GEN_13120;
  wire [13:0] _GEN_13122 = 14'h3342 == index ? 14'ha4 : _GEN_13121;
  wire [13:0] _GEN_13123 = 14'h3343 == index ? 14'ha3 : _GEN_13122;
  wire [13:0] _GEN_13124 = 14'h3344 == index ? 14'ha2 : _GEN_13123;
  wire [13:0] _GEN_13125 = 14'h3345 == index ? 14'ha1 : _GEN_13124;
  wire [13:0] _GEN_13126 = 14'h3346 == index ? 14'ha0 : _GEN_13125;
  wire [13:0] _GEN_13127 = 14'h3347 == index ? 14'h9f : _GEN_13126;
  wire [13:0] _GEN_13128 = 14'h3348 == index ? 14'h9e : _GEN_13127;
  wire [13:0] _GEN_13129 = 14'h3349 == index ? 14'h9d : _GEN_13128;
  wire [13:0] _GEN_13130 = 14'h334a == index ? 14'h9c : _GEN_13129;
  wire [13:0] _GEN_13131 = 14'h334b == index ? 14'h9b : _GEN_13130;
  wire [13:0] _GEN_13132 = 14'h334c == index ? 14'h9a : _GEN_13131;
  wire [13:0] _GEN_13133 = 14'h334d == index ? 14'h99 : _GEN_13132;
  wire [13:0] _GEN_13134 = 14'h334e == index ? 14'h98 : _GEN_13133;
  wire [13:0] _GEN_13135 = 14'h334f == index ? 14'h97 : _GEN_13134;
  wire [13:0] _GEN_13136 = 14'h3350 == index ? 14'h96 : _GEN_13135;
  wire [13:0] _GEN_13137 = 14'h3351 == index ? 14'h95 : _GEN_13136;
  wire [13:0] _GEN_13138 = 14'h3352 == index ? 14'h94 : _GEN_13137;
  wire [13:0] _GEN_13139 = 14'h3353 == index ? 14'h93 : _GEN_13138;
  wire [13:0] _GEN_13140 = 14'h3354 == index ? 14'h92 : _GEN_13139;
  wire [13:0] _GEN_13141 = 14'h3355 == index ? 14'h91 : _GEN_13140;
  wire [13:0] _GEN_13142 = 14'h3356 == index ? 14'h90 : _GEN_13141;
  wire [13:0] _GEN_13143 = 14'h3357 == index ? 14'h8f : _GEN_13142;
  wire [13:0] _GEN_13144 = 14'h3358 == index ? 14'h8e : _GEN_13143;
  wire [13:0] _GEN_13145 = 14'h3359 == index ? 14'h8d : _GEN_13144;
  wire [13:0] _GEN_13146 = 14'h335a == index ? 14'h8c : _GEN_13145;
  wire [13:0] _GEN_13147 = 14'h335b == index ? 14'h8b : _GEN_13146;
  wire [13:0] _GEN_13148 = 14'h335c == index ? 14'h8a : _GEN_13147;
  wire [13:0] _GEN_13149 = 14'h335d == index ? 14'h89 : _GEN_13148;
  wire [13:0] _GEN_13150 = 14'h335e == index ? 14'h88 : _GEN_13149;
  wire [13:0] _GEN_13151 = 14'h335f == index ? 14'h87 : _GEN_13150;
  wire [13:0] _GEN_13152 = 14'h3360 == index ? 14'h86 : _GEN_13151;
  wire [13:0] _GEN_13153 = 14'h3361 == index ? 14'h85 : _GEN_13152;
  wire [13:0] _GEN_13154 = 14'h3362 == index ? 14'h84 : _GEN_13153;
  wire [13:0] _GEN_13155 = 14'h3363 == index ? 14'h83 : _GEN_13154;
  wire [13:0] _GEN_13156 = 14'h3364 == index ? 14'h82 : _GEN_13155;
  wire [13:0] _GEN_13157 = 14'h3365 == index ? 14'h81 : _GEN_13156;
  wire [13:0] _GEN_13158 = 14'h3366 == index ? 14'h80 : _GEN_13157;
  wire [13:0] _GEN_13159 = 14'h3367 == index ? 14'h66 : _GEN_13158;
  wire [13:0] _GEN_13160 = 14'h3368 == index ? 14'h66 : _GEN_13159;
  wire [13:0] _GEN_13161 = 14'h3369 == index ? 14'h66 : _GEN_13160;
  wire [13:0] _GEN_13162 = 14'h336a == index ? 14'h66 : _GEN_13161;
  wire [13:0] _GEN_13163 = 14'h336b == index ? 14'h66 : _GEN_13162;
  wire [13:0] _GEN_13164 = 14'h336c == index ? 14'h66 : _GEN_13163;
  wire [13:0] _GEN_13165 = 14'h336d == index ? 14'h66 : _GEN_13164;
  wire [13:0] _GEN_13166 = 14'h336e == index ? 14'h66 : _GEN_13165;
  wire [13:0] _GEN_13167 = 14'h336f == index ? 14'h66 : _GEN_13166;
  wire [13:0] _GEN_13168 = 14'h3370 == index ? 14'h66 : _GEN_13167;
  wire [13:0] _GEN_13169 = 14'h3371 == index ? 14'h66 : _GEN_13168;
  wire [13:0] _GEN_13170 = 14'h3372 == index ? 14'h66 : _GEN_13169;
  wire [13:0] _GEN_13171 = 14'h3373 == index ? 14'h66 : _GEN_13170;
  wire [13:0] _GEN_13172 = 14'h3374 == index ? 14'h66 : _GEN_13171;
  wire [13:0] _GEN_13173 = 14'h3375 == index ? 14'h66 : _GEN_13172;
  wire [13:0] _GEN_13174 = 14'h3376 == index ? 14'h66 : _GEN_13173;
  wire [13:0] _GEN_13175 = 14'h3377 == index ? 14'h66 : _GEN_13174;
  wire [13:0] _GEN_13176 = 14'h3378 == index ? 14'h66 : _GEN_13175;
  wire [13:0] _GEN_13177 = 14'h3379 == index ? 14'h66 : _GEN_13176;
  wire [13:0] _GEN_13178 = 14'h337a == index ? 14'h66 : _GEN_13177;
  wire [13:0] _GEN_13179 = 14'h337b == index ? 14'h66 : _GEN_13178;
  wire [13:0] _GEN_13180 = 14'h337c == index ? 14'h66 : _GEN_13179;
  wire [13:0] _GEN_13181 = 14'h337d == index ? 14'h66 : _GEN_13180;
  wire [13:0] _GEN_13182 = 14'h337e == index ? 14'h66 : _GEN_13181;
  wire [13:0] _GEN_13183 = 14'h337f == index ? 14'h66 : _GEN_13182;
  wire [13:0] _GEN_13184 = 14'h3380 == index ? 14'h0 : _GEN_13183;
  wire [13:0] _GEN_13185 = 14'h3381 == index ? 14'h3380 : _GEN_13184;
  wire [13:0] _GEN_13186 = 14'h3382 == index ? 14'h1981 : _GEN_13185;
  wire [13:0] _GEN_13187 = 14'h3383 == index ? 14'h1101 : _GEN_13186;
  wire [13:0] _GEN_13188 = 14'h3384 == index ? 14'hc83 : _GEN_13187;
  wire [13:0] _GEN_13189 = 14'h3385 == index ? 14'ha03 : _GEN_13188;
  wire [13:0] _GEN_13190 = 14'h3386 == index ? 14'h881 : _GEN_13189;
  wire [13:0] _GEN_13191 = 14'h3387 == index ? 14'h705 : _GEN_13190;
  wire [13:0] _GEN_13192 = 14'h3388 == index ? 14'h607 : _GEN_13191;
  wire [13:0] _GEN_13193 = 14'h3389 == index ? 14'h584 : _GEN_13192;
  wire [13:0] _GEN_13194 = 14'h338a == index ? 14'h503 : _GEN_13193;
  wire [13:0] _GEN_13195 = 14'h338b == index ? 14'h484 : _GEN_13194;
  wire [13:0] _GEN_13196 = 14'h338c == index ? 14'h407 : _GEN_13195;
  wire [13:0] _GEN_13197 = 14'h338d == index ? 14'h38c : _GEN_13196;
  wire [13:0] _GEN_13198 = 14'h338e == index ? 14'h385 : _GEN_13197;
  wire [13:0] _GEN_13199 = 14'h338f == index ? 14'h30d : _GEN_13198;
  wire [13:0] _GEN_13200 = 14'h3390 == index ? 14'h307 : _GEN_13199;
  wire [13:0] _GEN_13201 = 14'h3391 == index ? 14'h301 : _GEN_13200;
  wire [13:0] _GEN_13202 = 14'h3392 == index ? 14'h28d : _GEN_13201;
  wire [13:0] _GEN_13203 = 14'h3393 == index ? 14'h288 : _GEN_13202;
  wire [13:0] _GEN_13204 = 14'h3394 == index ? 14'h283 : _GEN_13203;
  wire [13:0] _GEN_13205 = 14'h3395 == index ? 14'h213 : _GEN_13204;
  wire [13:0] _GEN_13206 = 14'h3396 == index ? 14'h20f : _GEN_13205;
  wire [13:0] _GEN_13207 = 14'h3397 == index ? 14'h20b : _GEN_13206;
  wire [13:0] _GEN_13208 = 14'h3398 == index ? 14'h207 : _GEN_13207;
  wire [13:0] _GEN_13209 = 14'h3399 == index ? 14'h203 : _GEN_13208;
  wire [13:0] _GEN_13210 = 14'h339a == index ? 14'h199 : _GEN_13209;
  wire [13:0] _GEN_13211 = 14'h339b == index ? 14'h196 : _GEN_13210;
  wire [13:0] _GEN_13212 = 14'h339c == index ? 14'h193 : _GEN_13211;
  wire [13:0] _GEN_13213 = 14'h339d == index ? 14'h190 : _GEN_13212;
  wire [13:0] _GEN_13214 = 14'h339e == index ? 14'h18d : _GEN_13213;
  wire [13:0] _GEN_13215 = 14'h339f == index ? 14'h18a : _GEN_13214;
  wire [13:0] _GEN_13216 = 14'h33a0 == index ? 14'h187 : _GEN_13215;
  wire [13:0] _GEN_13217 = 14'h33a1 == index ? 14'h184 : _GEN_13216;
  wire [13:0] _GEN_13218 = 14'h33a2 == index ? 14'h181 : _GEN_13217;
  wire [13:0] _GEN_13219 = 14'h33a3 == index ? 14'h121 : _GEN_13218;
  wire [13:0] _GEN_13220 = 14'h33a4 == index ? 14'h11f : _GEN_13219;
  wire [13:0] _GEN_13221 = 14'h33a5 == index ? 14'h11d : _GEN_13220;
  wire [13:0] _GEN_13222 = 14'h33a6 == index ? 14'h11b : _GEN_13221;
  wire [13:0] _GEN_13223 = 14'h33a7 == index ? 14'h119 : _GEN_13222;
  wire [13:0] _GEN_13224 = 14'h33a8 == index ? 14'h117 : _GEN_13223;
  wire [13:0] _GEN_13225 = 14'h33a9 == index ? 14'h115 : _GEN_13224;
  wire [13:0] _GEN_13226 = 14'h33aa == index ? 14'h113 : _GEN_13225;
  wire [13:0] _GEN_13227 = 14'h33ab == index ? 14'h111 : _GEN_13226;
  wire [13:0] _GEN_13228 = 14'h33ac == index ? 14'h10f : _GEN_13227;
  wire [13:0] _GEN_13229 = 14'h33ad == index ? 14'h10d : _GEN_13228;
  wire [13:0] _GEN_13230 = 14'h33ae == index ? 14'h10b : _GEN_13229;
  wire [13:0] _GEN_13231 = 14'h33af == index ? 14'h109 : _GEN_13230;
  wire [13:0] _GEN_13232 = 14'h33b0 == index ? 14'h107 : _GEN_13231;
  wire [13:0] _GEN_13233 = 14'h33b1 == index ? 14'h105 : _GEN_13232;
  wire [13:0] _GEN_13234 = 14'h33b2 == index ? 14'h103 : _GEN_13233;
  wire [13:0] _GEN_13235 = 14'h33b3 == index ? 14'h101 : _GEN_13234;
  wire [13:0] _GEN_13236 = 14'h33b4 == index ? 14'hb3 : _GEN_13235;
  wire [13:0] _GEN_13237 = 14'h33b5 == index ? 14'hb2 : _GEN_13236;
  wire [13:0] _GEN_13238 = 14'h33b6 == index ? 14'hb1 : _GEN_13237;
  wire [13:0] _GEN_13239 = 14'h33b7 == index ? 14'hb0 : _GEN_13238;
  wire [13:0] _GEN_13240 = 14'h33b8 == index ? 14'haf : _GEN_13239;
  wire [13:0] _GEN_13241 = 14'h33b9 == index ? 14'hae : _GEN_13240;
  wire [13:0] _GEN_13242 = 14'h33ba == index ? 14'had : _GEN_13241;
  wire [13:0] _GEN_13243 = 14'h33bb == index ? 14'hac : _GEN_13242;
  wire [13:0] _GEN_13244 = 14'h33bc == index ? 14'hab : _GEN_13243;
  wire [13:0] _GEN_13245 = 14'h33bd == index ? 14'haa : _GEN_13244;
  wire [13:0] _GEN_13246 = 14'h33be == index ? 14'ha9 : _GEN_13245;
  wire [13:0] _GEN_13247 = 14'h33bf == index ? 14'ha8 : _GEN_13246;
  wire [13:0] _GEN_13248 = 14'h33c0 == index ? 14'ha7 : _GEN_13247;
  wire [13:0] _GEN_13249 = 14'h33c1 == index ? 14'ha6 : _GEN_13248;
  wire [13:0] _GEN_13250 = 14'h33c2 == index ? 14'ha5 : _GEN_13249;
  wire [13:0] _GEN_13251 = 14'h33c3 == index ? 14'ha4 : _GEN_13250;
  wire [13:0] _GEN_13252 = 14'h33c4 == index ? 14'ha3 : _GEN_13251;
  wire [13:0] _GEN_13253 = 14'h33c5 == index ? 14'ha2 : _GEN_13252;
  wire [13:0] _GEN_13254 = 14'h33c6 == index ? 14'ha1 : _GEN_13253;
  wire [13:0] _GEN_13255 = 14'h33c7 == index ? 14'ha0 : _GEN_13254;
  wire [13:0] _GEN_13256 = 14'h33c8 == index ? 14'h9f : _GEN_13255;
  wire [13:0] _GEN_13257 = 14'h33c9 == index ? 14'h9e : _GEN_13256;
  wire [13:0] _GEN_13258 = 14'h33ca == index ? 14'h9d : _GEN_13257;
  wire [13:0] _GEN_13259 = 14'h33cb == index ? 14'h9c : _GEN_13258;
  wire [13:0] _GEN_13260 = 14'h33cc == index ? 14'h9b : _GEN_13259;
  wire [13:0] _GEN_13261 = 14'h33cd == index ? 14'h9a : _GEN_13260;
  wire [13:0] _GEN_13262 = 14'h33ce == index ? 14'h99 : _GEN_13261;
  wire [13:0] _GEN_13263 = 14'h33cf == index ? 14'h98 : _GEN_13262;
  wire [13:0] _GEN_13264 = 14'h33d0 == index ? 14'h97 : _GEN_13263;
  wire [13:0] _GEN_13265 = 14'h33d1 == index ? 14'h96 : _GEN_13264;
  wire [13:0] _GEN_13266 = 14'h33d2 == index ? 14'h95 : _GEN_13265;
  wire [13:0] _GEN_13267 = 14'h33d3 == index ? 14'h94 : _GEN_13266;
  wire [13:0] _GEN_13268 = 14'h33d4 == index ? 14'h93 : _GEN_13267;
  wire [13:0] _GEN_13269 = 14'h33d5 == index ? 14'h92 : _GEN_13268;
  wire [13:0] _GEN_13270 = 14'h33d6 == index ? 14'h91 : _GEN_13269;
  wire [13:0] _GEN_13271 = 14'h33d7 == index ? 14'h90 : _GEN_13270;
  wire [13:0] _GEN_13272 = 14'h33d8 == index ? 14'h8f : _GEN_13271;
  wire [13:0] _GEN_13273 = 14'h33d9 == index ? 14'h8e : _GEN_13272;
  wire [13:0] _GEN_13274 = 14'h33da == index ? 14'h8d : _GEN_13273;
  wire [13:0] _GEN_13275 = 14'h33db == index ? 14'h8c : _GEN_13274;
  wire [13:0] _GEN_13276 = 14'h33dc == index ? 14'h8b : _GEN_13275;
  wire [13:0] _GEN_13277 = 14'h33dd == index ? 14'h8a : _GEN_13276;
  wire [13:0] _GEN_13278 = 14'h33de == index ? 14'h89 : _GEN_13277;
  wire [13:0] _GEN_13279 = 14'h33df == index ? 14'h88 : _GEN_13278;
  wire [13:0] _GEN_13280 = 14'h33e0 == index ? 14'h87 : _GEN_13279;
  wire [13:0] _GEN_13281 = 14'h33e1 == index ? 14'h86 : _GEN_13280;
  wire [13:0] _GEN_13282 = 14'h33e2 == index ? 14'h85 : _GEN_13281;
  wire [13:0] _GEN_13283 = 14'h33e3 == index ? 14'h84 : _GEN_13282;
  wire [13:0] _GEN_13284 = 14'h33e4 == index ? 14'h83 : _GEN_13283;
  wire [13:0] _GEN_13285 = 14'h33e5 == index ? 14'h82 : _GEN_13284;
  wire [13:0] _GEN_13286 = 14'h33e6 == index ? 14'h81 : _GEN_13285;
  wire [13:0] _GEN_13287 = 14'h33e7 == index ? 14'h80 : _GEN_13286;
  wire [13:0] _GEN_13288 = 14'h33e8 == index ? 14'h67 : _GEN_13287;
  wire [13:0] _GEN_13289 = 14'h33e9 == index ? 14'h67 : _GEN_13288;
  wire [13:0] _GEN_13290 = 14'h33ea == index ? 14'h67 : _GEN_13289;
  wire [13:0] _GEN_13291 = 14'h33eb == index ? 14'h67 : _GEN_13290;
  wire [13:0] _GEN_13292 = 14'h33ec == index ? 14'h67 : _GEN_13291;
  wire [13:0] _GEN_13293 = 14'h33ed == index ? 14'h67 : _GEN_13292;
  wire [13:0] _GEN_13294 = 14'h33ee == index ? 14'h67 : _GEN_13293;
  wire [13:0] _GEN_13295 = 14'h33ef == index ? 14'h67 : _GEN_13294;
  wire [13:0] _GEN_13296 = 14'h33f0 == index ? 14'h67 : _GEN_13295;
  wire [13:0] _GEN_13297 = 14'h33f1 == index ? 14'h67 : _GEN_13296;
  wire [13:0] _GEN_13298 = 14'h33f2 == index ? 14'h67 : _GEN_13297;
  wire [13:0] _GEN_13299 = 14'h33f3 == index ? 14'h67 : _GEN_13298;
  wire [13:0] _GEN_13300 = 14'h33f4 == index ? 14'h67 : _GEN_13299;
  wire [13:0] _GEN_13301 = 14'h33f5 == index ? 14'h67 : _GEN_13300;
  wire [13:0] _GEN_13302 = 14'h33f6 == index ? 14'h67 : _GEN_13301;
  wire [13:0] _GEN_13303 = 14'h33f7 == index ? 14'h67 : _GEN_13302;
  wire [13:0] _GEN_13304 = 14'h33f8 == index ? 14'h67 : _GEN_13303;
  wire [13:0] _GEN_13305 = 14'h33f9 == index ? 14'h67 : _GEN_13304;
  wire [13:0] _GEN_13306 = 14'h33fa == index ? 14'h67 : _GEN_13305;
  wire [13:0] _GEN_13307 = 14'h33fb == index ? 14'h67 : _GEN_13306;
  wire [13:0] _GEN_13308 = 14'h33fc == index ? 14'h67 : _GEN_13307;
  wire [13:0] _GEN_13309 = 14'h33fd == index ? 14'h67 : _GEN_13308;
  wire [13:0] _GEN_13310 = 14'h33fe == index ? 14'h67 : _GEN_13309;
  wire [13:0] _GEN_13311 = 14'h33ff == index ? 14'h67 : _GEN_13310;
  wire [13:0] _GEN_13312 = 14'h3400 == index ? 14'h0 : _GEN_13311;
  wire [13:0] _GEN_13313 = 14'h3401 == index ? 14'h3400 : _GEN_13312;
  wire [13:0] _GEN_13314 = 14'h3402 == index ? 14'h1a00 : _GEN_13313;
  wire [13:0] _GEN_13315 = 14'h3403 == index ? 14'h1102 : _GEN_13314;
  wire [13:0] _GEN_13316 = 14'h3404 == index ? 14'hd00 : _GEN_13315;
  wire [13:0] _GEN_13317 = 14'h3405 == index ? 14'ha04 : _GEN_13316;
  wire [13:0] _GEN_13318 = 14'h3406 == index ? 14'h882 : _GEN_13317;
  wire [13:0] _GEN_13319 = 14'h3407 == index ? 14'h706 : _GEN_13318;
  wire [13:0] _GEN_13320 = 14'h3408 == index ? 14'h680 : _GEN_13319;
  wire [13:0] _GEN_13321 = 14'h3409 == index ? 14'h585 : _GEN_13320;
  wire [13:0] _GEN_13322 = 14'h340a == index ? 14'h504 : _GEN_13321;
  wire [13:0] _GEN_13323 = 14'h340b == index ? 14'h485 : _GEN_13322;
  wire [13:0] _GEN_13324 = 14'h340c == index ? 14'h408 : _GEN_13323;
  wire [13:0] _GEN_13325 = 14'h340d == index ? 14'h400 : _GEN_13324;
  wire [13:0] _GEN_13326 = 14'h340e == index ? 14'h386 : _GEN_13325;
  wire [13:0] _GEN_13327 = 14'h340f == index ? 14'h30e : _GEN_13326;
  wire [13:0] _GEN_13328 = 14'h3410 == index ? 14'h308 : _GEN_13327;
  wire [13:0] _GEN_13329 = 14'h3411 == index ? 14'h302 : _GEN_13328;
  wire [13:0] _GEN_13330 = 14'h3412 == index ? 14'h28e : _GEN_13329;
  wire [13:0] _GEN_13331 = 14'h3413 == index ? 14'h289 : _GEN_13330;
  wire [13:0] _GEN_13332 = 14'h3414 == index ? 14'h284 : _GEN_13331;
  wire [13:0] _GEN_13333 = 14'h3415 == index ? 14'h214 : _GEN_13332;
  wire [13:0] _GEN_13334 = 14'h3416 == index ? 14'h210 : _GEN_13333;
  wire [13:0] _GEN_13335 = 14'h3417 == index ? 14'h20c : _GEN_13334;
  wire [13:0] _GEN_13336 = 14'h3418 == index ? 14'h208 : _GEN_13335;
  wire [13:0] _GEN_13337 = 14'h3419 == index ? 14'h204 : _GEN_13336;
  wire [13:0] _GEN_13338 = 14'h341a == index ? 14'h200 : _GEN_13337;
  wire [13:0] _GEN_13339 = 14'h341b == index ? 14'h197 : _GEN_13338;
  wire [13:0] _GEN_13340 = 14'h341c == index ? 14'h194 : _GEN_13339;
  wire [13:0] _GEN_13341 = 14'h341d == index ? 14'h191 : _GEN_13340;
  wire [13:0] _GEN_13342 = 14'h341e == index ? 14'h18e : _GEN_13341;
  wire [13:0] _GEN_13343 = 14'h341f == index ? 14'h18b : _GEN_13342;
  wire [13:0] _GEN_13344 = 14'h3420 == index ? 14'h188 : _GEN_13343;
  wire [13:0] _GEN_13345 = 14'h3421 == index ? 14'h185 : _GEN_13344;
  wire [13:0] _GEN_13346 = 14'h3422 == index ? 14'h182 : _GEN_13345;
  wire [13:0] _GEN_13347 = 14'h3423 == index ? 14'h122 : _GEN_13346;
  wire [13:0] _GEN_13348 = 14'h3424 == index ? 14'h120 : _GEN_13347;
  wire [13:0] _GEN_13349 = 14'h3425 == index ? 14'h11e : _GEN_13348;
  wire [13:0] _GEN_13350 = 14'h3426 == index ? 14'h11c : _GEN_13349;
  wire [13:0] _GEN_13351 = 14'h3427 == index ? 14'h11a : _GEN_13350;
  wire [13:0] _GEN_13352 = 14'h3428 == index ? 14'h118 : _GEN_13351;
  wire [13:0] _GEN_13353 = 14'h3429 == index ? 14'h116 : _GEN_13352;
  wire [13:0] _GEN_13354 = 14'h342a == index ? 14'h114 : _GEN_13353;
  wire [13:0] _GEN_13355 = 14'h342b == index ? 14'h112 : _GEN_13354;
  wire [13:0] _GEN_13356 = 14'h342c == index ? 14'h110 : _GEN_13355;
  wire [13:0] _GEN_13357 = 14'h342d == index ? 14'h10e : _GEN_13356;
  wire [13:0] _GEN_13358 = 14'h342e == index ? 14'h10c : _GEN_13357;
  wire [13:0] _GEN_13359 = 14'h342f == index ? 14'h10a : _GEN_13358;
  wire [13:0] _GEN_13360 = 14'h3430 == index ? 14'h108 : _GEN_13359;
  wire [13:0] _GEN_13361 = 14'h3431 == index ? 14'h106 : _GEN_13360;
  wire [13:0] _GEN_13362 = 14'h3432 == index ? 14'h104 : _GEN_13361;
  wire [13:0] _GEN_13363 = 14'h3433 == index ? 14'h102 : _GEN_13362;
  wire [13:0] _GEN_13364 = 14'h3434 == index ? 14'h100 : _GEN_13363;
  wire [13:0] _GEN_13365 = 14'h3435 == index ? 14'hb3 : _GEN_13364;
  wire [13:0] _GEN_13366 = 14'h3436 == index ? 14'hb2 : _GEN_13365;
  wire [13:0] _GEN_13367 = 14'h3437 == index ? 14'hb1 : _GEN_13366;
  wire [13:0] _GEN_13368 = 14'h3438 == index ? 14'hb0 : _GEN_13367;
  wire [13:0] _GEN_13369 = 14'h3439 == index ? 14'haf : _GEN_13368;
  wire [13:0] _GEN_13370 = 14'h343a == index ? 14'hae : _GEN_13369;
  wire [13:0] _GEN_13371 = 14'h343b == index ? 14'had : _GEN_13370;
  wire [13:0] _GEN_13372 = 14'h343c == index ? 14'hac : _GEN_13371;
  wire [13:0] _GEN_13373 = 14'h343d == index ? 14'hab : _GEN_13372;
  wire [13:0] _GEN_13374 = 14'h343e == index ? 14'haa : _GEN_13373;
  wire [13:0] _GEN_13375 = 14'h343f == index ? 14'ha9 : _GEN_13374;
  wire [13:0] _GEN_13376 = 14'h3440 == index ? 14'ha8 : _GEN_13375;
  wire [13:0] _GEN_13377 = 14'h3441 == index ? 14'ha7 : _GEN_13376;
  wire [13:0] _GEN_13378 = 14'h3442 == index ? 14'ha6 : _GEN_13377;
  wire [13:0] _GEN_13379 = 14'h3443 == index ? 14'ha5 : _GEN_13378;
  wire [13:0] _GEN_13380 = 14'h3444 == index ? 14'ha4 : _GEN_13379;
  wire [13:0] _GEN_13381 = 14'h3445 == index ? 14'ha3 : _GEN_13380;
  wire [13:0] _GEN_13382 = 14'h3446 == index ? 14'ha2 : _GEN_13381;
  wire [13:0] _GEN_13383 = 14'h3447 == index ? 14'ha1 : _GEN_13382;
  wire [13:0] _GEN_13384 = 14'h3448 == index ? 14'ha0 : _GEN_13383;
  wire [13:0] _GEN_13385 = 14'h3449 == index ? 14'h9f : _GEN_13384;
  wire [13:0] _GEN_13386 = 14'h344a == index ? 14'h9e : _GEN_13385;
  wire [13:0] _GEN_13387 = 14'h344b == index ? 14'h9d : _GEN_13386;
  wire [13:0] _GEN_13388 = 14'h344c == index ? 14'h9c : _GEN_13387;
  wire [13:0] _GEN_13389 = 14'h344d == index ? 14'h9b : _GEN_13388;
  wire [13:0] _GEN_13390 = 14'h344e == index ? 14'h9a : _GEN_13389;
  wire [13:0] _GEN_13391 = 14'h344f == index ? 14'h99 : _GEN_13390;
  wire [13:0] _GEN_13392 = 14'h3450 == index ? 14'h98 : _GEN_13391;
  wire [13:0] _GEN_13393 = 14'h3451 == index ? 14'h97 : _GEN_13392;
  wire [13:0] _GEN_13394 = 14'h3452 == index ? 14'h96 : _GEN_13393;
  wire [13:0] _GEN_13395 = 14'h3453 == index ? 14'h95 : _GEN_13394;
  wire [13:0] _GEN_13396 = 14'h3454 == index ? 14'h94 : _GEN_13395;
  wire [13:0] _GEN_13397 = 14'h3455 == index ? 14'h93 : _GEN_13396;
  wire [13:0] _GEN_13398 = 14'h3456 == index ? 14'h92 : _GEN_13397;
  wire [13:0] _GEN_13399 = 14'h3457 == index ? 14'h91 : _GEN_13398;
  wire [13:0] _GEN_13400 = 14'h3458 == index ? 14'h90 : _GEN_13399;
  wire [13:0] _GEN_13401 = 14'h3459 == index ? 14'h8f : _GEN_13400;
  wire [13:0] _GEN_13402 = 14'h345a == index ? 14'h8e : _GEN_13401;
  wire [13:0] _GEN_13403 = 14'h345b == index ? 14'h8d : _GEN_13402;
  wire [13:0] _GEN_13404 = 14'h345c == index ? 14'h8c : _GEN_13403;
  wire [13:0] _GEN_13405 = 14'h345d == index ? 14'h8b : _GEN_13404;
  wire [13:0] _GEN_13406 = 14'h345e == index ? 14'h8a : _GEN_13405;
  wire [13:0] _GEN_13407 = 14'h345f == index ? 14'h89 : _GEN_13406;
  wire [13:0] _GEN_13408 = 14'h3460 == index ? 14'h88 : _GEN_13407;
  wire [13:0] _GEN_13409 = 14'h3461 == index ? 14'h87 : _GEN_13408;
  wire [13:0] _GEN_13410 = 14'h3462 == index ? 14'h86 : _GEN_13409;
  wire [13:0] _GEN_13411 = 14'h3463 == index ? 14'h85 : _GEN_13410;
  wire [13:0] _GEN_13412 = 14'h3464 == index ? 14'h84 : _GEN_13411;
  wire [13:0] _GEN_13413 = 14'h3465 == index ? 14'h83 : _GEN_13412;
  wire [13:0] _GEN_13414 = 14'h3466 == index ? 14'h82 : _GEN_13413;
  wire [13:0] _GEN_13415 = 14'h3467 == index ? 14'h81 : _GEN_13414;
  wire [13:0] _GEN_13416 = 14'h3468 == index ? 14'h80 : _GEN_13415;
  wire [13:0] _GEN_13417 = 14'h3469 == index ? 14'h68 : _GEN_13416;
  wire [13:0] _GEN_13418 = 14'h346a == index ? 14'h68 : _GEN_13417;
  wire [13:0] _GEN_13419 = 14'h346b == index ? 14'h68 : _GEN_13418;
  wire [13:0] _GEN_13420 = 14'h346c == index ? 14'h68 : _GEN_13419;
  wire [13:0] _GEN_13421 = 14'h346d == index ? 14'h68 : _GEN_13420;
  wire [13:0] _GEN_13422 = 14'h346e == index ? 14'h68 : _GEN_13421;
  wire [13:0] _GEN_13423 = 14'h346f == index ? 14'h68 : _GEN_13422;
  wire [13:0] _GEN_13424 = 14'h3470 == index ? 14'h68 : _GEN_13423;
  wire [13:0] _GEN_13425 = 14'h3471 == index ? 14'h68 : _GEN_13424;
  wire [13:0] _GEN_13426 = 14'h3472 == index ? 14'h68 : _GEN_13425;
  wire [13:0] _GEN_13427 = 14'h3473 == index ? 14'h68 : _GEN_13426;
  wire [13:0] _GEN_13428 = 14'h3474 == index ? 14'h68 : _GEN_13427;
  wire [13:0] _GEN_13429 = 14'h3475 == index ? 14'h68 : _GEN_13428;
  wire [13:0] _GEN_13430 = 14'h3476 == index ? 14'h68 : _GEN_13429;
  wire [13:0] _GEN_13431 = 14'h3477 == index ? 14'h68 : _GEN_13430;
  wire [13:0] _GEN_13432 = 14'h3478 == index ? 14'h68 : _GEN_13431;
  wire [13:0] _GEN_13433 = 14'h3479 == index ? 14'h68 : _GEN_13432;
  wire [13:0] _GEN_13434 = 14'h347a == index ? 14'h68 : _GEN_13433;
  wire [13:0] _GEN_13435 = 14'h347b == index ? 14'h68 : _GEN_13434;
  wire [13:0] _GEN_13436 = 14'h347c == index ? 14'h68 : _GEN_13435;
  wire [13:0] _GEN_13437 = 14'h347d == index ? 14'h68 : _GEN_13436;
  wire [13:0] _GEN_13438 = 14'h347e == index ? 14'h68 : _GEN_13437;
  wire [13:0] _GEN_13439 = 14'h347f == index ? 14'h68 : _GEN_13438;
  wire [13:0] _GEN_13440 = 14'h3480 == index ? 14'h0 : _GEN_13439;
  wire [13:0] _GEN_13441 = 14'h3481 == index ? 14'h3480 : _GEN_13440;
  wire [13:0] _GEN_13442 = 14'h3482 == index ? 14'h1a01 : _GEN_13441;
  wire [13:0] _GEN_13443 = 14'h3483 == index ? 14'h1180 : _GEN_13442;
  wire [13:0] _GEN_13444 = 14'h3484 == index ? 14'hd01 : _GEN_13443;
  wire [13:0] _GEN_13445 = 14'h3485 == index ? 14'ha80 : _GEN_13444;
  wire [13:0] _GEN_13446 = 14'h3486 == index ? 14'h883 : _GEN_13445;
  wire [13:0] _GEN_13447 = 14'h3487 == index ? 14'h780 : _GEN_13446;
  wire [13:0] _GEN_13448 = 14'h3488 == index ? 14'h681 : _GEN_13447;
  wire [13:0] _GEN_13449 = 14'h3489 == index ? 14'h586 : _GEN_13448;
  wire [13:0] _GEN_13450 = 14'h348a == index ? 14'h505 : _GEN_13449;
  wire [13:0] _GEN_13451 = 14'h348b == index ? 14'h486 : _GEN_13450;
  wire [13:0] _GEN_13452 = 14'h348c == index ? 14'h409 : _GEN_13451;
  wire [13:0] _GEN_13453 = 14'h348d == index ? 14'h401 : _GEN_13452;
  wire [13:0] _GEN_13454 = 14'h348e == index ? 14'h387 : _GEN_13453;
  wire [13:0] _GEN_13455 = 14'h348f == index ? 14'h380 : _GEN_13454;
  wire [13:0] _GEN_13456 = 14'h3490 == index ? 14'h309 : _GEN_13455;
  wire [13:0] _GEN_13457 = 14'h3491 == index ? 14'h303 : _GEN_13456;
  wire [13:0] _GEN_13458 = 14'h3492 == index ? 14'h28f : _GEN_13457;
  wire [13:0] _GEN_13459 = 14'h3493 == index ? 14'h28a : _GEN_13458;
  wire [13:0] _GEN_13460 = 14'h3494 == index ? 14'h285 : _GEN_13459;
  wire [13:0] _GEN_13461 = 14'h3495 == index ? 14'h280 : _GEN_13460;
  wire [13:0] _GEN_13462 = 14'h3496 == index ? 14'h211 : _GEN_13461;
  wire [13:0] _GEN_13463 = 14'h3497 == index ? 14'h20d : _GEN_13462;
  wire [13:0] _GEN_13464 = 14'h3498 == index ? 14'h209 : _GEN_13463;
  wire [13:0] _GEN_13465 = 14'h3499 == index ? 14'h205 : _GEN_13464;
  wire [13:0] _GEN_13466 = 14'h349a == index ? 14'h201 : _GEN_13465;
  wire [13:0] _GEN_13467 = 14'h349b == index ? 14'h198 : _GEN_13466;
  wire [13:0] _GEN_13468 = 14'h349c == index ? 14'h195 : _GEN_13467;
  wire [13:0] _GEN_13469 = 14'h349d == index ? 14'h192 : _GEN_13468;
  wire [13:0] _GEN_13470 = 14'h349e == index ? 14'h18f : _GEN_13469;
  wire [13:0] _GEN_13471 = 14'h349f == index ? 14'h18c : _GEN_13470;
  wire [13:0] _GEN_13472 = 14'h34a0 == index ? 14'h189 : _GEN_13471;
  wire [13:0] _GEN_13473 = 14'h34a1 == index ? 14'h186 : _GEN_13472;
  wire [13:0] _GEN_13474 = 14'h34a2 == index ? 14'h183 : _GEN_13473;
  wire [13:0] _GEN_13475 = 14'h34a3 == index ? 14'h180 : _GEN_13474;
  wire [13:0] _GEN_13476 = 14'h34a4 == index ? 14'h121 : _GEN_13475;
  wire [13:0] _GEN_13477 = 14'h34a5 == index ? 14'h11f : _GEN_13476;
  wire [13:0] _GEN_13478 = 14'h34a6 == index ? 14'h11d : _GEN_13477;
  wire [13:0] _GEN_13479 = 14'h34a7 == index ? 14'h11b : _GEN_13478;
  wire [13:0] _GEN_13480 = 14'h34a8 == index ? 14'h119 : _GEN_13479;
  wire [13:0] _GEN_13481 = 14'h34a9 == index ? 14'h117 : _GEN_13480;
  wire [13:0] _GEN_13482 = 14'h34aa == index ? 14'h115 : _GEN_13481;
  wire [13:0] _GEN_13483 = 14'h34ab == index ? 14'h113 : _GEN_13482;
  wire [13:0] _GEN_13484 = 14'h34ac == index ? 14'h111 : _GEN_13483;
  wire [13:0] _GEN_13485 = 14'h34ad == index ? 14'h10f : _GEN_13484;
  wire [13:0] _GEN_13486 = 14'h34ae == index ? 14'h10d : _GEN_13485;
  wire [13:0] _GEN_13487 = 14'h34af == index ? 14'h10b : _GEN_13486;
  wire [13:0] _GEN_13488 = 14'h34b0 == index ? 14'h109 : _GEN_13487;
  wire [13:0] _GEN_13489 = 14'h34b1 == index ? 14'h107 : _GEN_13488;
  wire [13:0] _GEN_13490 = 14'h34b2 == index ? 14'h105 : _GEN_13489;
  wire [13:0] _GEN_13491 = 14'h34b3 == index ? 14'h103 : _GEN_13490;
  wire [13:0] _GEN_13492 = 14'h34b4 == index ? 14'h101 : _GEN_13491;
  wire [13:0] _GEN_13493 = 14'h34b5 == index ? 14'hb4 : _GEN_13492;
  wire [13:0] _GEN_13494 = 14'h34b6 == index ? 14'hb3 : _GEN_13493;
  wire [13:0] _GEN_13495 = 14'h34b7 == index ? 14'hb2 : _GEN_13494;
  wire [13:0] _GEN_13496 = 14'h34b8 == index ? 14'hb1 : _GEN_13495;
  wire [13:0] _GEN_13497 = 14'h34b9 == index ? 14'hb0 : _GEN_13496;
  wire [13:0] _GEN_13498 = 14'h34ba == index ? 14'haf : _GEN_13497;
  wire [13:0] _GEN_13499 = 14'h34bb == index ? 14'hae : _GEN_13498;
  wire [13:0] _GEN_13500 = 14'h34bc == index ? 14'had : _GEN_13499;
  wire [13:0] _GEN_13501 = 14'h34bd == index ? 14'hac : _GEN_13500;
  wire [13:0] _GEN_13502 = 14'h34be == index ? 14'hab : _GEN_13501;
  wire [13:0] _GEN_13503 = 14'h34bf == index ? 14'haa : _GEN_13502;
  wire [13:0] _GEN_13504 = 14'h34c0 == index ? 14'ha9 : _GEN_13503;
  wire [13:0] _GEN_13505 = 14'h34c1 == index ? 14'ha8 : _GEN_13504;
  wire [13:0] _GEN_13506 = 14'h34c2 == index ? 14'ha7 : _GEN_13505;
  wire [13:0] _GEN_13507 = 14'h34c3 == index ? 14'ha6 : _GEN_13506;
  wire [13:0] _GEN_13508 = 14'h34c4 == index ? 14'ha5 : _GEN_13507;
  wire [13:0] _GEN_13509 = 14'h34c5 == index ? 14'ha4 : _GEN_13508;
  wire [13:0] _GEN_13510 = 14'h34c6 == index ? 14'ha3 : _GEN_13509;
  wire [13:0] _GEN_13511 = 14'h34c7 == index ? 14'ha2 : _GEN_13510;
  wire [13:0] _GEN_13512 = 14'h34c8 == index ? 14'ha1 : _GEN_13511;
  wire [13:0] _GEN_13513 = 14'h34c9 == index ? 14'ha0 : _GEN_13512;
  wire [13:0] _GEN_13514 = 14'h34ca == index ? 14'h9f : _GEN_13513;
  wire [13:0] _GEN_13515 = 14'h34cb == index ? 14'h9e : _GEN_13514;
  wire [13:0] _GEN_13516 = 14'h34cc == index ? 14'h9d : _GEN_13515;
  wire [13:0] _GEN_13517 = 14'h34cd == index ? 14'h9c : _GEN_13516;
  wire [13:0] _GEN_13518 = 14'h34ce == index ? 14'h9b : _GEN_13517;
  wire [13:0] _GEN_13519 = 14'h34cf == index ? 14'h9a : _GEN_13518;
  wire [13:0] _GEN_13520 = 14'h34d0 == index ? 14'h99 : _GEN_13519;
  wire [13:0] _GEN_13521 = 14'h34d1 == index ? 14'h98 : _GEN_13520;
  wire [13:0] _GEN_13522 = 14'h34d2 == index ? 14'h97 : _GEN_13521;
  wire [13:0] _GEN_13523 = 14'h34d3 == index ? 14'h96 : _GEN_13522;
  wire [13:0] _GEN_13524 = 14'h34d4 == index ? 14'h95 : _GEN_13523;
  wire [13:0] _GEN_13525 = 14'h34d5 == index ? 14'h94 : _GEN_13524;
  wire [13:0] _GEN_13526 = 14'h34d6 == index ? 14'h93 : _GEN_13525;
  wire [13:0] _GEN_13527 = 14'h34d7 == index ? 14'h92 : _GEN_13526;
  wire [13:0] _GEN_13528 = 14'h34d8 == index ? 14'h91 : _GEN_13527;
  wire [13:0] _GEN_13529 = 14'h34d9 == index ? 14'h90 : _GEN_13528;
  wire [13:0] _GEN_13530 = 14'h34da == index ? 14'h8f : _GEN_13529;
  wire [13:0] _GEN_13531 = 14'h34db == index ? 14'h8e : _GEN_13530;
  wire [13:0] _GEN_13532 = 14'h34dc == index ? 14'h8d : _GEN_13531;
  wire [13:0] _GEN_13533 = 14'h34dd == index ? 14'h8c : _GEN_13532;
  wire [13:0] _GEN_13534 = 14'h34de == index ? 14'h8b : _GEN_13533;
  wire [13:0] _GEN_13535 = 14'h34df == index ? 14'h8a : _GEN_13534;
  wire [13:0] _GEN_13536 = 14'h34e0 == index ? 14'h89 : _GEN_13535;
  wire [13:0] _GEN_13537 = 14'h34e1 == index ? 14'h88 : _GEN_13536;
  wire [13:0] _GEN_13538 = 14'h34e2 == index ? 14'h87 : _GEN_13537;
  wire [13:0] _GEN_13539 = 14'h34e3 == index ? 14'h86 : _GEN_13538;
  wire [13:0] _GEN_13540 = 14'h34e4 == index ? 14'h85 : _GEN_13539;
  wire [13:0] _GEN_13541 = 14'h34e5 == index ? 14'h84 : _GEN_13540;
  wire [13:0] _GEN_13542 = 14'h34e6 == index ? 14'h83 : _GEN_13541;
  wire [13:0] _GEN_13543 = 14'h34e7 == index ? 14'h82 : _GEN_13542;
  wire [13:0] _GEN_13544 = 14'h34e8 == index ? 14'h81 : _GEN_13543;
  wire [13:0] _GEN_13545 = 14'h34e9 == index ? 14'h80 : _GEN_13544;
  wire [13:0] _GEN_13546 = 14'h34ea == index ? 14'h69 : _GEN_13545;
  wire [13:0] _GEN_13547 = 14'h34eb == index ? 14'h69 : _GEN_13546;
  wire [13:0] _GEN_13548 = 14'h34ec == index ? 14'h69 : _GEN_13547;
  wire [13:0] _GEN_13549 = 14'h34ed == index ? 14'h69 : _GEN_13548;
  wire [13:0] _GEN_13550 = 14'h34ee == index ? 14'h69 : _GEN_13549;
  wire [13:0] _GEN_13551 = 14'h34ef == index ? 14'h69 : _GEN_13550;
  wire [13:0] _GEN_13552 = 14'h34f0 == index ? 14'h69 : _GEN_13551;
  wire [13:0] _GEN_13553 = 14'h34f1 == index ? 14'h69 : _GEN_13552;
  wire [13:0] _GEN_13554 = 14'h34f2 == index ? 14'h69 : _GEN_13553;
  wire [13:0] _GEN_13555 = 14'h34f3 == index ? 14'h69 : _GEN_13554;
  wire [13:0] _GEN_13556 = 14'h34f4 == index ? 14'h69 : _GEN_13555;
  wire [13:0] _GEN_13557 = 14'h34f5 == index ? 14'h69 : _GEN_13556;
  wire [13:0] _GEN_13558 = 14'h34f6 == index ? 14'h69 : _GEN_13557;
  wire [13:0] _GEN_13559 = 14'h34f7 == index ? 14'h69 : _GEN_13558;
  wire [13:0] _GEN_13560 = 14'h34f8 == index ? 14'h69 : _GEN_13559;
  wire [13:0] _GEN_13561 = 14'h34f9 == index ? 14'h69 : _GEN_13560;
  wire [13:0] _GEN_13562 = 14'h34fa == index ? 14'h69 : _GEN_13561;
  wire [13:0] _GEN_13563 = 14'h34fb == index ? 14'h69 : _GEN_13562;
  wire [13:0] _GEN_13564 = 14'h34fc == index ? 14'h69 : _GEN_13563;
  wire [13:0] _GEN_13565 = 14'h34fd == index ? 14'h69 : _GEN_13564;
  wire [13:0] _GEN_13566 = 14'h34fe == index ? 14'h69 : _GEN_13565;
  wire [13:0] _GEN_13567 = 14'h34ff == index ? 14'h69 : _GEN_13566;
  wire [13:0] _GEN_13568 = 14'h3500 == index ? 14'h0 : _GEN_13567;
  wire [13:0] _GEN_13569 = 14'h3501 == index ? 14'h3500 : _GEN_13568;
  wire [13:0] _GEN_13570 = 14'h3502 == index ? 14'h1a80 : _GEN_13569;
  wire [13:0] _GEN_13571 = 14'h3503 == index ? 14'h1181 : _GEN_13570;
  wire [13:0] _GEN_13572 = 14'h3504 == index ? 14'hd02 : _GEN_13571;
  wire [13:0] _GEN_13573 = 14'h3505 == index ? 14'ha81 : _GEN_13572;
  wire [13:0] _GEN_13574 = 14'h3506 == index ? 14'h884 : _GEN_13573;
  wire [13:0] _GEN_13575 = 14'h3507 == index ? 14'h781 : _GEN_13574;
  wire [13:0] _GEN_13576 = 14'h3508 == index ? 14'h682 : _GEN_13575;
  wire [13:0] _GEN_13577 = 14'h3509 == index ? 14'h587 : _GEN_13576;
  wire [13:0] _GEN_13578 = 14'h350a == index ? 14'h506 : _GEN_13577;
  wire [13:0] _GEN_13579 = 14'h350b == index ? 14'h487 : _GEN_13578;
  wire [13:0] _GEN_13580 = 14'h350c == index ? 14'h40a : _GEN_13579;
  wire [13:0] _GEN_13581 = 14'h350d == index ? 14'h402 : _GEN_13580;
  wire [13:0] _GEN_13582 = 14'h350e == index ? 14'h388 : _GEN_13581;
  wire [13:0] _GEN_13583 = 14'h350f == index ? 14'h381 : _GEN_13582;
  wire [13:0] _GEN_13584 = 14'h3510 == index ? 14'h30a : _GEN_13583;
  wire [13:0] _GEN_13585 = 14'h3511 == index ? 14'h304 : _GEN_13584;
  wire [13:0] _GEN_13586 = 14'h3512 == index ? 14'h290 : _GEN_13585;
  wire [13:0] _GEN_13587 = 14'h3513 == index ? 14'h28b : _GEN_13586;
  wire [13:0] _GEN_13588 = 14'h3514 == index ? 14'h286 : _GEN_13587;
  wire [13:0] _GEN_13589 = 14'h3515 == index ? 14'h281 : _GEN_13588;
  wire [13:0] _GEN_13590 = 14'h3516 == index ? 14'h212 : _GEN_13589;
  wire [13:0] _GEN_13591 = 14'h3517 == index ? 14'h20e : _GEN_13590;
  wire [13:0] _GEN_13592 = 14'h3518 == index ? 14'h20a : _GEN_13591;
  wire [13:0] _GEN_13593 = 14'h3519 == index ? 14'h206 : _GEN_13592;
  wire [13:0] _GEN_13594 = 14'h351a == index ? 14'h202 : _GEN_13593;
  wire [13:0] _GEN_13595 = 14'h351b == index ? 14'h199 : _GEN_13594;
  wire [13:0] _GEN_13596 = 14'h351c == index ? 14'h196 : _GEN_13595;
  wire [13:0] _GEN_13597 = 14'h351d == index ? 14'h193 : _GEN_13596;
  wire [13:0] _GEN_13598 = 14'h351e == index ? 14'h190 : _GEN_13597;
  wire [13:0] _GEN_13599 = 14'h351f == index ? 14'h18d : _GEN_13598;
  wire [13:0] _GEN_13600 = 14'h3520 == index ? 14'h18a : _GEN_13599;
  wire [13:0] _GEN_13601 = 14'h3521 == index ? 14'h187 : _GEN_13600;
  wire [13:0] _GEN_13602 = 14'h3522 == index ? 14'h184 : _GEN_13601;
  wire [13:0] _GEN_13603 = 14'h3523 == index ? 14'h181 : _GEN_13602;
  wire [13:0] _GEN_13604 = 14'h3524 == index ? 14'h122 : _GEN_13603;
  wire [13:0] _GEN_13605 = 14'h3525 == index ? 14'h120 : _GEN_13604;
  wire [13:0] _GEN_13606 = 14'h3526 == index ? 14'h11e : _GEN_13605;
  wire [13:0] _GEN_13607 = 14'h3527 == index ? 14'h11c : _GEN_13606;
  wire [13:0] _GEN_13608 = 14'h3528 == index ? 14'h11a : _GEN_13607;
  wire [13:0] _GEN_13609 = 14'h3529 == index ? 14'h118 : _GEN_13608;
  wire [13:0] _GEN_13610 = 14'h352a == index ? 14'h116 : _GEN_13609;
  wire [13:0] _GEN_13611 = 14'h352b == index ? 14'h114 : _GEN_13610;
  wire [13:0] _GEN_13612 = 14'h352c == index ? 14'h112 : _GEN_13611;
  wire [13:0] _GEN_13613 = 14'h352d == index ? 14'h110 : _GEN_13612;
  wire [13:0] _GEN_13614 = 14'h352e == index ? 14'h10e : _GEN_13613;
  wire [13:0] _GEN_13615 = 14'h352f == index ? 14'h10c : _GEN_13614;
  wire [13:0] _GEN_13616 = 14'h3530 == index ? 14'h10a : _GEN_13615;
  wire [13:0] _GEN_13617 = 14'h3531 == index ? 14'h108 : _GEN_13616;
  wire [13:0] _GEN_13618 = 14'h3532 == index ? 14'h106 : _GEN_13617;
  wire [13:0] _GEN_13619 = 14'h3533 == index ? 14'h104 : _GEN_13618;
  wire [13:0] _GEN_13620 = 14'h3534 == index ? 14'h102 : _GEN_13619;
  wire [13:0] _GEN_13621 = 14'h3535 == index ? 14'h100 : _GEN_13620;
  wire [13:0] _GEN_13622 = 14'h3536 == index ? 14'hb4 : _GEN_13621;
  wire [13:0] _GEN_13623 = 14'h3537 == index ? 14'hb3 : _GEN_13622;
  wire [13:0] _GEN_13624 = 14'h3538 == index ? 14'hb2 : _GEN_13623;
  wire [13:0] _GEN_13625 = 14'h3539 == index ? 14'hb1 : _GEN_13624;
  wire [13:0] _GEN_13626 = 14'h353a == index ? 14'hb0 : _GEN_13625;
  wire [13:0] _GEN_13627 = 14'h353b == index ? 14'haf : _GEN_13626;
  wire [13:0] _GEN_13628 = 14'h353c == index ? 14'hae : _GEN_13627;
  wire [13:0] _GEN_13629 = 14'h353d == index ? 14'had : _GEN_13628;
  wire [13:0] _GEN_13630 = 14'h353e == index ? 14'hac : _GEN_13629;
  wire [13:0] _GEN_13631 = 14'h353f == index ? 14'hab : _GEN_13630;
  wire [13:0] _GEN_13632 = 14'h3540 == index ? 14'haa : _GEN_13631;
  wire [13:0] _GEN_13633 = 14'h3541 == index ? 14'ha9 : _GEN_13632;
  wire [13:0] _GEN_13634 = 14'h3542 == index ? 14'ha8 : _GEN_13633;
  wire [13:0] _GEN_13635 = 14'h3543 == index ? 14'ha7 : _GEN_13634;
  wire [13:0] _GEN_13636 = 14'h3544 == index ? 14'ha6 : _GEN_13635;
  wire [13:0] _GEN_13637 = 14'h3545 == index ? 14'ha5 : _GEN_13636;
  wire [13:0] _GEN_13638 = 14'h3546 == index ? 14'ha4 : _GEN_13637;
  wire [13:0] _GEN_13639 = 14'h3547 == index ? 14'ha3 : _GEN_13638;
  wire [13:0] _GEN_13640 = 14'h3548 == index ? 14'ha2 : _GEN_13639;
  wire [13:0] _GEN_13641 = 14'h3549 == index ? 14'ha1 : _GEN_13640;
  wire [13:0] _GEN_13642 = 14'h354a == index ? 14'ha0 : _GEN_13641;
  wire [13:0] _GEN_13643 = 14'h354b == index ? 14'h9f : _GEN_13642;
  wire [13:0] _GEN_13644 = 14'h354c == index ? 14'h9e : _GEN_13643;
  wire [13:0] _GEN_13645 = 14'h354d == index ? 14'h9d : _GEN_13644;
  wire [13:0] _GEN_13646 = 14'h354e == index ? 14'h9c : _GEN_13645;
  wire [13:0] _GEN_13647 = 14'h354f == index ? 14'h9b : _GEN_13646;
  wire [13:0] _GEN_13648 = 14'h3550 == index ? 14'h9a : _GEN_13647;
  wire [13:0] _GEN_13649 = 14'h3551 == index ? 14'h99 : _GEN_13648;
  wire [13:0] _GEN_13650 = 14'h3552 == index ? 14'h98 : _GEN_13649;
  wire [13:0] _GEN_13651 = 14'h3553 == index ? 14'h97 : _GEN_13650;
  wire [13:0] _GEN_13652 = 14'h3554 == index ? 14'h96 : _GEN_13651;
  wire [13:0] _GEN_13653 = 14'h3555 == index ? 14'h95 : _GEN_13652;
  wire [13:0] _GEN_13654 = 14'h3556 == index ? 14'h94 : _GEN_13653;
  wire [13:0] _GEN_13655 = 14'h3557 == index ? 14'h93 : _GEN_13654;
  wire [13:0] _GEN_13656 = 14'h3558 == index ? 14'h92 : _GEN_13655;
  wire [13:0] _GEN_13657 = 14'h3559 == index ? 14'h91 : _GEN_13656;
  wire [13:0] _GEN_13658 = 14'h355a == index ? 14'h90 : _GEN_13657;
  wire [13:0] _GEN_13659 = 14'h355b == index ? 14'h8f : _GEN_13658;
  wire [13:0] _GEN_13660 = 14'h355c == index ? 14'h8e : _GEN_13659;
  wire [13:0] _GEN_13661 = 14'h355d == index ? 14'h8d : _GEN_13660;
  wire [13:0] _GEN_13662 = 14'h355e == index ? 14'h8c : _GEN_13661;
  wire [13:0] _GEN_13663 = 14'h355f == index ? 14'h8b : _GEN_13662;
  wire [13:0] _GEN_13664 = 14'h3560 == index ? 14'h8a : _GEN_13663;
  wire [13:0] _GEN_13665 = 14'h3561 == index ? 14'h89 : _GEN_13664;
  wire [13:0] _GEN_13666 = 14'h3562 == index ? 14'h88 : _GEN_13665;
  wire [13:0] _GEN_13667 = 14'h3563 == index ? 14'h87 : _GEN_13666;
  wire [13:0] _GEN_13668 = 14'h3564 == index ? 14'h86 : _GEN_13667;
  wire [13:0] _GEN_13669 = 14'h3565 == index ? 14'h85 : _GEN_13668;
  wire [13:0] _GEN_13670 = 14'h3566 == index ? 14'h84 : _GEN_13669;
  wire [13:0] _GEN_13671 = 14'h3567 == index ? 14'h83 : _GEN_13670;
  wire [13:0] _GEN_13672 = 14'h3568 == index ? 14'h82 : _GEN_13671;
  wire [13:0] _GEN_13673 = 14'h3569 == index ? 14'h81 : _GEN_13672;
  wire [13:0] _GEN_13674 = 14'h356a == index ? 14'h80 : _GEN_13673;
  wire [13:0] _GEN_13675 = 14'h356b == index ? 14'h6a : _GEN_13674;
  wire [13:0] _GEN_13676 = 14'h356c == index ? 14'h6a : _GEN_13675;
  wire [13:0] _GEN_13677 = 14'h356d == index ? 14'h6a : _GEN_13676;
  wire [13:0] _GEN_13678 = 14'h356e == index ? 14'h6a : _GEN_13677;
  wire [13:0] _GEN_13679 = 14'h356f == index ? 14'h6a : _GEN_13678;
  wire [13:0] _GEN_13680 = 14'h3570 == index ? 14'h6a : _GEN_13679;
  wire [13:0] _GEN_13681 = 14'h3571 == index ? 14'h6a : _GEN_13680;
  wire [13:0] _GEN_13682 = 14'h3572 == index ? 14'h6a : _GEN_13681;
  wire [13:0] _GEN_13683 = 14'h3573 == index ? 14'h6a : _GEN_13682;
  wire [13:0] _GEN_13684 = 14'h3574 == index ? 14'h6a : _GEN_13683;
  wire [13:0] _GEN_13685 = 14'h3575 == index ? 14'h6a : _GEN_13684;
  wire [13:0] _GEN_13686 = 14'h3576 == index ? 14'h6a : _GEN_13685;
  wire [13:0] _GEN_13687 = 14'h3577 == index ? 14'h6a : _GEN_13686;
  wire [13:0] _GEN_13688 = 14'h3578 == index ? 14'h6a : _GEN_13687;
  wire [13:0] _GEN_13689 = 14'h3579 == index ? 14'h6a : _GEN_13688;
  wire [13:0] _GEN_13690 = 14'h357a == index ? 14'h6a : _GEN_13689;
  wire [13:0] _GEN_13691 = 14'h357b == index ? 14'h6a : _GEN_13690;
  wire [13:0] _GEN_13692 = 14'h357c == index ? 14'h6a : _GEN_13691;
  wire [13:0] _GEN_13693 = 14'h357d == index ? 14'h6a : _GEN_13692;
  wire [13:0] _GEN_13694 = 14'h357e == index ? 14'h6a : _GEN_13693;
  wire [13:0] _GEN_13695 = 14'h357f == index ? 14'h6a : _GEN_13694;
  wire [13:0] _GEN_13696 = 14'h3580 == index ? 14'h0 : _GEN_13695;
  wire [13:0] _GEN_13697 = 14'h3581 == index ? 14'h3580 : _GEN_13696;
  wire [13:0] _GEN_13698 = 14'h3582 == index ? 14'h1a81 : _GEN_13697;
  wire [13:0] _GEN_13699 = 14'h3583 == index ? 14'h1182 : _GEN_13698;
  wire [13:0] _GEN_13700 = 14'h3584 == index ? 14'hd03 : _GEN_13699;
  wire [13:0] _GEN_13701 = 14'h3585 == index ? 14'ha82 : _GEN_13700;
  wire [13:0] _GEN_13702 = 14'h3586 == index ? 14'h885 : _GEN_13701;
  wire [13:0] _GEN_13703 = 14'h3587 == index ? 14'h782 : _GEN_13702;
  wire [13:0] _GEN_13704 = 14'h3588 == index ? 14'h683 : _GEN_13703;
  wire [13:0] _GEN_13705 = 14'h3589 == index ? 14'h588 : _GEN_13704;
  wire [13:0] _GEN_13706 = 14'h358a == index ? 14'h507 : _GEN_13705;
  wire [13:0] _GEN_13707 = 14'h358b == index ? 14'h488 : _GEN_13706;
  wire [13:0] _GEN_13708 = 14'h358c == index ? 14'h40b : _GEN_13707;
  wire [13:0] _GEN_13709 = 14'h358d == index ? 14'h403 : _GEN_13708;
  wire [13:0] _GEN_13710 = 14'h358e == index ? 14'h389 : _GEN_13709;
  wire [13:0] _GEN_13711 = 14'h358f == index ? 14'h382 : _GEN_13710;
  wire [13:0] _GEN_13712 = 14'h3590 == index ? 14'h30b : _GEN_13711;
  wire [13:0] _GEN_13713 = 14'h3591 == index ? 14'h305 : _GEN_13712;
  wire [13:0] _GEN_13714 = 14'h3592 == index ? 14'h291 : _GEN_13713;
  wire [13:0] _GEN_13715 = 14'h3593 == index ? 14'h28c : _GEN_13714;
  wire [13:0] _GEN_13716 = 14'h3594 == index ? 14'h287 : _GEN_13715;
  wire [13:0] _GEN_13717 = 14'h3595 == index ? 14'h282 : _GEN_13716;
  wire [13:0] _GEN_13718 = 14'h3596 == index ? 14'h213 : _GEN_13717;
  wire [13:0] _GEN_13719 = 14'h3597 == index ? 14'h20f : _GEN_13718;
  wire [13:0] _GEN_13720 = 14'h3598 == index ? 14'h20b : _GEN_13719;
  wire [13:0] _GEN_13721 = 14'h3599 == index ? 14'h207 : _GEN_13720;
  wire [13:0] _GEN_13722 = 14'h359a == index ? 14'h203 : _GEN_13721;
  wire [13:0] _GEN_13723 = 14'h359b == index ? 14'h19a : _GEN_13722;
  wire [13:0] _GEN_13724 = 14'h359c == index ? 14'h197 : _GEN_13723;
  wire [13:0] _GEN_13725 = 14'h359d == index ? 14'h194 : _GEN_13724;
  wire [13:0] _GEN_13726 = 14'h359e == index ? 14'h191 : _GEN_13725;
  wire [13:0] _GEN_13727 = 14'h359f == index ? 14'h18e : _GEN_13726;
  wire [13:0] _GEN_13728 = 14'h35a0 == index ? 14'h18b : _GEN_13727;
  wire [13:0] _GEN_13729 = 14'h35a1 == index ? 14'h188 : _GEN_13728;
  wire [13:0] _GEN_13730 = 14'h35a2 == index ? 14'h185 : _GEN_13729;
  wire [13:0] _GEN_13731 = 14'h35a3 == index ? 14'h182 : _GEN_13730;
  wire [13:0] _GEN_13732 = 14'h35a4 == index ? 14'h123 : _GEN_13731;
  wire [13:0] _GEN_13733 = 14'h35a5 == index ? 14'h121 : _GEN_13732;
  wire [13:0] _GEN_13734 = 14'h35a6 == index ? 14'h11f : _GEN_13733;
  wire [13:0] _GEN_13735 = 14'h35a7 == index ? 14'h11d : _GEN_13734;
  wire [13:0] _GEN_13736 = 14'h35a8 == index ? 14'h11b : _GEN_13735;
  wire [13:0] _GEN_13737 = 14'h35a9 == index ? 14'h119 : _GEN_13736;
  wire [13:0] _GEN_13738 = 14'h35aa == index ? 14'h117 : _GEN_13737;
  wire [13:0] _GEN_13739 = 14'h35ab == index ? 14'h115 : _GEN_13738;
  wire [13:0] _GEN_13740 = 14'h35ac == index ? 14'h113 : _GEN_13739;
  wire [13:0] _GEN_13741 = 14'h35ad == index ? 14'h111 : _GEN_13740;
  wire [13:0] _GEN_13742 = 14'h35ae == index ? 14'h10f : _GEN_13741;
  wire [13:0] _GEN_13743 = 14'h35af == index ? 14'h10d : _GEN_13742;
  wire [13:0] _GEN_13744 = 14'h35b0 == index ? 14'h10b : _GEN_13743;
  wire [13:0] _GEN_13745 = 14'h35b1 == index ? 14'h109 : _GEN_13744;
  wire [13:0] _GEN_13746 = 14'h35b2 == index ? 14'h107 : _GEN_13745;
  wire [13:0] _GEN_13747 = 14'h35b3 == index ? 14'h105 : _GEN_13746;
  wire [13:0] _GEN_13748 = 14'h35b4 == index ? 14'h103 : _GEN_13747;
  wire [13:0] _GEN_13749 = 14'h35b5 == index ? 14'h101 : _GEN_13748;
  wire [13:0] _GEN_13750 = 14'h35b6 == index ? 14'hb5 : _GEN_13749;
  wire [13:0] _GEN_13751 = 14'h35b7 == index ? 14'hb4 : _GEN_13750;
  wire [13:0] _GEN_13752 = 14'h35b8 == index ? 14'hb3 : _GEN_13751;
  wire [13:0] _GEN_13753 = 14'h35b9 == index ? 14'hb2 : _GEN_13752;
  wire [13:0] _GEN_13754 = 14'h35ba == index ? 14'hb1 : _GEN_13753;
  wire [13:0] _GEN_13755 = 14'h35bb == index ? 14'hb0 : _GEN_13754;
  wire [13:0] _GEN_13756 = 14'h35bc == index ? 14'haf : _GEN_13755;
  wire [13:0] _GEN_13757 = 14'h35bd == index ? 14'hae : _GEN_13756;
  wire [13:0] _GEN_13758 = 14'h35be == index ? 14'had : _GEN_13757;
  wire [13:0] _GEN_13759 = 14'h35bf == index ? 14'hac : _GEN_13758;
  wire [13:0] _GEN_13760 = 14'h35c0 == index ? 14'hab : _GEN_13759;
  wire [13:0] _GEN_13761 = 14'h35c1 == index ? 14'haa : _GEN_13760;
  wire [13:0] _GEN_13762 = 14'h35c2 == index ? 14'ha9 : _GEN_13761;
  wire [13:0] _GEN_13763 = 14'h35c3 == index ? 14'ha8 : _GEN_13762;
  wire [13:0] _GEN_13764 = 14'h35c4 == index ? 14'ha7 : _GEN_13763;
  wire [13:0] _GEN_13765 = 14'h35c5 == index ? 14'ha6 : _GEN_13764;
  wire [13:0] _GEN_13766 = 14'h35c6 == index ? 14'ha5 : _GEN_13765;
  wire [13:0] _GEN_13767 = 14'h35c7 == index ? 14'ha4 : _GEN_13766;
  wire [13:0] _GEN_13768 = 14'h35c8 == index ? 14'ha3 : _GEN_13767;
  wire [13:0] _GEN_13769 = 14'h35c9 == index ? 14'ha2 : _GEN_13768;
  wire [13:0] _GEN_13770 = 14'h35ca == index ? 14'ha1 : _GEN_13769;
  wire [13:0] _GEN_13771 = 14'h35cb == index ? 14'ha0 : _GEN_13770;
  wire [13:0] _GEN_13772 = 14'h35cc == index ? 14'h9f : _GEN_13771;
  wire [13:0] _GEN_13773 = 14'h35cd == index ? 14'h9e : _GEN_13772;
  wire [13:0] _GEN_13774 = 14'h35ce == index ? 14'h9d : _GEN_13773;
  wire [13:0] _GEN_13775 = 14'h35cf == index ? 14'h9c : _GEN_13774;
  wire [13:0] _GEN_13776 = 14'h35d0 == index ? 14'h9b : _GEN_13775;
  wire [13:0] _GEN_13777 = 14'h35d1 == index ? 14'h9a : _GEN_13776;
  wire [13:0] _GEN_13778 = 14'h35d2 == index ? 14'h99 : _GEN_13777;
  wire [13:0] _GEN_13779 = 14'h35d3 == index ? 14'h98 : _GEN_13778;
  wire [13:0] _GEN_13780 = 14'h35d4 == index ? 14'h97 : _GEN_13779;
  wire [13:0] _GEN_13781 = 14'h35d5 == index ? 14'h96 : _GEN_13780;
  wire [13:0] _GEN_13782 = 14'h35d6 == index ? 14'h95 : _GEN_13781;
  wire [13:0] _GEN_13783 = 14'h35d7 == index ? 14'h94 : _GEN_13782;
  wire [13:0] _GEN_13784 = 14'h35d8 == index ? 14'h93 : _GEN_13783;
  wire [13:0] _GEN_13785 = 14'h35d9 == index ? 14'h92 : _GEN_13784;
  wire [13:0] _GEN_13786 = 14'h35da == index ? 14'h91 : _GEN_13785;
  wire [13:0] _GEN_13787 = 14'h35db == index ? 14'h90 : _GEN_13786;
  wire [13:0] _GEN_13788 = 14'h35dc == index ? 14'h8f : _GEN_13787;
  wire [13:0] _GEN_13789 = 14'h35dd == index ? 14'h8e : _GEN_13788;
  wire [13:0] _GEN_13790 = 14'h35de == index ? 14'h8d : _GEN_13789;
  wire [13:0] _GEN_13791 = 14'h35df == index ? 14'h8c : _GEN_13790;
  wire [13:0] _GEN_13792 = 14'h35e0 == index ? 14'h8b : _GEN_13791;
  wire [13:0] _GEN_13793 = 14'h35e1 == index ? 14'h8a : _GEN_13792;
  wire [13:0] _GEN_13794 = 14'h35e2 == index ? 14'h89 : _GEN_13793;
  wire [13:0] _GEN_13795 = 14'h35e3 == index ? 14'h88 : _GEN_13794;
  wire [13:0] _GEN_13796 = 14'h35e4 == index ? 14'h87 : _GEN_13795;
  wire [13:0] _GEN_13797 = 14'h35e5 == index ? 14'h86 : _GEN_13796;
  wire [13:0] _GEN_13798 = 14'h35e6 == index ? 14'h85 : _GEN_13797;
  wire [13:0] _GEN_13799 = 14'h35e7 == index ? 14'h84 : _GEN_13798;
  wire [13:0] _GEN_13800 = 14'h35e8 == index ? 14'h83 : _GEN_13799;
  wire [13:0] _GEN_13801 = 14'h35e9 == index ? 14'h82 : _GEN_13800;
  wire [13:0] _GEN_13802 = 14'h35ea == index ? 14'h81 : _GEN_13801;
  wire [13:0] _GEN_13803 = 14'h35eb == index ? 14'h80 : _GEN_13802;
  wire [13:0] _GEN_13804 = 14'h35ec == index ? 14'h6b : _GEN_13803;
  wire [13:0] _GEN_13805 = 14'h35ed == index ? 14'h6b : _GEN_13804;
  wire [13:0] _GEN_13806 = 14'h35ee == index ? 14'h6b : _GEN_13805;
  wire [13:0] _GEN_13807 = 14'h35ef == index ? 14'h6b : _GEN_13806;
  wire [13:0] _GEN_13808 = 14'h35f0 == index ? 14'h6b : _GEN_13807;
  wire [13:0] _GEN_13809 = 14'h35f1 == index ? 14'h6b : _GEN_13808;
  wire [13:0] _GEN_13810 = 14'h35f2 == index ? 14'h6b : _GEN_13809;
  wire [13:0] _GEN_13811 = 14'h35f3 == index ? 14'h6b : _GEN_13810;
  wire [13:0] _GEN_13812 = 14'h35f4 == index ? 14'h6b : _GEN_13811;
  wire [13:0] _GEN_13813 = 14'h35f5 == index ? 14'h6b : _GEN_13812;
  wire [13:0] _GEN_13814 = 14'h35f6 == index ? 14'h6b : _GEN_13813;
  wire [13:0] _GEN_13815 = 14'h35f7 == index ? 14'h6b : _GEN_13814;
  wire [13:0] _GEN_13816 = 14'h35f8 == index ? 14'h6b : _GEN_13815;
  wire [13:0] _GEN_13817 = 14'h35f9 == index ? 14'h6b : _GEN_13816;
  wire [13:0] _GEN_13818 = 14'h35fa == index ? 14'h6b : _GEN_13817;
  wire [13:0] _GEN_13819 = 14'h35fb == index ? 14'h6b : _GEN_13818;
  wire [13:0] _GEN_13820 = 14'h35fc == index ? 14'h6b : _GEN_13819;
  wire [13:0] _GEN_13821 = 14'h35fd == index ? 14'h6b : _GEN_13820;
  wire [13:0] _GEN_13822 = 14'h35fe == index ? 14'h6b : _GEN_13821;
  wire [13:0] _GEN_13823 = 14'h35ff == index ? 14'h6b : _GEN_13822;
  wire [13:0] _GEN_13824 = 14'h3600 == index ? 14'h0 : _GEN_13823;
  wire [13:0] _GEN_13825 = 14'h3601 == index ? 14'h3600 : _GEN_13824;
  wire [13:0] _GEN_13826 = 14'h3602 == index ? 14'h1b00 : _GEN_13825;
  wire [13:0] _GEN_13827 = 14'h3603 == index ? 14'h1200 : _GEN_13826;
  wire [13:0] _GEN_13828 = 14'h3604 == index ? 14'hd80 : _GEN_13827;
  wire [13:0] _GEN_13829 = 14'h3605 == index ? 14'ha83 : _GEN_13828;
  wire [13:0] _GEN_13830 = 14'h3606 == index ? 14'h900 : _GEN_13829;
  wire [13:0] _GEN_13831 = 14'h3607 == index ? 14'h783 : _GEN_13830;
  wire [13:0] _GEN_13832 = 14'h3608 == index ? 14'h684 : _GEN_13831;
  wire [13:0] _GEN_13833 = 14'h3609 == index ? 14'h600 : _GEN_13832;
  wire [13:0] _GEN_13834 = 14'h360a == index ? 14'h508 : _GEN_13833;
  wire [13:0] _GEN_13835 = 14'h360b == index ? 14'h489 : _GEN_13834;
  wire [13:0] _GEN_13836 = 14'h360c == index ? 14'h480 : _GEN_13835;
  wire [13:0] _GEN_13837 = 14'h360d == index ? 14'h404 : _GEN_13836;
  wire [13:0] _GEN_13838 = 14'h360e == index ? 14'h38a : _GEN_13837;
  wire [13:0] _GEN_13839 = 14'h360f == index ? 14'h383 : _GEN_13838;
  wire [13:0] _GEN_13840 = 14'h3610 == index ? 14'h30c : _GEN_13839;
  wire [13:0] _GEN_13841 = 14'h3611 == index ? 14'h306 : _GEN_13840;
  wire [13:0] _GEN_13842 = 14'h3612 == index ? 14'h300 : _GEN_13841;
  wire [13:0] _GEN_13843 = 14'h3613 == index ? 14'h28d : _GEN_13842;
  wire [13:0] _GEN_13844 = 14'h3614 == index ? 14'h288 : _GEN_13843;
  wire [13:0] _GEN_13845 = 14'h3615 == index ? 14'h283 : _GEN_13844;
  wire [13:0] _GEN_13846 = 14'h3616 == index ? 14'h214 : _GEN_13845;
  wire [13:0] _GEN_13847 = 14'h3617 == index ? 14'h210 : _GEN_13846;
  wire [13:0] _GEN_13848 = 14'h3618 == index ? 14'h20c : _GEN_13847;
  wire [13:0] _GEN_13849 = 14'h3619 == index ? 14'h208 : _GEN_13848;
  wire [13:0] _GEN_13850 = 14'h361a == index ? 14'h204 : _GEN_13849;
  wire [13:0] _GEN_13851 = 14'h361b == index ? 14'h200 : _GEN_13850;
  wire [13:0] _GEN_13852 = 14'h361c == index ? 14'h198 : _GEN_13851;
  wire [13:0] _GEN_13853 = 14'h361d == index ? 14'h195 : _GEN_13852;
  wire [13:0] _GEN_13854 = 14'h361e == index ? 14'h192 : _GEN_13853;
  wire [13:0] _GEN_13855 = 14'h361f == index ? 14'h18f : _GEN_13854;
  wire [13:0] _GEN_13856 = 14'h3620 == index ? 14'h18c : _GEN_13855;
  wire [13:0] _GEN_13857 = 14'h3621 == index ? 14'h189 : _GEN_13856;
  wire [13:0] _GEN_13858 = 14'h3622 == index ? 14'h186 : _GEN_13857;
  wire [13:0] _GEN_13859 = 14'h3623 == index ? 14'h183 : _GEN_13858;
  wire [13:0] _GEN_13860 = 14'h3624 == index ? 14'h180 : _GEN_13859;
  wire [13:0] _GEN_13861 = 14'h3625 == index ? 14'h122 : _GEN_13860;
  wire [13:0] _GEN_13862 = 14'h3626 == index ? 14'h120 : _GEN_13861;
  wire [13:0] _GEN_13863 = 14'h3627 == index ? 14'h11e : _GEN_13862;
  wire [13:0] _GEN_13864 = 14'h3628 == index ? 14'h11c : _GEN_13863;
  wire [13:0] _GEN_13865 = 14'h3629 == index ? 14'h11a : _GEN_13864;
  wire [13:0] _GEN_13866 = 14'h362a == index ? 14'h118 : _GEN_13865;
  wire [13:0] _GEN_13867 = 14'h362b == index ? 14'h116 : _GEN_13866;
  wire [13:0] _GEN_13868 = 14'h362c == index ? 14'h114 : _GEN_13867;
  wire [13:0] _GEN_13869 = 14'h362d == index ? 14'h112 : _GEN_13868;
  wire [13:0] _GEN_13870 = 14'h362e == index ? 14'h110 : _GEN_13869;
  wire [13:0] _GEN_13871 = 14'h362f == index ? 14'h10e : _GEN_13870;
  wire [13:0] _GEN_13872 = 14'h3630 == index ? 14'h10c : _GEN_13871;
  wire [13:0] _GEN_13873 = 14'h3631 == index ? 14'h10a : _GEN_13872;
  wire [13:0] _GEN_13874 = 14'h3632 == index ? 14'h108 : _GEN_13873;
  wire [13:0] _GEN_13875 = 14'h3633 == index ? 14'h106 : _GEN_13874;
  wire [13:0] _GEN_13876 = 14'h3634 == index ? 14'h104 : _GEN_13875;
  wire [13:0] _GEN_13877 = 14'h3635 == index ? 14'h102 : _GEN_13876;
  wire [13:0] _GEN_13878 = 14'h3636 == index ? 14'h100 : _GEN_13877;
  wire [13:0] _GEN_13879 = 14'h3637 == index ? 14'hb5 : _GEN_13878;
  wire [13:0] _GEN_13880 = 14'h3638 == index ? 14'hb4 : _GEN_13879;
  wire [13:0] _GEN_13881 = 14'h3639 == index ? 14'hb3 : _GEN_13880;
  wire [13:0] _GEN_13882 = 14'h363a == index ? 14'hb2 : _GEN_13881;
  wire [13:0] _GEN_13883 = 14'h363b == index ? 14'hb1 : _GEN_13882;
  wire [13:0] _GEN_13884 = 14'h363c == index ? 14'hb0 : _GEN_13883;
  wire [13:0] _GEN_13885 = 14'h363d == index ? 14'haf : _GEN_13884;
  wire [13:0] _GEN_13886 = 14'h363e == index ? 14'hae : _GEN_13885;
  wire [13:0] _GEN_13887 = 14'h363f == index ? 14'had : _GEN_13886;
  wire [13:0] _GEN_13888 = 14'h3640 == index ? 14'hac : _GEN_13887;
  wire [13:0] _GEN_13889 = 14'h3641 == index ? 14'hab : _GEN_13888;
  wire [13:0] _GEN_13890 = 14'h3642 == index ? 14'haa : _GEN_13889;
  wire [13:0] _GEN_13891 = 14'h3643 == index ? 14'ha9 : _GEN_13890;
  wire [13:0] _GEN_13892 = 14'h3644 == index ? 14'ha8 : _GEN_13891;
  wire [13:0] _GEN_13893 = 14'h3645 == index ? 14'ha7 : _GEN_13892;
  wire [13:0] _GEN_13894 = 14'h3646 == index ? 14'ha6 : _GEN_13893;
  wire [13:0] _GEN_13895 = 14'h3647 == index ? 14'ha5 : _GEN_13894;
  wire [13:0] _GEN_13896 = 14'h3648 == index ? 14'ha4 : _GEN_13895;
  wire [13:0] _GEN_13897 = 14'h3649 == index ? 14'ha3 : _GEN_13896;
  wire [13:0] _GEN_13898 = 14'h364a == index ? 14'ha2 : _GEN_13897;
  wire [13:0] _GEN_13899 = 14'h364b == index ? 14'ha1 : _GEN_13898;
  wire [13:0] _GEN_13900 = 14'h364c == index ? 14'ha0 : _GEN_13899;
  wire [13:0] _GEN_13901 = 14'h364d == index ? 14'h9f : _GEN_13900;
  wire [13:0] _GEN_13902 = 14'h364e == index ? 14'h9e : _GEN_13901;
  wire [13:0] _GEN_13903 = 14'h364f == index ? 14'h9d : _GEN_13902;
  wire [13:0] _GEN_13904 = 14'h3650 == index ? 14'h9c : _GEN_13903;
  wire [13:0] _GEN_13905 = 14'h3651 == index ? 14'h9b : _GEN_13904;
  wire [13:0] _GEN_13906 = 14'h3652 == index ? 14'h9a : _GEN_13905;
  wire [13:0] _GEN_13907 = 14'h3653 == index ? 14'h99 : _GEN_13906;
  wire [13:0] _GEN_13908 = 14'h3654 == index ? 14'h98 : _GEN_13907;
  wire [13:0] _GEN_13909 = 14'h3655 == index ? 14'h97 : _GEN_13908;
  wire [13:0] _GEN_13910 = 14'h3656 == index ? 14'h96 : _GEN_13909;
  wire [13:0] _GEN_13911 = 14'h3657 == index ? 14'h95 : _GEN_13910;
  wire [13:0] _GEN_13912 = 14'h3658 == index ? 14'h94 : _GEN_13911;
  wire [13:0] _GEN_13913 = 14'h3659 == index ? 14'h93 : _GEN_13912;
  wire [13:0] _GEN_13914 = 14'h365a == index ? 14'h92 : _GEN_13913;
  wire [13:0] _GEN_13915 = 14'h365b == index ? 14'h91 : _GEN_13914;
  wire [13:0] _GEN_13916 = 14'h365c == index ? 14'h90 : _GEN_13915;
  wire [13:0] _GEN_13917 = 14'h365d == index ? 14'h8f : _GEN_13916;
  wire [13:0] _GEN_13918 = 14'h365e == index ? 14'h8e : _GEN_13917;
  wire [13:0] _GEN_13919 = 14'h365f == index ? 14'h8d : _GEN_13918;
  wire [13:0] _GEN_13920 = 14'h3660 == index ? 14'h8c : _GEN_13919;
  wire [13:0] _GEN_13921 = 14'h3661 == index ? 14'h8b : _GEN_13920;
  wire [13:0] _GEN_13922 = 14'h3662 == index ? 14'h8a : _GEN_13921;
  wire [13:0] _GEN_13923 = 14'h3663 == index ? 14'h89 : _GEN_13922;
  wire [13:0] _GEN_13924 = 14'h3664 == index ? 14'h88 : _GEN_13923;
  wire [13:0] _GEN_13925 = 14'h3665 == index ? 14'h87 : _GEN_13924;
  wire [13:0] _GEN_13926 = 14'h3666 == index ? 14'h86 : _GEN_13925;
  wire [13:0] _GEN_13927 = 14'h3667 == index ? 14'h85 : _GEN_13926;
  wire [13:0] _GEN_13928 = 14'h3668 == index ? 14'h84 : _GEN_13927;
  wire [13:0] _GEN_13929 = 14'h3669 == index ? 14'h83 : _GEN_13928;
  wire [13:0] _GEN_13930 = 14'h366a == index ? 14'h82 : _GEN_13929;
  wire [13:0] _GEN_13931 = 14'h366b == index ? 14'h81 : _GEN_13930;
  wire [13:0] _GEN_13932 = 14'h366c == index ? 14'h80 : _GEN_13931;
  wire [13:0] _GEN_13933 = 14'h366d == index ? 14'h6c : _GEN_13932;
  wire [13:0] _GEN_13934 = 14'h366e == index ? 14'h6c : _GEN_13933;
  wire [13:0] _GEN_13935 = 14'h366f == index ? 14'h6c : _GEN_13934;
  wire [13:0] _GEN_13936 = 14'h3670 == index ? 14'h6c : _GEN_13935;
  wire [13:0] _GEN_13937 = 14'h3671 == index ? 14'h6c : _GEN_13936;
  wire [13:0] _GEN_13938 = 14'h3672 == index ? 14'h6c : _GEN_13937;
  wire [13:0] _GEN_13939 = 14'h3673 == index ? 14'h6c : _GEN_13938;
  wire [13:0] _GEN_13940 = 14'h3674 == index ? 14'h6c : _GEN_13939;
  wire [13:0] _GEN_13941 = 14'h3675 == index ? 14'h6c : _GEN_13940;
  wire [13:0] _GEN_13942 = 14'h3676 == index ? 14'h6c : _GEN_13941;
  wire [13:0] _GEN_13943 = 14'h3677 == index ? 14'h6c : _GEN_13942;
  wire [13:0] _GEN_13944 = 14'h3678 == index ? 14'h6c : _GEN_13943;
  wire [13:0] _GEN_13945 = 14'h3679 == index ? 14'h6c : _GEN_13944;
  wire [13:0] _GEN_13946 = 14'h367a == index ? 14'h6c : _GEN_13945;
  wire [13:0] _GEN_13947 = 14'h367b == index ? 14'h6c : _GEN_13946;
  wire [13:0] _GEN_13948 = 14'h367c == index ? 14'h6c : _GEN_13947;
  wire [13:0] _GEN_13949 = 14'h367d == index ? 14'h6c : _GEN_13948;
  wire [13:0] _GEN_13950 = 14'h367e == index ? 14'h6c : _GEN_13949;
  wire [13:0] _GEN_13951 = 14'h367f == index ? 14'h6c : _GEN_13950;
  wire [13:0] _GEN_13952 = 14'h3680 == index ? 14'h0 : _GEN_13951;
  wire [13:0] _GEN_13953 = 14'h3681 == index ? 14'h3680 : _GEN_13952;
  wire [13:0] _GEN_13954 = 14'h3682 == index ? 14'h1b01 : _GEN_13953;
  wire [13:0] _GEN_13955 = 14'h3683 == index ? 14'h1201 : _GEN_13954;
  wire [13:0] _GEN_13956 = 14'h3684 == index ? 14'hd81 : _GEN_13955;
  wire [13:0] _GEN_13957 = 14'h3685 == index ? 14'ha84 : _GEN_13956;
  wire [13:0] _GEN_13958 = 14'h3686 == index ? 14'h901 : _GEN_13957;
  wire [13:0] _GEN_13959 = 14'h3687 == index ? 14'h784 : _GEN_13958;
  wire [13:0] _GEN_13960 = 14'h3688 == index ? 14'h685 : _GEN_13959;
  wire [13:0] _GEN_13961 = 14'h3689 == index ? 14'h601 : _GEN_13960;
  wire [13:0] _GEN_13962 = 14'h368a == index ? 14'h509 : _GEN_13961;
  wire [13:0] _GEN_13963 = 14'h368b == index ? 14'h48a : _GEN_13962;
  wire [13:0] _GEN_13964 = 14'h368c == index ? 14'h481 : _GEN_13963;
  wire [13:0] _GEN_13965 = 14'h368d == index ? 14'h405 : _GEN_13964;
  wire [13:0] _GEN_13966 = 14'h368e == index ? 14'h38b : _GEN_13965;
  wire [13:0] _GEN_13967 = 14'h368f == index ? 14'h384 : _GEN_13966;
  wire [13:0] _GEN_13968 = 14'h3690 == index ? 14'h30d : _GEN_13967;
  wire [13:0] _GEN_13969 = 14'h3691 == index ? 14'h307 : _GEN_13968;
  wire [13:0] _GEN_13970 = 14'h3692 == index ? 14'h301 : _GEN_13969;
  wire [13:0] _GEN_13971 = 14'h3693 == index ? 14'h28e : _GEN_13970;
  wire [13:0] _GEN_13972 = 14'h3694 == index ? 14'h289 : _GEN_13971;
  wire [13:0] _GEN_13973 = 14'h3695 == index ? 14'h284 : _GEN_13972;
  wire [13:0] _GEN_13974 = 14'h3696 == index ? 14'h215 : _GEN_13973;
  wire [13:0] _GEN_13975 = 14'h3697 == index ? 14'h211 : _GEN_13974;
  wire [13:0] _GEN_13976 = 14'h3698 == index ? 14'h20d : _GEN_13975;
  wire [13:0] _GEN_13977 = 14'h3699 == index ? 14'h209 : _GEN_13976;
  wire [13:0] _GEN_13978 = 14'h369a == index ? 14'h205 : _GEN_13977;
  wire [13:0] _GEN_13979 = 14'h369b == index ? 14'h201 : _GEN_13978;
  wire [13:0] _GEN_13980 = 14'h369c == index ? 14'h199 : _GEN_13979;
  wire [13:0] _GEN_13981 = 14'h369d == index ? 14'h196 : _GEN_13980;
  wire [13:0] _GEN_13982 = 14'h369e == index ? 14'h193 : _GEN_13981;
  wire [13:0] _GEN_13983 = 14'h369f == index ? 14'h190 : _GEN_13982;
  wire [13:0] _GEN_13984 = 14'h36a0 == index ? 14'h18d : _GEN_13983;
  wire [13:0] _GEN_13985 = 14'h36a1 == index ? 14'h18a : _GEN_13984;
  wire [13:0] _GEN_13986 = 14'h36a2 == index ? 14'h187 : _GEN_13985;
  wire [13:0] _GEN_13987 = 14'h36a3 == index ? 14'h184 : _GEN_13986;
  wire [13:0] _GEN_13988 = 14'h36a4 == index ? 14'h181 : _GEN_13987;
  wire [13:0] _GEN_13989 = 14'h36a5 == index ? 14'h123 : _GEN_13988;
  wire [13:0] _GEN_13990 = 14'h36a6 == index ? 14'h121 : _GEN_13989;
  wire [13:0] _GEN_13991 = 14'h36a7 == index ? 14'h11f : _GEN_13990;
  wire [13:0] _GEN_13992 = 14'h36a8 == index ? 14'h11d : _GEN_13991;
  wire [13:0] _GEN_13993 = 14'h36a9 == index ? 14'h11b : _GEN_13992;
  wire [13:0] _GEN_13994 = 14'h36aa == index ? 14'h119 : _GEN_13993;
  wire [13:0] _GEN_13995 = 14'h36ab == index ? 14'h117 : _GEN_13994;
  wire [13:0] _GEN_13996 = 14'h36ac == index ? 14'h115 : _GEN_13995;
  wire [13:0] _GEN_13997 = 14'h36ad == index ? 14'h113 : _GEN_13996;
  wire [13:0] _GEN_13998 = 14'h36ae == index ? 14'h111 : _GEN_13997;
  wire [13:0] _GEN_13999 = 14'h36af == index ? 14'h10f : _GEN_13998;
  wire [13:0] _GEN_14000 = 14'h36b0 == index ? 14'h10d : _GEN_13999;
  wire [13:0] _GEN_14001 = 14'h36b1 == index ? 14'h10b : _GEN_14000;
  wire [13:0] _GEN_14002 = 14'h36b2 == index ? 14'h109 : _GEN_14001;
  wire [13:0] _GEN_14003 = 14'h36b3 == index ? 14'h107 : _GEN_14002;
  wire [13:0] _GEN_14004 = 14'h36b4 == index ? 14'h105 : _GEN_14003;
  wire [13:0] _GEN_14005 = 14'h36b5 == index ? 14'h103 : _GEN_14004;
  wire [13:0] _GEN_14006 = 14'h36b6 == index ? 14'h101 : _GEN_14005;
  wire [13:0] _GEN_14007 = 14'h36b7 == index ? 14'hb6 : _GEN_14006;
  wire [13:0] _GEN_14008 = 14'h36b8 == index ? 14'hb5 : _GEN_14007;
  wire [13:0] _GEN_14009 = 14'h36b9 == index ? 14'hb4 : _GEN_14008;
  wire [13:0] _GEN_14010 = 14'h36ba == index ? 14'hb3 : _GEN_14009;
  wire [13:0] _GEN_14011 = 14'h36bb == index ? 14'hb2 : _GEN_14010;
  wire [13:0] _GEN_14012 = 14'h36bc == index ? 14'hb1 : _GEN_14011;
  wire [13:0] _GEN_14013 = 14'h36bd == index ? 14'hb0 : _GEN_14012;
  wire [13:0] _GEN_14014 = 14'h36be == index ? 14'haf : _GEN_14013;
  wire [13:0] _GEN_14015 = 14'h36bf == index ? 14'hae : _GEN_14014;
  wire [13:0] _GEN_14016 = 14'h36c0 == index ? 14'had : _GEN_14015;
  wire [13:0] _GEN_14017 = 14'h36c1 == index ? 14'hac : _GEN_14016;
  wire [13:0] _GEN_14018 = 14'h36c2 == index ? 14'hab : _GEN_14017;
  wire [13:0] _GEN_14019 = 14'h36c3 == index ? 14'haa : _GEN_14018;
  wire [13:0] _GEN_14020 = 14'h36c4 == index ? 14'ha9 : _GEN_14019;
  wire [13:0] _GEN_14021 = 14'h36c5 == index ? 14'ha8 : _GEN_14020;
  wire [13:0] _GEN_14022 = 14'h36c6 == index ? 14'ha7 : _GEN_14021;
  wire [13:0] _GEN_14023 = 14'h36c7 == index ? 14'ha6 : _GEN_14022;
  wire [13:0] _GEN_14024 = 14'h36c8 == index ? 14'ha5 : _GEN_14023;
  wire [13:0] _GEN_14025 = 14'h36c9 == index ? 14'ha4 : _GEN_14024;
  wire [13:0] _GEN_14026 = 14'h36ca == index ? 14'ha3 : _GEN_14025;
  wire [13:0] _GEN_14027 = 14'h36cb == index ? 14'ha2 : _GEN_14026;
  wire [13:0] _GEN_14028 = 14'h36cc == index ? 14'ha1 : _GEN_14027;
  wire [13:0] _GEN_14029 = 14'h36cd == index ? 14'ha0 : _GEN_14028;
  wire [13:0] _GEN_14030 = 14'h36ce == index ? 14'h9f : _GEN_14029;
  wire [13:0] _GEN_14031 = 14'h36cf == index ? 14'h9e : _GEN_14030;
  wire [13:0] _GEN_14032 = 14'h36d0 == index ? 14'h9d : _GEN_14031;
  wire [13:0] _GEN_14033 = 14'h36d1 == index ? 14'h9c : _GEN_14032;
  wire [13:0] _GEN_14034 = 14'h36d2 == index ? 14'h9b : _GEN_14033;
  wire [13:0] _GEN_14035 = 14'h36d3 == index ? 14'h9a : _GEN_14034;
  wire [13:0] _GEN_14036 = 14'h36d4 == index ? 14'h99 : _GEN_14035;
  wire [13:0] _GEN_14037 = 14'h36d5 == index ? 14'h98 : _GEN_14036;
  wire [13:0] _GEN_14038 = 14'h36d6 == index ? 14'h97 : _GEN_14037;
  wire [13:0] _GEN_14039 = 14'h36d7 == index ? 14'h96 : _GEN_14038;
  wire [13:0] _GEN_14040 = 14'h36d8 == index ? 14'h95 : _GEN_14039;
  wire [13:0] _GEN_14041 = 14'h36d9 == index ? 14'h94 : _GEN_14040;
  wire [13:0] _GEN_14042 = 14'h36da == index ? 14'h93 : _GEN_14041;
  wire [13:0] _GEN_14043 = 14'h36db == index ? 14'h92 : _GEN_14042;
  wire [13:0] _GEN_14044 = 14'h36dc == index ? 14'h91 : _GEN_14043;
  wire [13:0] _GEN_14045 = 14'h36dd == index ? 14'h90 : _GEN_14044;
  wire [13:0] _GEN_14046 = 14'h36de == index ? 14'h8f : _GEN_14045;
  wire [13:0] _GEN_14047 = 14'h36df == index ? 14'h8e : _GEN_14046;
  wire [13:0] _GEN_14048 = 14'h36e0 == index ? 14'h8d : _GEN_14047;
  wire [13:0] _GEN_14049 = 14'h36e1 == index ? 14'h8c : _GEN_14048;
  wire [13:0] _GEN_14050 = 14'h36e2 == index ? 14'h8b : _GEN_14049;
  wire [13:0] _GEN_14051 = 14'h36e3 == index ? 14'h8a : _GEN_14050;
  wire [13:0] _GEN_14052 = 14'h36e4 == index ? 14'h89 : _GEN_14051;
  wire [13:0] _GEN_14053 = 14'h36e5 == index ? 14'h88 : _GEN_14052;
  wire [13:0] _GEN_14054 = 14'h36e6 == index ? 14'h87 : _GEN_14053;
  wire [13:0] _GEN_14055 = 14'h36e7 == index ? 14'h86 : _GEN_14054;
  wire [13:0] _GEN_14056 = 14'h36e8 == index ? 14'h85 : _GEN_14055;
  wire [13:0] _GEN_14057 = 14'h36e9 == index ? 14'h84 : _GEN_14056;
  wire [13:0] _GEN_14058 = 14'h36ea == index ? 14'h83 : _GEN_14057;
  wire [13:0] _GEN_14059 = 14'h36eb == index ? 14'h82 : _GEN_14058;
  wire [13:0] _GEN_14060 = 14'h36ec == index ? 14'h81 : _GEN_14059;
  wire [13:0] _GEN_14061 = 14'h36ed == index ? 14'h80 : _GEN_14060;
  wire [13:0] _GEN_14062 = 14'h36ee == index ? 14'h6d : _GEN_14061;
  wire [13:0] _GEN_14063 = 14'h36ef == index ? 14'h6d : _GEN_14062;
  wire [13:0] _GEN_14064 = 14'h36f0 == index ? 14'h6d : _GEN_14063;
  wire [13:0] _GEN_14065 = 14'h36f1 == index ? 14'h6d : _GEN_14064;
  wire [13:0] _GEN_14066 = 14'h36f2 == index ? 14'h6d : _GEN_14065;
  wire [13:0] _GEN_14067 = 14'h36f3 == index ? 14'h6d : _GEN_14066;
  wire [13:0] _GEN_14068 = 14'h36f4 == index ? 14'h6d : _GEN_14067;
  wire [13:0] _GEN_14069 = 14'h36f5 == index ? 14'h6d : _GEN_14068;
  wire [13:0] _GEN_14070 = 14'h36f6 == index ? 14'h6d : _GEN_14069;
  wire [13:0] _GEN_14071 = 14'h36f7 == index ? 14'h6d : _GEN_14070;
  wire [13:0] _GEN_14072 = 14'h36f8 == index ? 14'h6d : _GEN_14071;
  wire [13:0] _GEN_14073 = 14'h36f9 == index ? 14'h6d : _GEN_14072;
  wire [13:0] _GEN_14074 = 14'h36fa == index ? 14'h6d : _GEN_14073;
  wire [13:0] _GEN_14075 = 14'h36fb == index ? 14'h6d : _GEN_14074;
  wire [13:0] _GEN_14076 = 14'h36fc == index ? 14'h6d : _GEN_14075;
  wire [13:0] _GEN_14077 = 14'h36fd == index ? 14'h6d : _GEN_14076;
  wire [13:0] _GEN_14078 = 14'h36fe == index ? 14'h6d : _GEN_14077;
  wire [13:0] _GEN_14079 = 14'h36ff == index ? 14'h6d : _GEN_14078;
  wire [13:0] _GEN_14080 = 14'h3700 == index ? 14'h0 : _GEN_14079;
  wire [13:0] _GEN_14081 = 14'h3701 == index ? 14'h3700 : _GEN_14080;
  wire [13:0] _GEN_14082 = 14'h3702 == index ? 14'h1b80 : _GEN_14081;
  wire [13:0] _GEN_14083 = 14'h3703 == index ? 14'h1202 : _GEN_14082;
  wire [13:0] _GEN_14084 = 14'h3704 == index ? 14'hd82 : _GEN_14083;
  wire [13:0] _GEN_14085 = 14'h3705 == index ? 14'hb00 : _GEN_14084;
  wire [13:0] _GEN_14086 = 14'h3706 == index ? 14'h902 : _GEN_14085;
  wire [13:0] _GEN_14087 = 14'h3707 == index ? 14'h785 : _GEN_14086;
  wire [13:0] _GEN_14088 = 14'h3708 == index ? 14'h686 : _GEN_14087;
  wire [13:0] _GEN_14089 = 14'h3709 == index ? 14'h602 : _GEN_14088;
  wire [13:0] _GEN_14090 = 14'h370a == index ? 14'h580 : _GEN_14089;
  wire [13:0] _GEN_14091 = 14'h370b == index ? 14'h500 : _GEN_14090;
  wire [13:0] _GEN_14092 = 14'h370c == index ? 14'h482 : _GEN_14091;
  wire [13:0] _GEN_14093 = 14'h370d == index ? 14'h406 : _GEN_14092;
  wire [13:0] _GEN_14094 = 14'h370e == index ? 14'h38c : _GEN_14093;
  wire [13:0] _GEN_14095 = 14'h370f == index ? 14'h385 : _GEN_14094;
  wire [13:0] _GEN_14096 = 14'h3710 == index ? 14'h30e : _GEN_14095;
  wire [13:0] _GEN_14097 = 14'h3711 == index ? 14'h308 : _GEN_14096;
  wire [13:0] _GEN_14098 = 14'h3712 == index ? 14'h302 : _GEN_14097;
  wire [13:0] _GEN_14099 = 14'h3713 == index ? 14'h28f : _GEN_14098;
  wire [13:0] _GEN_14100 = 14'h3714 == index ? 14'h28a : _GEN_14099;
  wire [13:0] _GEN_14101 = 14'h3715 == index ? 14'h285 : _GEN_14100;
  wire [13:0] _GEN_14102 = 14'h3716 == index ? 14'h280 : _GEN_14101;
  wire [13:0] _GEN_14103 = 14'h3717 == index ? 14'h212 : _GEN_14102;
  wire [13:0] _GEN_14104 = 14'h3718 == index ? 14'h20e : _GEN_14103;
  wire [13:0] _GEN_14105 = 14'h3719 == index ? 14'h20a : _GEN_14104;
  wire [13:0] _GEN_14106 = 14'h371a == index ? 14'h206 : _GEN_14105;
  wire [13:0] _GEN_14107 = 14'h371b == index ? 14'h202 : _GEN_14106;
  wire [13:0] _GEN_14108 = 14'h371c == index ? 14'h19a : _GEN_14107;
  wire [13:0] _GEN_14109 = 14'h371d == index ? 14'h197 : _GEN_14108;
  wire [13:0] _GEN_14110 = 14'h371e == index ? 14'h194 : _GEN_14109;
  wire [13:0] _GEN_14111 = 14'h371f == index ? 14'h191 : _GEN_14110;
  wire [13:0] _GEN_14112 = 14'h3720 == index ? 14'h18e : _GEN_14111;
  wire [13:0] _GEN_14113 = 14'h3721 == index ? 14'h18b : _GEN_14112;
  wire [13:0] _GEN_14114 = 14'h3722 == index ? 14'h188 : _GEN_14113;
  wire [13:0] _GEN_14115 = 14'h3723 == index ? 14'h185 : _GEN_14114;
  wire [13:0] _GEN_14116 = 14'h3724 == index ? 14'h182 : _GEN_14115;
  wire [13:0] _GEN_14117 = 14'h3725 == index ? 14'h124 : _GEN_14116;
  wire [13:0] _GEN_14118 = 14'h3726 == index ? 14'h122 : _GEN_14117;
  wire [13:0] _GEN_14119 = 14'h3727 == index ? 14'h120 : _GEN_14118;
  wire [13:0] _GEN_14120 = 14'h3728 == index ? 14'h11e : _GEN_14119;
  wire [13:0] _GEN_14121 = 14'h3729 == index ? 14'h11c : _GEN_14120;
  wire [13:0] _GEN_14122 = 14'h372a == index ? 14'h11a : _GEN_14121;
  wire [13:0] _GEN_14123 = 14'h372b == index ? 14'h118 : _GEN_14122;
  wire [13:0] _GEN_14124 = 14'h372c == index ? 14'h116 : _GEN_14123;
  wire [13:0] _GEN_14125 = 14'h372d == index ? 14'h114 : _GEN_14124;
  wire [13:0] _GEN_14126 = 14'h372e == index ? 14'h112 : _GEN_14125;
  wire [13:0] _GEN_14127 = 14'h372f == index ? 14'h110 : _GEN_14126;
  wire [13:0] _GEN_14128 = 14'h3730 == index ? 14'h10e : _GEN_14127;
  wire [13:0] _GEN_14129 = 14'h3731 == index ? 14'h10c : _GEN_14128;
  wire [13:0] _GEN_14130 = 14'h3732 == index ? 14'h10a : _GEN_14129;
  wire [13:0] _GEN_14131 = 14'h3733 == index ? 14'h108 : _GEN_14130;
  wire [13:0] _GEN_14132 = 14'h3734 == index ? 14'h106 : _GEN_14131;
  wire [13:0] _GEN_14133 = 14'h3735 == index ? 14'h104 : _GEN_14132;
  wire [13:0] _GEN_14134 = 14'h3736 == index ? 14'h102 : _GEN_14133;
  wire [13:0] _GEN_14135 = 14'h3737 == index ? 14'h100 : _GEN_14134;
  wire [13:0] _GEN_14136 = 14'h3738 == index ? 14'hb6 : _GEN_14135;
  wire [13:0] _GEN_14137 = 14'h3739 == index ? 14'hb5 : _GEN_14136;
  wire [13:0] _GEN_14138 = 14'h373a == index ? 14'hb4 : _GEN_14137;
  wire [13:0] _GEN_14139 = 14'h373b == index ? 14'hb3 : _GEN_14138;
  wire [13:0] _GEN_14140 = 14'h373c == index ? 14'hb2 : _GEN_14139;
  wire [13:0] _GEN_14141 = 14'h373d == index ? 14'hb1 : _GEN_14140;
  wire [13:0] _GEN_14142 = 14'h373e == index ? 14'hb0 : _GEN_14141;
  wire [13:0] _GEN_14143 = 14'h373f == index ? 14'haf : _GEN_14142;
  wire [13:0] _GEN_14144 = 14'h3740 == index ? 14'hae : _GEN_14143;
  wire [13:0] _GEN_14145 = 14'h3741 == index ? 14'had : _GEN_14144;
  wire [13:0] _GEN_14146 = 14'h3742 == index ? 14'hac : _GEN_14145;
  wire [13:0] _GEN_14147 = 14'h3743 == index ? 14'hab : _GEN_14146;
  wire [13:0] _GEN_14148 = 14'h3744 == index ? 14'haa : _GEN_14147;
  wire [13:0] _GEN_14149 = 14'h3745 == index ? 14'ha9 : _GEN_14148;
  wire [13:0] _GEN_14150 = 14'h3746 == index ? 14'ha8 : _GEN_14149;
  wire [13:0] _GEN_14151 = 14'h3747 == index ? 14'ha7 : _GEN_14150;
  wire [13:0] _GEN_14152 = 14'h3748 == index ? 14'ha6 : _GEN_14151;
  wire [13:0] _GEN_14153 = 14'h3749 == index ? 14'ha5 : _GEN_14152;
  wire [13:0] _GEN_14154 = 14'h374a == index ? 14'ha4 : _GEN_14153;
  wire [13:0] _GEN_14155 = 14'h374b == index ? 14'ha3 : _GEN_14154;
  wire [13:0] _GEN_14156 = 14'h374c == index ? 14'ha2 : _GEN_14155;
  wire [13:0] _GEN_14157 = 14'h374d == index ? 14'ha1 : _GEN_14156;
  wire [13:0] _GEN_14158 = 14'h374e == index ? 14'ha0 : _GEN_14157;
  wire [13:0] _GEN_14159 = 14'h374f == index ? 14'h9f : _GEN_14158;
  wire [13:0] _GEN_14160 = 14'h3750 == index ? 14'h9e : _GEN_14159;
  wire [13:0] _GEN_14161 = 14'h3751 == index ? 14'h9d : _GEN_14160;
  wire [13:0] _GEN_14162 = 14'h3752 == index ? 14'h9c : _GEN_14161;
  wire [13:0] _GEN_14163 = 14'h3753 == index ? 14'h9b : _GEN_14162;
  wire [13:0] _GEN_14164 = 14'h3754 == index ? 14'h9a : _GEN_14163;
  wire [13:0] _GEN_14165 = 14'h3755 == index ? 14'h99 : _GEN_14164;
  wire [13:0] _GEN_14166 = 14'h3756 == index ? 14'h98 : _GEN_14165;
  wire [13:0] _GEN_14167 = 14'h3757 == index ? 14'h97 : _GEN_14166;
  wire [13:0] _GEN_14168 = 14'h3758 == index ? 14'h96 : _GEN_14167;
  wire [13:0] _GEN_14169 = 14'h3759 == index ? 14'h95 : _GEN_14168;
  wire [13:0] _GEN_14170 = 14'h375a == index ? 14'h94 : _GEN_14169;
  wire [13:0] _GEN_14171 = 14'h375b == index ? 14'h93 : _GEN_14170;
  wire [13:0] _GEN_14172 = 14'h375c == index ? 14'h92 : _GEN_14171;
  wire [13:0] _GEN_14173 = 14'h375d == index ? 14'h91 : _GEN_14172;
  wire [13:0] _GEN_14174 = 14'h375e == index ? 14'h90 : _GEN_14173;
  wire [13:0] _GEN_14175 = 14'h375f == index ? 14'h8f : _GEN_14174;
  wire [13:0] _GEN_14176 = 14'h3760 == index ? 14'h8e : _GEN_14175;
  wire [13:0] _GEN_14177 = 14'h3761 == index ? 14'h8d : _GEN_14176;
  wire [13:0] _GEN_14178 = 14'h3762 == index ? 14'h8c : _GEN_14177;
  wire [13:0] _GEN_14179 = 14'h3763 == index ? 14'h8b : _GEN_14178;
  wire [13:0] _GEN_14180 = 14'h3764 == index ? 14'h8a : _GEN_14179;
  wire [13:0] _GEN_14181 = 14'h3765 == index ? 14'h89 : _GEN_14180;
  wire [13:0] _GEN_14182 = 14'h3766 == index ? 14'h88 : _GEN_14181;
  wire [13:0] _GEN_14183 = 14'h3767 == index ? 14'h87 : _GEN_14182;
  wire [13:0] _GEN_14184 = 14'h3768 == index ? 14'h86 : _GEN_14183;
  wire [13:0] _GEN_14185 = 14'h3769 == index ? 14'h85 : _GEN_14184;
  wire [13:0] _GEN_14186 = 14'h376a == index ? 14'h84 : _GEN_14185;
  wire [13:0] _GEN_14187 = 14'h376b == index ? 14'h83 : _GEN_14186;
  wire [13:0] _GEN_14188 = 14'h376c == index ? 14'h82 : _GEN_14187;
  wire [13:0] _GEN_14189 = 14'h376d == index ? 14'h81 : _GEN_14188;
  wire [13:0] _GEN_14190 = 14'h376e == index ? 14'h80 : _GEN_14189;
  wire [13:0] _GEN_14191 = 14'h376f == index ? 14'h6e : _GEN_14190;
  wire [13:0] _GEN_14192 = 14'h3770 == index ? 14'h6e : _GEN_14191;
  wire [13:0] _GEN_14193 = 14'h3771 == index ? 14'h6e : _GEN_14192;
  wire [13:0] _GEN_14194 = 14'h3772 == index ? 14'h6e : _GEN_14193;
  wire [13:0] _GEN_14195 = 14'h3773 == index ? 14'h6e : _GEN_14194;
  wire [13:0] _GEN_14196 = 14'h3774 == index ? 14'h6e : _GEN_14195;
  wire [13:0] _GEN_14197 = 14'h3775 == index ? 14'h6e : _GEN_14196;
  wire [13:0] _GEN_14198 = 14'h3776 == index ? 14'h6e : _GEN_14197;
  wire [13:0] _GEN_14199 = 14'h3777 == index ? 14'h6e : _GEN_14198;
  wire [13:0] _GEN_14200 = 14'h3778 == index ? 14'h6e : _GEN_14199;
  wire [13:0] _GEN_14201 = 14'h3779 == index ? 14'h6e : _GEN_14200;
  wire [13:0] _GEN_14202 = 14'h377a == index ? 14'h6e : _GEN_14201;
  wire [13:0] _GEN_14203 = 14'h377b == index ? 14'h6e : _GEN_14202;
  wire [13:0] _GEN_14204 = 14'h377c == index ? 14'h6e : _GEN_14203;
  wire [13:0] _GEN_14205 = 14'h377d == index ? 14'h6e : _GEN_14204;
  wire [13:0] _GEN_14206 = 14'h377e == index ? 14'h6e : _GEN_14205;
  wire [13:0] _GEN_14207 = 14'h377f == index ? 14'h6e : _GEN_14206;
  wire [13:0] _GEN_14208 = 14'h3780 == index ? 14'h0 : _GEN_14207;
  wire [13:0] _GEN_14209 = 14'h3781 == index ? 14'h3780 : _GEN_14208;
  wire [13:0] _GEN_14210 = 14'h3782 == index ? 14'h1b81 : _GEN_14209;
  wire [13:0] _GEN_14211 = 14'h3783 == index ? 14'h1280 : _GEN_14210;
  wire [13:0] _GEN_14212 = 14'h3784 == index ? 14'hd83 : _GEN_14211;
  wire [13:0] _GEN_14213 = 14'h3785 == index ? 14'hb01 : _GEN_14212;
  wire [13:0] _GEN_14214 = 14'h3786 == index ? 14'h903 : _GEN_14213;
  wire [13:0] _GEN_14215 = 14'h3787 == index ? 14'h786 : _GEN_14214;
  wire [13:0] _GEN_14216 = 14'h3788 == index ? 14'h687 : _GEN_14215;
  wire [13:0] _GEN_14217 = 14'h3789 == index ? 14'h603 : _GEN_14216;
  wire [13:0] _GEN_14218 = 14'h378a == index ? 14'h581 : _GEN_14217;
  wire [13:0] _GEN_14219 = 14'h378b == index ? 14'h501 : _GEN_14218;
  wire [13:0] _GEN_14220 = 14'h378c == index ? 14'h483 : _GEN_14219;
  wire [13:0] _GEN_14221 = 14'h378d == index ? 14'h407 : _GEN_14220;
  wire [13:0] _GEN_14222 = 14'h378e == index ? 14'h38d : _GEN_14221;
  wire [13:0] _GEN_14223 = 14'h378f == index ? 14'h386 : _GEN_14222;
  wire [13:0] _GEN_14224 = 14'h3790 == index ? 14'h30f : _GEN_14223;
  wire [13:0] _GEN_14225 = 14'h3791 == index ? 14'h309 : _GEN_14224;
  wire [13:0] _GEN_14226 = 14'h3792 == index ? 14'h303 : _GEN_14225;
  wire [13:0] _GEN_14227 = 14'h3793 == index ? 14'h290 : _GEN_14226;
  wire [13:0] _GEN_14228 = 14'h3794 == index ? 14'h28b : _GEN_14227;
  wire [13:0] _GEN_14229 = 14'h3795 == index ? 14'h286 : _GEN_14228;
  wire [13:0] _GEN_14230 = 14'h3796 == index ? 14'h281 : _GEN_14229;
  wire [13:0] _GEN_14231 = 14'h3797 == index ? 14'h213 : _GEN_14230;
  wire [13:0] _GEN_14232 = 14'h3798 == index ? 14'h20f : _GEN_14231;
  wire [13:0] _GEN_14233 = 14'h3799 == index ? 14'h20b : _GEN_14232;
  wire [13:0] _GEN_14234 = 14'h379a == index ? 14'h207 : _GEN_14233;
  wire [13:0] _GEN_14235 = 14'h379b == index ? 14'h203 : _GEN_14234;
  wire [13:0] _GEN_14236 = 14'h379c == index ? 14'h19b : _GEN_14235;
  wire [13:0] _GEN_14237 = 14'h379d == index ? 14'h198 : _GEN_14236;
  wire [13:0] _GEN_14238 = 14'h379e == index ? 14'h195 : _GEN_14237;
  wire [13:0] _GEN_14239 = 14'h379f == index ? 14'h192 : _GEN_14238;
  wire [13:0] _GEN_14240 = 14'h37a0 == index ? 14'h18f : _GEN_14239;
  wire [13:0] _GEN_14241 = 14'h37a1 == index ? 14'h18c : _GEN_14240;
  wire [13:0] _GEN_14242 = 14'h37a2 == index ? 14'h189 : _GEN_14241;
  wire [13:0] _GEN_14243 = 14'h37a3 == index ? 14'h186 : _GEN_14242;
  wire [13:0] _GEN_14244 = 14'h37a4 == index ? 14'h183 : _GEN_14243;
  wire [13:0] _GEN_14245 = 14'h37a5 == index ? 14'h180 : _GEN_14244;
  wire [13:0] _GEN_14246 = 14'h37a6 == index ? 14'h123 : _GEN_14245;
  wire [13:0] _GEN_14247 = 14'h37a7 == index ? 14'h121 : _GEN_14246;
  wire [13:0] _GEN_14248 = 14'h37a8 == index ? 14'h11f : _GEN_14247;
  wire [13:0] _GEN_14249 = 14'h37a9 == index ? 14'h11d : _GEN_14248;
  wire [13:0] _GEN_14250 = 14'h37aa == index ? 14'h11b : _GEN_14249;
  wire [13:0] _GEN_14251 = 14'h37ab == index ? 14'h119 : _GEN_14250;
  wire [13:0] _GEN_14252 = 14'h37ac == index ? 14'h117 : _GEN_14251;
  wire [13:0] _GEN_14253 = 14'h37ad == index ? 14'h115 : _GEN_14252;
  wire [13:0] _GEN_14254 = 14'h37ae == index ? 14'h113 : _GEN_14253;
  wire [13:0] _GEN_14255 = 14'h37af == index ? 14'h111 : _GEN_14254;
  wire [13:0] _GEN_14256 = 14'h37b0 == index ? 14'h10f : _GEN_14255;
  wire [13:0] _GEN_14257 = 14'h37b1 == index ? 14'h10d : _GEN_14256;
  wire [13:0] _GEN_14258 = 14'h37b2 == index ? 14'h10b : _GEN_14257;
  wire [13:0] _GEN_14259 = 14'h37b3 == index ? 14'h109 : _GEN_14258;
  wire [13:0] _GEN_14260 = 14'h37b4 == index ? 14'h107 : _GEN_14259;
  wire [13:0] _GEN_14261 = 14'h37b5 == index ? 14'h105 : _GEN_14260;
  wire [13:0] _GEN_14262 = 14'h37b6 == index ? 14'h103 : _GEN_14261;
  wire [13:0] _GEN_14263 = 14'h37b7 == index ? 14'h101 : _GEN_14262;
  wire [13:0] _GEN_14264 = 14'h37b8 == index ? 14'hb7 : _GEN_14263;
  wire [13:0] _GEN_14265 = 14'h37b9 == index ? 14'hb6 : _GEN_14264;
  wire [13:0] _GEN_14266 = 14'h37ba == index ? 14'hb5 : _GEN_14265;
  wire [13:0] _GEN_14267 = 14'h37bb == index ? 14'hb4 : _GEN_14266;
  wire [13:0] _GEN_14268 = 14'h37bc == index ? 14'hb3 : _GEN_14267;
  wire [13:0] _GEN_14269 = 14'h37bd == index ? 14'hb2 : _GEN_14268;
  wire [13:0] _GEN_14270 = 14'h37be == index ? 14'hb1 : _GEN_14269;
  wire [13:0] _GEN_14271 = 14'h37bf == index ? 14'hb0 : _GEN_14270;
  wire [13:0] _GEN_14272 = 14'h37c0 == index ? 14'haf : _GEN_14271;
  wire [13:0] _GEN_14273 = 14'h37c1 == index ? 14'hae : _GEN_14272;
  wire [13:0] _GEN_14274 = 14'h37c2 == index ? 14'had : _GEN_14273;
  wire [13:0] _GEN_14275 = 14'h37c3 == index ? 14'hac : _GEN_14274;
  wire [13:0] _GEN_14276 = 14'h37c4 == index ? 14'hab : _GEN_14275;
  wire [13:0] _GEN_14277 = 14'h37c5 == index ? 14'haa : _GEN_14276;
  wire [13:0] _GEN_14278 = 14'h37c6 == index ? 14'ha9 : _GEN_14277;
  wire [13:0] _GEN_14279 = 14'h37c7 == index ? 14'ha8 : _GEN_14278;
  wire [13:0] _GEN_14280 = 14'h37c8 == index ? 14'ha7 : _GEN_14279;
  wire [13:0] _GEN_14281 = 14'h37c9 == index ? 14'ha6 : _GEN_14280;
  wire [13:0] _GEN_14282 = 14'h37ca == index ? 14'ha5 : _GEN_14281;
  wire [13:0] _GEN_14283 = 14'h37cb == index ? 14'ha4 : _GEN_14282;
  wire [13:0] _GEN_14284 = 14'h37cc == index ? 14'ha3 : _GEN_14283;
  wire [13:0] _GEN_14285 = 14'h37cd == index ? 14'ha2 : _GEN_14284;
  wire [13:0] _GEN_14286 = 14'h37ce == index ? 14'ha1 : _GEN_14285;
  wire [13:0] _GEN_14287 = 14'h37cf == index ? 14'ha0 : _GEN_14286;
  wire [13:0] _GEN_14288 = 14'h37d0 == index ? 14'h9f : _GEN_14287;
  wire [13:0] _GEN_14289 = 14'h37d1 == index ? 14'h9e : _GEN_14288;
  wire [13:0] _GEN_14290 = 14'h37d2 == index ? 14'h9d : _GEN_14289;
  wire [13:0] _GEN_14291 = 14'h37d3 == index ? 14'h9c : _GEN_14290;
  wire [13:0] _GEN_14292 = 14'h37d4 == index ? 14'h9b : _GEN_14291;
  wire [13:0] _GEN_14293 = 14'h37d5 == index ? 14'h9a : _GEN_14292;
  wire [13:0] _GEN_14294 = 14'h37d6 == index ? 14'h99 : _GEN_14293;
  wire [13:0] _GEN_14295 = 14'h37d7 == index ? 14'h98 : _GEN_14294;
  wire [13:0] _GEN_14296 = 14'h37d8 == index ? 14'h97 : _GEN_14295;
  wire [13:0] _GEN_14297 = 14'h37d9 == index ? 14'h96 : _GEN_14296;
  wire [13:0] _GEN_14298 = 14'h37da == index ? 14'h95 : _GEN_14297;
  wire [13:0] _GEN_14299 = 14'h37db == index ? 14'h94 : _GEN_14298;
  wire [13:0] _GEN_14300 = 14'h37dc == index ? 14'h93 : _GEN_14299;
  wire [13:0] _GEN_14301 = 14'h37dd == index ? 14'h92 : _GEN_14300;
  wire [13:0] _GEN_14302 = 14'h37de == index ? 14'h91 : _GEN_14301;
  wire [13:0] _GEN_14303 = 14'h37df == index ? 14'h90 : _GEN_14302;
  wire [13:0] _GEN_14304 = 14'h37e0 == index ? 14'h8f : _GEN_14303;
  wire [13:0] _GEN_14305 = 14'h37e1 == index ? 14'h8e : _GEN_14304;
  wire [13:0] _GEN_14306 = 14'h37e2 == index ? 14'h8d : _GEN_14305;
  wire [13:0] _GEN_14307 = 14'h37e3 == index ? 14'h8c : _GEN_14306;
  wire [13:0] _GEN_14308 = 14'h37e4 == index ? 14'h8b : _GEN_14307;
  wire [13:0] _GEN_14309 = 14'h37e5 == index ? 14'h8a : _GEN_14308;
  wire [13:0] _GEN_14310 = 14'h37e6 == index ? 14'h89 : _GEN_14309;
  wire [13:0] _GEN_14311 = 14'h37e7 == index ? 14'h88 : _GEN_14310;
  wire [13:0] _GEN_14312 = 14'h37e8 == index ? 14'h87 : _GEN_14311;
  wire [13:0] _GEN_14313 = 14'h37e9 == index ? 14'h86 : _GEN_14312;
  wire [13:0] _GEN_14314 = 14'h37ea == index ? 14'h85 : _GEN_14313;
  wire [13:0] _GEN_14315 = 14'h37eb == index ? 14'h84 : _GEN_14314;
  wire [13:0] _GEN_14316 = 14'h37ec == index ? 14'h83 : _GEN_14315;
  wire [13:0] _GEN_14317 = 14'h37ed == index ? 14'h82 : _GEN_14316;
  wire [13:0] _GEN_14318 = 14'h37ee == index ? 14'h81 : _GEN_14317;
  wire [13:0] _GEN_14319 = 14'h37ef == index ? 14'h80 : _GEN_14318;
  wire [13:0] _GEN_14320 = 14'h37f0 == index ? 14'h6f : _GEN_14319;
  wire [13:0] _GEN_14321 = 14'h37f1 == index ? 14'h6f : _GEN_14320;
  wire [13:0] _GEN_14322 = 14'h37f2 == index ? 14'h6f : _GEN_14321;
  wire [13:0] _GEN_14323 = 14'h37f3 == index ? 14'h6f : _GEN_14322;
  wire [13:0] _GEN_14324 = 14'h37f4 == index ? 14'h6f : _GEN_14323;
  wire [13:0] _GEN_14325 = 14'h37f5 == index ? 14'h6f : _GEN_14324;
  wire [13:0] _GEN_14326 = 14'h37f6 == index ? 14'h6f : _GEN_14325;
  wire [13:0] _GEN_14327 = 14'h37f7 == index ? 14'h6f : _GEN_14326;
  wire [13:0] _GEN_14328 = 14'h37f8 == index ? 14'h6f : _GEN_14327;
  wire [13:0] _GEN_14329 = 14'h37f9 == index ? 14'h6f : _GEN_14328;
  wire [13:0] _GEN_14330 = 14'h37fa == index ? 14'h6f : _GEN_14329;
  wire [13:0] _GEN_14331 = 14'h37fb == index ? 14'h6f : _GEN_14330;
  wire [13:0] _GEN_14332 = 14'h37fc == index ? 14'h6f : _GEN_14331;
  wire [13:0] _GEN_14333 = 14'h37fd == index ? 14'h6f : _GEN_14332;
  wire [13:0] _GEN_14334 = 14'h37fe == index ? 14'h6f : _GEN_14333;
  wire [13:0] _GEN_14335 = 14'h37ff == index ? 14'h6f : _GEN_14334;
  wire [13:0] _GEN_14336 = 14'h3800 == index ? 14'h0 : _GEN_14335;
  wire [13:0] _GEN_14337 = 14'h3801 == index ? 14'h3800 : _GEN_14336;
  wire [13:0] _GEN_14338 = 14'h3802 == index ? 14'h1c00 : _GEN_14337;
  wire [13:0] _GEN_14339 = 14'h3803 == index ? 14'h1281 : _GEN_14338;
  wire [13:0] _GEN_14340 = 14'h3804 == index ? 14'he00 : _GEN_14339;
  wire [13:0] _GEN_14341 = 14'h3805 == index ? 14'hb02 : _GEN_14340;
  wire [13:0] _GEN_14342 = 14'h3806 == index ? 14'h904 : _GEN_14341;
  wire [13:0] _GEN_14343 = 14'h3807 == index ? 14'h800 : _GEN_14342;
  wire [13:0] _GEN_14344 = 14'h3808 == index ? 14'h700 : _GEN_14343;
  wire [13:0] _GEN_14345 = 14'h3809 == index ? 14'h604 : _GEN_14344;
  wire [13:0] _GEN_14346 = 14'h380a == index ? 14'h582 : _GEN_14345;
  wire [13:0] _GEN_14347 = 14'h380b == index ? 14'h502 : _GEN_14346;
  wire [13:0] _GEN_14348 = 14'h380c == index ? 14'h484 : _GEN_14347;
  wire [13:0] _GEN_14349 = 14'h380d == index ? 14'h408 : _GEN_14348;
  wire [13:0] _GEN_14350 = 14'h380e == index ? 14'h400 : _GEN_14349;
  wire [13:0] _GEN_14351 = 14'h380f == index ? 14'h387 : _GEN_14350;
  wire [13:0] _GEN_14352 = 14'h3810 == index ? 14'h380 : _GEN_14351;
  wire [13:0] _GEN_14353 = 14'h3811 == index ? 14'h30a : _GEN_14352;
  wire [13:0] _GEN_14354 = 14'h3812 == index ? 14'h304 : _GEN_14353;
  wire [13:0] _GEN_14355 = 14'h3813 == index ? 14'h291 : _GEN_14354;
  wire [13:0] _GEN_14356 = 14'h3814 == index ? 14'h28c : _GEN_14355;
  wire [13:0] _GEN_14357 = 14'h3815 == index ? 14'h287 : _GEN_14356;
  wire [13:0] _GEN_14358 = 14'h3816 == index ? 14'h282 : _GEN_14357;
  wire [13:0] _GEN_14359 = 14'h3817 == index ? 14'h214 : _GEN_14358;
  wire [13:0] _GEN_14360 = 14'h3818 == index ? 14'h210 : _GEN_14359;
  wire [13:0] _GEN_14361 = 14'h3819 == index ? 14'h20c : _GEN_14360;
  wire [13:0] _GEN_14362 = 14'h381a == index ? 14'h208 : _GEN_14361;
  wire [13:0] _GEN_14363 = 14'h381b == index ? 14'h204 : _GEN_14362;
  wire [13:0] _GEN_14364 = 14'h381c == index ? 14'h200 : _GEN_14363;
  wire [13:0] _GEN_14365 = 14'h381d == index ? 14'h199 : _GEN_14364;
  wire [13:0] _GEN_14366 = 14'h381e == index ? 14'h196 : _GEN_14365;
  wire [13:0] _GEN_14367 = 14'h381f == index ? 14'h193 : _GEN_14366;
  wire [13:0] _GEN_14368 = 14'h3820 == index ? 14'h190 : _GEN_14367;
  wire [13:0] _GEN_14369 = 14'h3821 == index ? 14'h18d : _GEN_14368;
  wire [13:0] _GEN_14370 = 14'h3822 == index ? 14'h18a : _GEN_14369;
  wire [13:0] _GEN_14371 = 14'h3823 == index ? 14'h187 : _GEN_14370;
  wire [13:0] _GEN_14372 = 14'h3824 == index ? 14'h184 : _GEN_14371;
  wire [13:0] _GEN_14373 = 14'h3825 == index ? 14'h181 : _GEN_14372;
  wire [13:0] _GEN_14374 = 14'h3826 == index ? 14'h124 : _GEN_14373;
  wire [13:0] _GEN_14375 = 14'h3827 == index ? 14'h122 : _GEN_14374;
  wire [13:0] _GEN_14376 = 14'h3828 == index ? 14'h120 : _GEN_14375;
  wire [13:0] _GEN_14377 = 14'h3829 == index ? 14'h11e : _GEN_14376;
  wire [13:0] _GEN_14378 = 14'h382a == index ? 14'h11c : _GEN_14377;
  wire [13:0] _GEN_14379 = 14'h382b == index ? 14'h11a : _GEN_14378;
  wire [13:0] _GEN_14380 = 14'h382c == index ? 14'h118 : _GEN_14379;
  wire [13:0] _GEN_14381 = 14'h382d == index ? 14'h116 : _GEN_14380;
  wire [13:0] _GEN_14382 = 14'h382e == index ? 14'h114 : _GEN_14381;
  wire [13:0] _GEN_14383 = 14'h382f == index ? 14'h112 : _GEN_14382;
  wire [13:0] _GEN_14384 = 14'h3830 == index ? 14'h110 : _GEN_14383;
  wire [13:0] _GEN_14385 = 14'h3831 == index ? 14'h10e : _GEN_14384;
  wire [13:0] _GEN_14386 = 14'h3832 == index ? 14'h10c : _GEN_14385;
  wire [13:0] _GEN_14387 = 14'h3833 == index ? 14'h10a : _GEN_14386;
  wire [13:0] _GEN_14388 = 14'h3834 == index ? 14'h108 : _GEN_14387;
  wire [13:0] _GEN_14389 = 14'h3835 == index ? 14'h106 : _GEN_14388;
  wire [13:0] _GEN_14390 = 14'h3836 == index ? 14'h104 : _GEN_14389;
  wire [13:0] _GEN_14391 = 14'h3837 == index ? 14'h102 : _GEN_14390;
  wire [13:0] _GEN_14392 = 14'h3838 == index ? 14'h100 : _GEN_14391;
  wire [13:0] _GEN_14393 = 14'h3839 == index ? 14'hb7 : _GEN_14392;
  wire [13:0] _GEN_14394 = 14'h383a == index ? 14'hb6 : _GEN_14393;
  wire [13:0] _GEN_14395 = 14'h383b == index ? 14'hb5 : _GEN_14394;
  wire [13:0] _GEN_14396 = 14'h383c == index ? 14'hb4 : _GEN_14395;
  wire [13:0] _GEN_14397 = 14'h383d == index ? 14'hb3 : _GEN_14396;
  wire [13:0] _GEN_14398 = 14'h383e == index ? 14'hb2 : _GEN_14397;
  wire [13:0] _GEN_14399 = 14'h383f == index ? 14'hb1 : _GEN_14398;
  wire [13:0] _GEN_14400 = 14'h3840 == index ? 14'hb0 : _GEN_14399;
  wire [13:0] _GEN_14401 = 14'h3841 == index ? 14'haf : _GEN_14400;
  wire [13:0] _GEN_14402 = 14'h3842 == index ? 14'hae : _GEN_14401;
  wire [13:0] _GEN_14403 = 14'h3843 == index ? 14'had : _GEN_14402;
  wire [13:0] _GEN_14404 = 14'h3844 == index ? 14'hac : _GEN_14403;
  wire [13:0] _GEN_14405 = 14'h3845 == index ? 14'hab : _GEN_14404;
  wire [13:0] _GEN_14406 = 14'h3846 == index ? 14'haa : _GEN_14405;
  wire [13:0] _GEN_14407 = 14'h3847 == index ? 14'ha9 : _GEN_14406;
  wire [13:0] _GEN_14408 = 14'h3848 == index ? 14'ha8 : _GEN_14407;
  wire [13:0] _GEN_14409 = 14'h3849 == index ? 14'ha7 : _GEN_14408;
  wire [13:0] _GEN_14410 = 14'h384a == index ? 14'ha6 : _GEN_14409;
  wire [13:0] _GEN_14411 = 14'h384b == index ? 14'ha5 : _GEN_14410;
  wire [13:0] _GEN_14412 = 14'h384c == index ? 14'ha4 : _GEN_14411;
  wire [13:0] _GEN_14413 = 14'h384d == index ? 14'ha3 : _GEN_14412;
  wire [13:0] _GEN_14414 = 14'h384e == index ? 14'ha2 : _GEN_14413;
  wire [13:0] _GEN_14415 = 14'h384f == index ? 14'ha1 : _GEN_14414;
  wire [13:0] _GEN_14416 = 14'h3850 == index ? 14'ha0 : _GEN_14415;
  wire [13:0] _GEN_14417 = 14'h3851 == index ? 14'h9f : _GEN_14416;
  wire [13:0] _GEN_14418 = 14'h3852 == index ? 14'h9e : _GEN_14417;
  wire [13:0] _GEN_14419 = 14'h3853 == index ? 14'h9d : _GEN_14418;
  wire [13:0] _GEN_14420 = 14'h3854 == index ? 14'h9c : _GEN_14419;
  wire [13:0] _GEN_14421 = 14'h3855 == index ? 14'h9b : _GEN_14420;
  wire [13:0] _GEN_14422 = 14'h3856 == index ? 14'h9a : _GEN_14421;
  wire [13:0] _GEN_14423 = 14'h3857 == index ? 14'h99 : _GEN_14422;
  wire [13:0] _GEN_14424 = 14'h3858 == index ? 14'h98 : _GEN_14423;
  wire [13:0] _GEN_14425 = 14'h3859 == index ? 14'h97 : _GEN_14424;
  wire [13:0] _GEN_14426 = 14'h385a == index ? 14'h96 : _GEN_14425;
  wire [13:0] _GEN_14427 = 14'h385b == index ? 14'h95 : _GEN_14426;
  wire [13:0] _GEN_14428 = 14'h385c == index ? 14'h94 : _GEN_14427;
  wire [13:0] _GEN_14429 = 14'h385d == index ? 14'h93 : _GEN_14428;
  wire [13:0] _GEN_14430 = 14'h385e == index ? 14'h92 : _GEN_14429;
  wire [13:0] _GEN_14431 = 14'h385f == index ? 14'h91 : _GEN_14430;
  wire [13:0] _GEN_14432 = 14'h3860 == index ? 14'h90 : _GEN_14431;
  wire [13:0] _GEN_14433 = 14'h3861 == index ? 14'h8f : _GEN_14432;
  wire [13:0] _GEN_14434 = 14'h3862 == index ? 14'h8e : _GEN_14433;
  wire [13:0] _GEN_14435 = 14'h3863 == index ? 14'h8d : _GEN_14434;
  wire [13:0] _GEN_14436 = 14'h3864 == index ? 14'h8c : _GEN_14435;
  wire [13:0] _GEN_14437 = 14'h3865 == index ? 14'h8b : _GEN_14436;
  wire [13:0] _GEN_14438 = 14'h3866 == index ? 14'h8a : _GEN_14437;
  wire [13:0] _GEN_14439 = 14'h3867 == index ? 14'h89 : _GEN_14438;
  wire [13:0] _GEN_14440 = 14'h3868 == index ? 14'h88 : _GEN_14439;
  wire [13:0] _GEN_14441 = 14'h3869 == index ? 14'h87 : _GEN_14440;
  wire [13:0] _GEN_14442 = 14'h386a == index ? 14'h86 : _GEN_14441;
  wire [13:0] _GEN_14443 = 14'h386b == index ? 14'h85 : _GEN_14442;
  wire [13:0] _GEN_14444 = 14'h386c == index ? 14'h84 : _GEN_14443;
  wire [13:0] _GEN_14445 = 14'h386d == index ? 14'h83 : _GEN_14444;
  wire [13:0] _GEN_14446 = 14'h386e == index ? 14'h82 : _GEN_14445;
  wire [13:0] _GEN_14447 = 14'h386f == index ? 14'h81 : _GEN_14446;
  wire [13:0] _GEN_14448 = 14'h3870 == index ? 14'h80 : _GEN_14447;
  wire [13:0] _GEN_14449 = 14'h3871 == index ? 14'h70 : _GEN_14448;
  wire [13:0] _GEN_14450 = 14'h3872 == index ? 14'h70 : _GEN_14449;
  wire [13:0] _GEN_14451 = 14'h3873 == index ? 14'h70 : _GEN_14450;
  wire [13:0] _GEN_14452 = 14'h3874 == index ? 14'h70 : _GEN_14451;
  wire [13:0] _GEN_14453 = 14'h3875 == index ? 14'h70 : _GEN_14452;
  wire [13:0] _GEN_14454 = 14'h3876 == index ? 14'h70 : _GEN_14453;
  wire [13:0] _GEN_14455 = 14'h3877 == index ? 14'h70 : _GEN_14454;
  wire [13:0] _GEN_14456 = 14'h3878 == index ? 14'h70 : _GEN_14455;
  wire [13:0] _GEN_14457 = 14'h3879 == index ? 14'h70 : _GEN_14456;
  wire [13:0] _GEN_14458 = 14'h387a == index ? 14'h70 : _GEN_14457;
  wire [13:0] _GEN_14459 = 14'h387b == index ? 14'h70 : _GEN_14458;
  wire [13:0] _GEN_14460 = 14'h387c == index ? 14'h70 : _GEN_14459;
  wire [13:0] _GEN_14461 = 14'h387d == index ? 14'h70 : _GEN_14460;
  wire [13:0] _GEN_14462 = 14'h387e == index ? 14'h70 : _GEN_14461;
  wire [13:0] _GEN_14463 = 14'h387f == index ? 14'h70 : _GEN_14462;
  wire [13:0] _GEN_14464 = 14'h3880 == index ? 14'h0 : _GEN_14463;
  wire [13:0] _GEN_14465 = 14'h3881 == index ? 14'h3880 : _GEN_14464;
  wire [13:0] _GEN_14466 = 14'h3882 == index ? 14'h1c01 : _GEN_14465;
  wire [13:0] _GEN_14467 = 14'h3883 == index ? 14'h1282 : _GEN_14466;
  wire [13:0] _GEN_14468 = 14'h3884 == index ? 14'he01 : _GEN_14467;
  wire [13:0] _GEN_14469 = 14'h3885 == index ? 14'hb03 : _GEN_14468;
  wire [13:0] _GEN_14470 = 14'h3886 == index ? 14'h905 : _GEN_14469;
  wire [13:0] _GEN_14471 = 14'h3887 == index ? 14'h801 : _GEN_14470;
  wire [13:0] _GEN_14472 = 14'h3888 == index ? 14'h701 : _GEN_14471;
  wire [13:0] _GEN_14473 = 14'h3889 == index ? 14'h605 : _GEN_14472;
  wire [13:0] _GEN_14474 = 14'h388a == index ? 14'h583 : _GEN_14473;
  wire [13:0] _GEN_14475 = 14'h388b == index ? 14'h503 : _GEN_14474;
  wire [13:0] _GEN_14476 = 14'h388c == index ? 14'h485 : _GEN_14475;
  wire [13:0] _GEN_14477 = 14'h388d == index ? 14'h409 : _GEN_14476;
  wire [13:0] _GEN_14478 = 14'h388e == index ? 14'h401 : _GEN_14477;
  wire [13:0] _GEN_14479 = 14'h388f == index ? 14'h388 : _GEN_14478;
  wire [13:0] _GEN_14480 = 14'h3890 == index ? 14'h381 : _GEN_14479;
  wire [13:0] _GEN_14481 = 14'h3891 == index ? 14'h30b : _GEN_14480;
  wire [13:0] _GEN_14482 = 14'h3892 == index ? 14'h305 : _GEN_14481;
  wire [13:0] _GEN_14483 = 14'h3893 == index ? 14'h292 : _GEN_14482;
  wire [13:0] _GEN_14484 = 14'h3894 == index ? 14'h28d : _GEN_14483;
  wire [13:0] _GEN_14485 = 14'h3895 == index ? 14'h288 : _GEN_14484;
  wire [13:0] _GEN_14486 = 14'h3896 == index ? 14'h283 : _GEN_14485;
  wire [13:0] _GEN_14487 = 14'h3897 == index ? 14'h215 : _GEN_14486;
  wire [13:0] _GEN_14488 = 14'h3898 == index ? 14'h211 : _GEN_14487;
  wire [13:0] _GEN_14489 = 14'h3899 == index ? 14'h20d : _GEN_14488;
  wire [13:0] _GEN_14490 = 14'h389a == index ? 14'h209 : _GEN_14489;
  wire [13:0] _GEN_14491 = 14'h389b == index ? 14'h205 : _GEN_14490;
  wire [13:0] _GEN_14492 = 14'h389c == index ? 14'h201 : _GEN_14491;
  wire [13:0] _GEN_14493 = 14'h389d == index ? 14'h19a : _GEN_14492;
  wire [13:0] _GEN_14494 = 14'h389e == index ? 14'h197 : _GEN_14493;
  wire [13:0] _GEN_14495 = 14'h389f == index ? 14'h194 : _GEN_14494;
  wire [13:0] _GEN_14496 = 14'h38a0 == index ? 14'h191 : _GEN_14495;
  wire [13:0] _GEN_14497 = 14'h38a1 == index ? 14'h18e : _GEN_14496;
  wire [13:0] _GEN_14498 = 14'h38a2 == index ? 14'h18b : _GEN_14497;
  wire [13:0] _GEN_14499 = 14'h38a3 == index ? 14'h188 : _GEN_14498;
  wire [13:0] _GEN_14500 = 14'h38a4 == index ? 14'h185 : _GEN_14499;
  wire [13:0] _GEN_14501 = 14'h38a5 == index ? 14'h182 : _GEN_14500;
  wire [13:0] _GEN_14502 = 14'h38a6 == index ? 14'h125 : _GEN_14501;
  wire [13:0] _GEN_14503 = 14'h38a7 == index ? 14'h123 : _GEN_14502;
  wire [13:0] _GEN_14504 = 14'h38a8 == index ? 14'h121 : _GEN_14503;
  wire [13:0] _GEN_14505 = 14'h38a9 == index ? 14'h11f : _GEN_14504;
  wire [13:0] _GEN_14506 = 14'h38aa == index ? 14'h11d : _GEN_14505;
  wire [13:0] _GEN_14507 = 14'h38ab == index ? 14'h11b : _GEN_14506;
  wire [13:0] _GEN_14508 = 14'h38ac == index ? 14'h119 : _GEN_14507;
  wire [13:0] _GEN_14509 = 14'h38ad == index ? 14'h117 : _GEN_14508;
  wire [13:0] _GEN_14510 = 14'h38ae == index ? 14'h115 : _GEN_14509;
  wire [13:0] _GEN_14511 = 14'h38af == index ? 14'h113 : _GEN_14510;
  wire [13:0] _GEN_14512 = 14'h38b0 == index ? 14'h111 : _GEN_14511;
  wire [13:0] _GEN_14513 = 14'h38b1 == index ? 14'h10f : _GEN_14512;
  wire [13:0] _GEN_14514 = 14'h38b2 == index ? 14'h10d : _GEN_14513;
  wire [13:0] _GEN_14515 = 14'h38b3 == index ? 14'h10b : _GEN_14514;
  wire [13:0] _GEN_14516 = 14'h38b4 == index ? 14'h109 : _GEN_14515;
  wire [13:0] _GEN_14517 = 14'h38b5 == index ? 14'h107 : _GEN_14516;
  wire [13:0] _GEN_14518 = 14'h38b6 == index ? 14'h105 : _GEN_14517;
  wire [13:0] _GEN_14519 = 14'h38b7 == index ? 14'h103 : _GEN_14518;
  wire [13:0] _GEN_14520 = 14'h38b8 == index ? 14'h101 : _GEN_14519;
  wire [13:0] _GEN_14521 = 14'h38b9 == index ? 14'hb8 : _GEN_14520;
  wire [13:0] _GEN_14522 = 14'h38ba == index ? 14'hb7 : _GEN_14521;
  wire [13:0] _GEN_14523 = 14'h38bb == index ? 14'hb6 : _GEN_14522;
  wire [13:0] _GEN_14524 = 14'h38bc == index ? 14'hb5 : _GEN_14523;
  wire [13:0] _GEN_14525 = 14'h38bd == index ? 14'hb4 : _GEN_14524;
  wire [13:0] _GEN_14526 = 14'h38be == index ? 14'hb3 : _GEN_14525;
  wire [13:0] _GEN_14527 = 14'h38bf == index ? 14'hb2 : _GEN_14526;
  wire [13:0] _GEN_14528 = 14'h38c0 == index ? 14'hb1 : _GEN_14527;
  wire [13:0] _GEN_14529 = 14'h38c1 == index ? 14'hb0 : _GEN_14528;
  wire [13:0] _GEN_14530 = 14'h38c2 == index ? 14'haf : _GEN_14529;
  wire [13:0] _GEN_14531 = 14'h38c3 == index ? 14'hae : _GEN_14530;
  wire [13:0] _GEN_14532 = 14'h38c4 == index ? 14'had : _GEN_14531;
  wire [13:0] _GEN_14533 = 14'h38c5 == index ? 14'hac : _GEN_14532;
  wire [13:0] _GEN_14534 = 14'h38c6 == index ? 14'hab : _GEN_14533;
  wire [13:0] _GEN_14535 = 14'h38c7 == index ? 14'haa : _GEN_14534;
  wire [13:0] _GEN_14536 = 14'h38c8 == index ? 14'ha9 : _GEN_14535;
  wire [13:0] _GEN_14537 = 14'h38c9 == index ? 14'ha8 : _GEN_14536;
  wire [13:0] _GEN_14538 = 14'h38ca == index ? 14'ha7 : _GEN_14537;
  wire [13:0] _GEN_14539 = 14'h38cb == index ? 14'ha6 : _GEN_14538;
  wire [13:0] _GEN_14540 = 14'h38cc == index ? 14'ha5 : _GEN_14539;
  wire [13:0] _GEN_14541 = 14'h38cd == index ? 14'ha4 : _GEN_14540;
  wire [13:0] _GEN_14542 = 14'h38ce == index ? 14'ha3 : _GEN_14541;
  wire [13:0] _GEN_14543 = 14'h38cf == index ? 14'ha2 : _GEN_14542;
  wire [13:0] _GEN_14544 = 14'h38d0 == index ? 14'ha1 : _GEN_14543;
  wire [13:0] _GEN_14545 = 14'h38d1 == index ? 14'ha0 : _GEN_14544;
  wire [13:0] _GEN_14546 = 14'h38d2 == index ? 14'h9f : _GEN_14545;
  wire [13:0] _GEN_14547 = 14'h38d3 == index ? 14'h9e : _GEN_14546;
  wire [13:0] _GEN_14548 = 14'h38d4 == index ? 14'h9d : _GEN_14547;
  wire [13:0] _GEN_14549 = 14'h38d5 == index ? 14'h9c : _GEN_14548;
  wire [13:0] _GEN_14550 = 14'h38d6 == index ? 14'h9b : _GEN_14549;
  wire [13:0] _GEN_14551 = 14'h38d7 == index ? 14'h9a : _GEN_14550;
  wire [13:0] _GEN_14552 = 14'h38d8 == index ? 14'h99 : _GEN_14551;
  wire [13:0] _GEN_14553 = 14'h38d9 == index ? 14'h98 : _GEN_14552;
  wire [13:0] _GEN_14554 = 14'h38da == index ? 14'h97 : _GEN_14553;
  wire [13:0] _GEN_14555 = 14'h38db == index ? 14'h96 : _GEN_14554;
  wire [13:0] _GEN_14556 = 14'h38dc == index ? 14'h95 : _GEN_14555;
  wire [13:0] _GEN_14557 = 14'h38dd == index ? 14'h94 : _GEN_14556;
  wire [13:0] _GEN_14558 = 14'h38de == index ? 14'h93 : _GEN_14557;
  wire [13:0] _GEN_14559 = 14'h38df == index ? 14'h92 : _GEN_14558;
  wire [13:0] _GEN_14560 = 14'h38e0 == index ? 14'h91 : _GEN_14559;
  wire [13:0] _GEN_14561 = 14'h38e1 == index ? 14'h90 : _GEN_14560;
  wire [13:0] _GEN_14562 = 14'h38e2 == index ? 14'h8f : _GEN_14561;
  wire [13:0] _GEN_14563 = 14'h38e3 == index ? 14'h8e : _GEN_14562;
  wire [13:0] _GEN_14564 = 14'h38e4 == index ? 14'h8d : _GEN_14563;
  wire [13:0] _GEN_14565 = 14'h38e5 == index ? 14'h8c : _GEN_14564;
  wire [13:0] _GEN_14566 = 14'h38e6 == index ? 14'h8b : _GEN_14565;
  wire [13:0] _GEN_14567 = 14'h38e7 == index ? 14'h8a : _GEN_14566;
  wire [13:0] _GEN_14568 = 14'h38e8 == index ? 14'h89 : _GEN_14567;
  wire [13:0] _GEN_14569 = 14'h38e9 == index ? 14'h88 : _GEN_14568;
  wire [13:0] _GEN_14570 = 14'h38ea == index ? 14'h87 : _GEN_14569;
  wire [13:0] _GEN_14571 = 14'h38eb == index ? 14'h86 : _GEN_14570;
  wire [13:0] _GEN_14572 = 14'h38ec == index ? 14'h85 : _GEN_14571;
  wire [13:0] _GEN_14573 = 14'h38ed == index ? 14'h84 : _GEN_14572;
  wire [13:0] _GEN_14574 = 14'h38ee == index ? 14'h83 : _GEN_14573;
  wire [13:0] _GEN_14575 = 14'h38ef == index ? 14'h82 : _GEN_14574;
  wire [13:0] _GEN_14576 = 14'h38f0 == index ? 14'h81 : _GEN_14575;
  wire [13:0] _GEN_14577 = 14'h38f1 == index ? 14'h80 : _GEN_14576;
  wire [13:0] _GEN_14578 = 14'h38f2 == index ? 14'h71 : _GEN_14577;
  wire [13:0] _GEN_14579 = 14'h38f3 == index ? 14'h71 : _GEN_14578;
  wire [13:0] _GEN_14580 = 14'h38f4 == index ? 14'h71 : _GEN_14579;
  wire [13:0] _GEN_14581 = 14'h38f5 == index ? 14'h71 : _GEN_14580;
  wire [13:0] _GEN_14582 = 14'h38f6 == index ? 14'h71 : _GEN_14581;
  wire [13:0] _GEN_14583 = 14'h38f7 == index ? 14'h71 : _GEN_14582;
  wire [13:0] _GEN_14584 = 14'h38f8 == index ? 14'h71 : _GEN_14583;
  wire [13:0] _GEN_14585 = 14'h38f9 == index ? 14'h71 : _GEN_14584;
  wire [13:0] _GEN_14586 = 14'h38fa == index ? 14'h71 : _GEN_14585;
  wire [13:0] _GEN_14587 = 14'h38fb == index ? 14'h71 : _GEN_14586;
  wire [13:0] _GEN_14588 = 14'h38fc == index ? 14'h71 : _GEN_14587;
  wire [13:0] _GEN_14589 = 14'h38fd == index ? 14'h71 : _GEN_14588;
  wire [13:0] _GEN_14590 = 14'h38fe == index ? 14'h71 : _GEN_14589;
  wire [13:0] _GEN_14591 = 14'h38ff == index ? 14'h71 : _GEN_14590;
  wire [13:0] _GEN_14592 = 14'h3900 == index ? 14'h0 : _GEN_14591;
  wire [13:0] _GEN_14593 = 14'h3901 == index ? 14'h3900 : _GEN_14592;
  wire [13:0] _GEN_14594 = 14'h3902 == index ? 14'h1c80 : _GEN_14593;
  wire [13:0] _GEN_14595 = 14'h3903 == index ? 14'h1300 : _GEN_14594;
  wire [13:0] _GEN_14596 = 14'h3904 == index ? 14'he02 : _GEN_14595;
  wire [13:0] _GEN_14597 = 14'h3905 == index ? 14'hb04 : _GEN_14596;
  wire [13:0] _GEN_14598 = 14'h3906 == index ? 14'h980 : _GEN_14597;
  wire [13:0] _GEN_14599 = 14'h3907 == index ? 14'h802 : _GEN_14598;
  wire [13:0] _GEN_14600 = 14'h3908 == index ? 14'h702 : _GEN_14599;
  wire [13:0] _GEN_14601 = 14'h3909 == index ? 14'h606 : _GEN_14600;
  wire [13:0] _GEN_14602 = 14'h390a == index ? 14'h584 : _GEN_14601;
  wire [13:0] _GEN_14603 = 14'h390b == index ? 14'h504 : _GEN_14602;
  wire [13:0] _GEN_14604 = 14'h390c == index ? 14'h486 : _GEN_14603;
  wire [13:0] _GEN_14605 = 14'h390d == index ? 14'h40a : _GEN_14604;
  wire [13:0] _GEN_14606 = 14'h390e == index ? 14'h402 : _GEN_14605;
  wire [13:0] _GEN_14607 = 14'h390f == index ? 14'h389 : _GEN_14606;
  wire [13:0] _GEN_14608 = 14'h3910 == index ? 14'h382 : _GEN_14607;
  wire [13:0] _GEN_14609 = 14'h3911 == index ? 14'h30c : _GEN_14608;
  wire [13:0] _GEN_14610 = 14'h3912 == index ? 14'h306 : _GEN_14609;
  wire [13:0] _GEN_14611 = 14'h3913 == index ? 14'h300 : _GEN_14610;
  wire [13:0] _GEN_14612 = 14'h3914 == index ? 14'h28e : _GEN_14611;
  wire [13:0] _GEN_14613 = 14'h3915 == index ? 14'h289 : _GEN_14612;
  wire [13:0] _GEN_14614 = 14'h3916 == index ? 14'h284 : _GEN_14613;
  wire [13:0] _GEN_14615 = 14'h3917 == index ? 14'h216 : _GEN_14614;
  wire [13:0] _GEN_14616 = 14'h3918 == index ? 14'h212 : _GEN_14615;
  wire [13:0] _GEN_14617 = 14'h3919 == index ? 14'h20e : _GEN_14616;
  wire [13:0] _GEN_14618 = 14'h391a == index ? 14'h20a : _GEN_14617;
  wire [13:0] _GEN_14619 = 14'h391b == index ? 14'h206 : _GEN_14618;
  wire [13:0] _GEN_14620 = 14'h391c == index ? 14'h202 : _GEN_14619;
  wire [13:0] _GEN_14621 = 14'h391d == index ? 14'h19b : _GEN_14620;
  wire [13:0] _GEN_14622 = 14'h391e == index ? 14'h198 : _GEN_14621;
  wire [13:0] _GEN_14623 = 14'h391f == index ? 14'h195 : _GEN_14622;
  wire [13:0] _GEN_14624 = 14'h3920 == index ? 14'h192 : _GEN_14623;
  wire [13:0] _GEN_14625 = 14'h3921 == index ? 14'h18f : _GEN_14624;
  wire [13:0] _GEN_14626 = 14'h3922 == index ? 14'h18c : _GEN_14625;
  wire [13:0] _GEN_14627 = 14'h3923 == index ? 14'h189 : _GEN_14626;
  wire [13:0] _GEN_14628 = 14'h3924 == index ? 14'h186 : _GEN_14627;
  wire [13:0] _GEN_14629 = 14'h3925 == index ? 14'h183 : _GEN_14628;
  wire [13:0] _GEN_14630 = 14'h3926 == index ? 14'h180 : _GEN_14629;
  wire [13:0] _GEN_14631 = 14'h3927 == index ? 14'h124 : _GEN_14630;
  wire [13:0] _GEN_14632 = 14'h3928 == index ? 14'h122 : _GEN_14631;
  wire [13:0] _GEN_14633 = 14'h3929 == index ? 14'h120 : _GEN_14632;
  wire [13:0] _GEN_14634 = 14'h392a == index ? 14'h11e : _GEN_14633;
  wire [13:0] _GEN_14635 = 14'h392b == index ? 14'h11c : _GEN_14634;
  wire [13:0] _GEN_14636 = 14'h392c == index ? 14'h11a : _GEN_14635;
  wire [13:0] _GEN_14637 = 14'h392d == index ? 14'h118 : _GEN_14636;
  wire [13:0] _GEN_14638 = 14'h392e == index ? 14'h116 : _GEN_14637;
  wire [13:0] _GEN_14639 = 14'h392f == index ? 14'h114 : _GEN_14638;
  wire [13:0] _GEN_14640 = 14'h3930 == index ? 14'h112 : _GEN_14639;
  wire [13:0] _GEN_14641 = 14'h3931 == index ? 14'h110 : _GEN_14640;
  wire [13:0] _GEN_14642 = 14'h3932 == index ? 14'h10e : _GEN_14641;
  wire [13:0] _GEN_14643 = 14'h3933 == index ? 14'h10c : _GEN_14642;
  wire [13:0] _GEN_14644 = 14'h3934 == index ? 14'h10a : _GEN_14643;
  wire [13:0] _GEN_14645 = 14'h3935 == index ? 14'h108 : _GEN_14644;
  wire [13:0] _GEN_14646 = 14'h3936 == index ? 14'h106 : _GEN_14645;
  wire [13:0] _GEN_14647 = 14'h3937 == index ? 14'h104 : _GEN_14646;
  wire [13:0] _GEN_14648 = 14'h3938 == index ? 14'h102 : _GEN_14647;
  wire [13:0] _GEN_14649 = 14'h3939 == index ? 14'h100 : _GEN_14648;
  wire [13:0] _GEN_14650 = 14'h393a == index ? 14'hb8 : _GEN_14649;
  wire [13:0] _GEN_14651 = 14'h393b == index ? 14'hb7 : _GEN_14650;
  wire [13:0] _GEN_14652 = 14'h393c == index ? 14'hb6 : _GEN_14651;
  wire [13:0] _GEN_14653 = 14'h393d == index ? 14'hb5 : _GEN_14652;
  wire [13:0] _GEN_14654 = 14'h393e == index ? 14'hb4 : _GEN_14653;
  wire [13:0] _GEN_14655 = 14'h393f == index ? 14'hb3 : _GEN_14654;
  wire [13:0] _GEN_14656 = 14'h3940 == index ? 14'hb2 : _GEN_14655;
  wire [13:0] _GEN_14657 = 14'h3941 == index ? 14'hb1 : _GEN_14656;
  wire [13:0] _GEN_14658 = 14'h3942 == index ? 14'hb0 : _GEN_14657;
  wire [13:0] _GEN_14659 = 14'h3943 == index ? 14'haf : _GEN_14658;
  wire [13:0] _GEN_14660 = 14'h3944 == index ? 14'hae : _GEN_14659;
  wire [13:0] _GEN_14661 = 14'h3945 == index ? 14'had : _GEN_14660;
  wire [13:0] _GEN_14662 = 14'h3946 == index ? 14'hac : _GEN_14661;
  wire [13:0] _GEN_14663 = 14'h3947 == index ? 14'hab : _GEN_14662;
  wire [13:0] _GEN_14664 = 14'h3948 == index ? 14'haa : _GEN_14663;
  wire [13:0] _GEN_14665 = 14'h3949 == index ? 14'ha9 : _GEN_14664;
  wire [13:0] _GEN_14666 = 14'h394a == index ? 14'ha8 : _GEN_14665;
  wire [13:0] _GEN_14667 = 14'h394b == index ? 14'ha7 : _GEN_14666;
  wire [13:0] _GEN_14668 = 14'h394c == index ? 14'ha6 : _GEN_14667;
  wire [13:0] _GEN_14669 = 14'h394d == index ? 14'ha5 : _GEN_14668;
  wire [13:0] _GEN_14670 = 14'h394e == index ? 14'ha4 : _GEN_14669;
  wire [13:0] _GEN_14671 = 14'h394f == index ? 14'ha3 : _GEN_14670;
  wire [13:0] _GEN_14672 = 14'h3950 == index ? 14'ha2 : _GEN_14671;
  wire [13:0] _GEN_14673 = 14'h3951 == index ? 14'ha1 : _GEN_14672;
  wire [13:0] _GEN_14674 = 14'h3952 == index ? 14'ha0 : _GEN_14673;
  wire [13:0] _GEN_14675 = 14'h3953 == index ? 14'h9f : _GEN_14674;
  wire [13:0] _GEN_14676 = 14'h3954 == index ? 14'h9e : _GEN_14675;
  wire [13:0] _GEN_14677 = 14'h3955 == index ? 14'h9d : _GEN_14676;
  wire [13:0] _GEN_14678 = 14'h3956 == index ? 14'h9c : _GEN_14677;
  wire [13:0] _GEN_14679 = 14'h3957 == index ? 14'h9b : _GEN_14678;
  wire [13:0] _GEN_14680 = 14'h3958 == index ? 14'h9a : _GEN_14679;
  wire [13:0] _GEN_14681 = 14'h3959 == index ? 14'h99 : _GEN_14680;
  wire [13:0] _GEN_14682 = 14'h395a == index ? 14'h98 : _GEN_14681;
  wire [13:0] _GEN_14683 = 14'h395b == index ? 14'h97 : _GEN_14682;
  wire [13:0] _GEN_14684 = 14'h395c == index ? 14'h96 : _GEN_14683;
  wire [13:0] _GEN_14685 = 14'h395d == index ? 14'h95 : _GEN_14684;
  wire [13:0] _GEN_14686 = 14'h395e == index ? 14'h94 : _GEN_14685;
  wire [13:0] _GEN_14687 = 14'h395f == index ? 14'h93 : _GEN_14686;
  wire [13:0] _GEN_14688 = 14'h3960 == index ? 14'h92 : _GEN_14687;
  wire [13:0] _GEN_14689 = 14'h3961 == index ? 14'h91 : _GEN_14688;
  wire [13:0] _GEN_14690 = 14'h3962 == index ? 14'h90 : _GEN_14689;
  wire [13:0] _GEN_14691 = 14'h3963 == index ? 14'h8f : _GEN_14690;
  wire [13:0] _GEN_14692 = 14'h3964 == index ? 14'h8e : _GEN_14691;
  wire [13:0] _GEN_14693 = 14'h3965 == index ? 14'h8d : _GEN_14692;
  wire [13:0] _GEN_14694 = 14'h3966 == index ? 14'h8c : _GEN_14693;
  wire [13:0] _GEN_14695 = 14'h3967 == index ? 14'h8b : _GEN_14694;
  wire [13:0] _GEN_14696 = 14'h3968 == index ? 14'h8a : _GEN_14695;
  wire [13:0] _GEN_14697 = 14'h3969 == index ? 14'h89 : _GEN_14696;
  wire [13:0] _GEN_14698 = 14'h396a == index ? 14'h88 : _GEN_14697;
  wire [13:0] _GEN_14699 = 14'h396b == index ? 14'h87 : _GEN_14698;
  wire [13:0] _GEN_14700 = 14'h396c == index ? 14'h86 : _GEN_14699;
  wire [13:0] _GEN_14701 = 14'h396d == index ? 14'h85 : _GEN_14700;
  wire [13:0] _GEN_14702 = 14'h396e == index ? 14'h84 : _GEN_14701;
  wire [13:0] _GEN_14703 = 14'h396f == index ? 14'h83 : _GEN_14702;
  wire [13:0] _GEN_14704 = 14'h3970 == index ? 14'h82 : _GEN_14703;
  wire [13:0] _GEN_14705 = 14'h3971 == index ? 14'h81 : _GEN_14704;
  wire [13:0] _GEN_14706 = 14'h3972 == index ? 14'h80 : _GEN_14705;
  wire [13:0] _GEN_14707 = 14'h3973 == index ? 14'h72 : _GEN_14706;
  wire [13:0] _GEN_14708 = 14'h3974 == index ? 14'h72 : _GEN_14707;
  wire [13:0] _GEN_14709 = 14'h3975 == index ? 14'h72 : _GEN_14708;
  wire [13:0] _GEN_14710 = 14'h3976 == index ? 14'h72 : _GEN_14709;
  wire [13:0] _GEN_14711 = 14'h3977 == index ? 14'h72 : _GEN_14710;
  wire [13:0] _GEN_14712 = 14'h3978 == index ? 14'h72 : _GEN_14711;
  wire [13:0] _GEN_14713 = 14'h3979 == index ? 14'h72 : _GEN_14712;
  wire [13:0] _GEN_14714 = 14'h397a == index ? 14'h72 : _GEN_14713;
  wire [13:0] _GEN_14715 = 14'h397b == index ? 14'h72 : _GEN_14714;
  wire [13:0] _GEN_14716 = 14'h397c == index ? 14'h72 : _GEN_14715;
  wire [13:0] _GEN_14717 = 14'h397d == index ? 14'h72 : _GEN_14716;
  wire [13:0] _GEN_14718 = 14'h397e == index ? 14'h72 : _GEN_14717;
  wire [13:0] _GEN_14719 = 14'h397f == index ? 14'h72 : _GEN_14718;
  wire [13:0] _GEN_14720 = 14'h3980 == index ? 14'h0 : _GEN_14719;
  wire [13:0] _GEN_14721 = 14'h3981 == index ? 14'h3980 : _GEN_14720;
  wire [13:0] _GEN_14722 = 14'h3982 == index ? 14'h1c81 : _GEN_14721;
  wire [13:0] _GEN_14723 = 14'h3983 == index ? 14'h1301 : _GEN_14722;
  wire [13:0] _GEN_14724 = 14'h3984 == index ? 14'he03 : _GEN_14723;
  wire [13:0] _GEN_14725 = 14'h3985 == index ? 14'hb80 : _GEN_14724;
  wire [13:0] _GEN_14726 = 14'h3986 == index ? 14'h981 : _GEN_14725;
  wire [13:0] _GEN_14727 = 14'h3987 == index ? 14'h803 : _GEN_14726;
  wire [13:0] _GEN_14728 = 14'h3988 == index ? 14'h703 : _GEN_14727;
  wire [13:0] _GEN_14729 = 14'h3989 == index ? 14'h607 : _GEN_14728;
  wire [13:0] _GEN_14730 = 14'h398a == index ? 14'h585 : _GEN_14729;
  wire [13:0] _GEN_14731 = 14'h398b == index ? 14'h505 : _GEN_14730;
  wire [13:0] _GEN_14732 = 14'h398c == index ? 14'h487 : _GEN_14731;
  wire [13:0] _GEN_14733 = 14'h398d == index ? 14'h40b : _GEN_14732;
  wire [13:0] _GEN_14734 = 14'h398e == index ? 14'h403 : _GEN_14733;
  wire [13:0] _GEN_14735 = 14'h398f == index ? 14'h38a : _GEN_14734;
  wire [13:0] _GEN_14736 = 14'h3990 == index ? 14'h383 : _GEN_14735;
  wire [13:0] _GEN_14737 = 14'h3991 == index ? 14'h30d : _GEN_14736;
  wire [13:0] _GEN_14738 = 14'h3992 == index ? 14'h307 : _GEN_14737;
  wire [13:0] _GEN_14739 = 14'h3993 == index ? 14'h301 : _GEN_14738;
  wire [13:0] _GEN_14740 = 14'h3994 == index ? 14'h28f : _GEN_14739;
  wire [13:0] _GEN_14741 = 14'h3995 == index ? 14'h28a : _GEN_14740;
  wire [13:0] _GEN_14742 = 14'h3996 == index ? 14'h285 : _GEN_14741;
  wire [13:0] _GEN_14743 = 14'h3997 == index ? 14'h280 : _GEN_14742;
  wire [13:0] _GEN_14744 = 14'h3998 == index ? 14'h213 : _GEN_14743;
  wire [13:0] _GEN_14745 = 14'h3999 == index ? 14'h20f : _GEN_14744;
  wire [13:0] _GEN_14746 = 14'h399a == index ? 14'h20b : _GEN_14745;
  wire [13:0] _GEN_14747 = 14'h399b == index ? 14'h207 : _GEN_14746;
  wire [13:0] _GEN_14748 = 14'h399c == index ? 14'h203 : _GEN_14747;
  wire [13:0] _GEN_14749 = 14'h399d == index ? 14'h19c : _GEN_14748;
  wire [13:0] _GEN_14750 = 14'h399e == index ? 14'h199 : _GEN_14749;
  wire [13:0] _GEN_14751 = 14'h399f == index ? 14'h196 : _GEN_14750;
  wire [13:0] _GEN_14752 = 14'h39a0 == index ? 14'h193 : _GEN_14751;
  wire [13:0] _GEN_14753 = 14'h39a1 == index ? 14'h190 : _GEN_14752;
  wire [13:0] _GEN_14754 = 14'h39a2 == index ? 14'h18d : _GEN_14753;
  wire [13:0] _GEN_14755 = 14'h39a3 == index ? 14'h18a : _GEN_14754;
  wire [13:0] _GEN_14756 = 14'h39a4 == index ? 14'h187 : _GEN_14755;
  wire [13:0] _GEN_14757 = 14'h39a5 == index ? 14'h184 : _GEN_14756;
  wire [13:0] _GEN_14758 = 14'h39a6 == index ? 14'h181 : _GEN_14757;
  wire [13:0] _GEN_14759 = 14'h39a7 == index ? 14'h125 : _GEN_14758;
  wire [13:0] _GEN_14760 = 14'h39a8 == index ? 14'h123 : _GEN_14759;
  wire [13:0] _GEN_14761 = 14'h39a9 == index ? 14'h121 : _GEN_14760;
  wire [13:0] _GEN_14762 = 14'h39aa == index ? 14'h11f : _GEN_14761;
  wire [13:0] _GEN_14763 = 14'h39ab == index ? 14'h11d : _GEN_14762;
  wire [13:0] _GEN_14764 = 14'h39ac == index ? 14'h11b : _GEN_14763;
  wire [13:0] _GEN_14765 = 14'h39ad == index ? 14'h119 : _GEN_14764;
  wire [13:0] _GEN_14766 = 14'h39ae == index ? 14'h117 : _GEN_14765;
  wire [13:0] _GEN_14767 = 14'h39af == index ? 14'h115 : _GEN_14766;
  wire [13:0] _GEN_14768 = 14'h39b0 == index ? 14'h113 : _GEN_14767;
  wire [13:0] _GEN_14769 = 14'h39b1 == index ? 14'h111 : _GEN_14768;
  wire [13:0] _GEN_14770 = 14'h39b2 == index ? 14'h10f : _GEN_14769;
  wire [13:0] _GEN_14771 = 14'h39b3 == index ? 14'h10d : _GEN_14770;
  wire [13:0] _GEN_14772 = 14'h39b4 == index ? 14'h10b : _GEN_14771;
  wire [13:0] _GEN_14773 = 14'h39b5 == index ? 14'h109 : _GEN_14772;
  wire [13:0] _GEN_14774 = 14'h39b6 == index ? 14'h107 : _GEN_14773;
  wire [13:0] _GEN_14775 = 14'h39b7 == index ? 14'h105 : _GEN_14774;
  wire [13:0] _GEN_14776 = 14'h39b8 == index ? 14'h103 : _GEN_14775;
  wire [13:0] _GEN_14777 = 14'h39b9 == index ? 14'h101 : _GEN_14776;
  wire [13:0] _GEN_14778 = 14'h39ba == index ? 14'hb9 : _GEN_14777;
  wire [13:0] _GEN_14779 = 14'h39bb == index ? 14'hb8 : _GEN_14778;
  wire [13:0] _GEN_14780 = 14'h39bc == index ? 14'hb7 : _GEN_14779;
  wire [13:0] _GEN_14781 = 14'h39bd == index ? 14'hb6 : _GEN_14780;
  wire [13:0] _GEN_14782 = 14'h39be == index ? 14'hb5 : _GEN_14781;
  wire [13:0] _GEN_14783 = 14'h39bf == index ? 14'hb4 : _GEN_14782;
  wire [13:0] _GEN_14784 = 14'h39c0 == index ? 14'hb3 : _GEN_14783;
  wire [13:0] _GEN_14785 = 14'h39c1 == index ? 14'hb2 : _GEN_14784;
  wire [13:0] _GEN_14786 = 14'h39c2 == index ? 14'hb1 : _GEN_14785;
  wire [13:0] _GEN_14787 = 14'h39c3 == index ? 14'hb0 : _GEN_14786;
  wire [13:0] _GEN_14788 = 14'h39c4 == index ? 14'haf : _GEN_14787;
  wire [13:0] _GEN_14789 = 14'h39c5 == index ? 14'hae : _GEN_14788;
  wire [13:0] _GEN_14790 = 14'h39c6 == index ? 14'had : _GEN_14789;
  wire [13:0] _GEN_14791 = 14'h39c7 == index ? 14'hac : _GEN_14790;
  wire [13:0] _GEN_14792 = 14'h39c8 == index ? 14'hab : _GEN_14791;
  wire [13:0] _GEN_14793 = 14'h39c9 == index ? 14'haa : _GEN_14792;
  wire [13:0] _GEN_14794 = 14'h39ca == index ? 14'ha9 : _GEN_14793;
  wire [13:0] _GEN_14795 = 14'h39cb == index ? 14'ha8 : _GEN_14794;
  wire [13:0] _GEN_14796 = 14'h39cc == index ? 14'ha7 : _GEN_14795;
  wire [13:0] _GEN_14797 = 14'h39cd == index ? 14'ha6 : _GEN_14796;
  wire [13:0] _GEN_14798 = 14'h39ce == index ? 14'ha5 : _GEN_14797;
  wire [13:0] _GEN_14799 = 14'h39cf == index ? 14'ha4 : _GEN_14798;
  wire [13:0] _GEN_14800 = 14'h39d0 == index ? 14'ha3 : _GEN_14799;
  wire [13:0] _GEN_14801 = 14'h39d1 == index ? 14'ha2 : _GEN_14800;
  wire [13:0] _GEN_14802 = 14'h39d2 == index ? 14'ha1 : _GEN_14801;
  wire [13:0] _GEN_14803 = 14'h39d3 == index ? 14'ha0 : _GEN_14802;
  wire [13:0] _GEN_14804 = 14'h39d4 == index ? 14'h9f : _GEN_14803;
  wire [13:0] _GEN_14805 = 14'h39d5 == index ? 14'h9e : _GEN_14804;
  wire [13:0] _GEN_14806 = 14'h39d6 == index ? 14'h9d : _GEN_14805;
  wire [13:0] _GEN_14807 = 14'h39d7 == index ? 14'h9c : _GEN_14806;
  wire [13:0] _GEN_14808 = 14'h39d8 == index ? 14'h9b : _GEN_14807;
  wire [13:0] _GEN_14809 = 14'h39d9 == index ? 14'h9a : _GEN_14808;
  wire [13:0] _GEN_14810 = 14'h39da == index ? 14'h99 : _GEN_14809;
  wire [13:0] _GEN_14811 = 14'h39db == index ? 14'h98 : _GEN_14810;
  wire [13:0] _GEN_14812 = 14'h39dc == index ? 14'h97 : _GEN_14811;
  wire [13:0] _GEN_14813 = 14'h39dd == index ? 14'h96 : _GEN_14812;
  wire [13:0] _GEN_14814 = 14'h39de == index ? 14'h95 : _GEN_14813;
  wire [13:0] _GEN_14815 = 14'h39df == index ? 14'h94 : _GEN_14814;
  wire [13:0] _GEN_14816 = 14'h39e0 == index ? 14'h93 : _GEN_14815;
  wire [13:0] _GEN_14817 = 14'h39e1 == index ? 14'h92 : _GEN_14816;
  wire [13:0] _GEN_14818 = 14'h39e2 == index ? 14'h91 : _GEN_14817;
  wire [13:0] _GEN_14819 = 14'h39e3 == index ? 14'h90 : _GEN_14818;
  wire [13:0] _GEN_14820 = 14'h39e4 == index ? 14'h8f : _GEN_14819;
  wire [13:0] _GEN_14821 = 14'h39e5 == index ? 14'h8e : _GEN_14820;
  wire [13:0] _GEN_14822 = 14'h39e6 == index ? 14'h8d : _GEN_14821;
  wire [13:0] _GEN_14823 = 14'h39e7 == index ? 14'h8c : _GEN_14822;
  wire [13:0] _GEN_14824 = 14'h39e8 == index ? 14'h8b : _GEN_14823;
  wire [13:0] _GEN_14825 = 14'h39e9 == index ? 14'h8a : _GEN_14824;
  wire [13:0] _GEN_14826 = 14'h39ea == index ? 14'h89 : _GEN_14825;
  wire [13:0] _GEN_14827 = 14'h39eb == index ? 14'h88 : _GEN_14826;
  wire [13:0] _GEN_14828 = 14'h39ec == index ? 14'h87 : _GEN_14827;
  wire [13:0] _GEN_14829 = 14'h39ed == index ? 14'h86 : _GEN_14828;
  wire [13:0] _GEN_14830 = 14'h39ee == index ? 14'h85 : _GEN_14829;
  wire [13:0] _GEN_14831 = 14'h39ef == index ? 14'h84 : _GEN_14830;
  wire [13:0] _GEN_14832 = 14'h39f0 == index ? 14'h83 : _GEN_14831;
  wire [13:0] _GEN_14833 = 14'h39f1 == index ? 14'h82 : _GEN_14832;
  wire [13:0] _GEN_14834 = 14'h39f2 == index ? 14'h81 : _GEN_14833;
  wire [13:0] _GEN_14835 = 14'h39f3 == index ? 14'h80 : _GEN_14834;
  wire [13:0] _GEN_14836 = 14'h39f4 == index ? 14'h73 : _GEN_14835;
  wire [13:0] _GEN_14837 = 14'h39f5 == index ? 14'h73 : _GEN_14836;
  wire [13:0] _GEN_14838 = 14'h39f6 == index ? 14'h73 : _GEN_14837;
  wire [13:0] _GEN_14839 = 14'h39f7 == index ? 14'h73 : _GEN_14838;
  wire [13:0] _GEN_14840 = 14'h39f8 == index ? 14'h73 : _GEN_14839;
  wire [13:0] _GEN_14841 = 14'h39f9 == index ? 14'h73 : _GEN_14840;
  wire [13:0] _GEN_14842 = 14'h39fa == index ? 14'h73 : _GEN_14841;
  wire [13:0] _GEN_14843 = 14'h39fb == index ? 14'h73 : _GEN_14842;
  wire [13:0] _GEN_14844 = 14'h39fc == index ? 14'h73 : _GEN_14843;
  wire [13:0] _GEN_14845 = 14'h39fd == index ? 14'h73 : _GEN_14844;
  wire [13:0] _GEN_14846 = 14'h39fe == index ? 14'h73 : _GEN_14845;
  wire [13:0] _GEN_14847 = 14'h39ff == index ? 14'h73 : _GEN_14846;
  wire [13:0] _GEN_14848 = 14'h3a00 == index ? 14'h0 : _GEN_14847;
  wire [13:0] _GEN_14849 = 14'h3a01 == index ? 14'h3a00 : _GEN_14848;
  wire [13:0] _GEN_14850 = 14'h3a02 == index ? 14'h1d00 : _GEN_14849;
  wire [13:0] _GEN_14851 = 14'h3a03 == index ? 14'h1302 : _GEN_14850;
  wire [13:0] _GEN_14852 = 14'h3a04 == index ? 14'he80 : _GEN_14851;
  wire [13:0] _GEN_14853 = 14'h3a05 == index ? 14'hb81 : _GEN_14852;
  wire [13:0] _GEN_14854 = 14'h3a06 == index ? 14'h982 : _GEN_14853;
  wire [13:0] _GEN_14855 = 14'h3a07 == index ? 14'h804 : _GEN_14854;
  wire [13:0] _GEN_14856 = 14'h3a08 == index ? 14'h704 : _GEN_14855;
  wire [13:0] _GEN_14857 = 14'h3a09 == index ? 14'h608 : _GEN_14856;
  wire [13:0] _GEN_14858 = 14'h3a0a == index ? 14'h586 : _GEN_14857;
  wire [13:0] _GEN_14859 = 14'h3a0b == index ? 14'h506 : _GEN_14858;
  wire [13:0] _GEN_14860 = 14'h3a0c == index ? 14'h488 : _GEN_14859;
  wire [13:0] _GEN_14861 = 14'h3a0d == index ? 14'h40c : _GEN_14860;
  wire [13:0] _GEN_14862 = 14'h3a0e == index ? 14'h404 : _GEN_14861;
  wire [13:0] _GEN_14863 = 14'h3a0f == index ? 14'h38b : _GEN_14862;
  wire [13:0] _GEN_14864 = 14'h3a10 == index ? 14'h384 : _GEN_14863;
  wire [13:0] _GEN_14865 = 14'h3a11 == index ? 14'h30e : _GEN_14864;
  wire [13:0] _GEN_14866 = 14'h3a12 == index ? 14'h308 : _GEN_14865;
  wire [13:0] _GEN_14867 = 14'h3a13 == index ? 14'h302 : _GEN_14866;
  wire [13:0] _GEN_14868 = 14'h3a14 == index ? 14'h290 : _GEN_14867;
  wire [13:0] _GEN_14869 = 14'h3a15 == index ? 14'h28b : _GEN_14868;
  wire [13:0] _GEN_14870 = 14'h3a16 == index ? 14'h286 : _GEN_14869;
  wire [13:0] _GEN_14871 = 14'h3a17 == index ? 14'h281 : _GEN_14870;
  wire [13:0] _GEN_14872 = 14'h3a18 == index ? 14'h214 : _GEN_14871;
  wire [13:0] _GEN_14873 = 14'h3a19 == index ? 14'h210 : _GEN_14872;
  wire [13:0] _GEN_14874 = 14'h3a1a == index ? 14'h20c : _GEN_14873;
  wire [13:0] _GEN_14875 = 14'h3a1b == index ? 14'h208 : _GEN_14874;
  wire [13:0] _GEN_14876 = 14'h3a1c == index ? 14'h204 : _GEN_14875;
  wire [13:0] _GEN_14877 = 14'h3a1d == index ? 14'h200 : _GEN_14876;
  wire [13:0] _GEN_14878 = 14'h3a1e == index ? 14'h19a : _GEN_14877;
  wire [13:0] _GEN_14879 = 14'h3a1f == index ? 14'h197 : _GEN_14878;
  wire [13:0] _GEN_14880 = 14'h3a20 == index ? 14'h194 : _GEN_14879;
  wire [13:0] _GEN_14881 = 14'h3a21 == index ? 14'h191 : _GEN_14880;
  wire [13:0] _GEN_14882 = 14'h3a22 == index ? 14'h18e : _GEN_14881;
  wire [13:0] _GEN_14883 = 14'h3a23 == index ? 14'h18b : _GEN_14882;
  wire [13:0] _GEN_14884 = 14'h3a24 == index ? 14'h188 : _GEN_14883;
  wire [13:0] _GEN_14885 = 14'h3a25 == index ? 14'h185 : _GEN_14884;
  wire [13:0] _GEN_14886 = 14'h3a26 == index ? 14'h182 : _GEN_14885;
  wire [13:0] _GEN_14887 = 14'h3a27 == index ? 14'h126 : _GEN_14886;
  wire [13:0] _GEN_14888 = 14'h3a28 == index ? 14'h124 : _GEN_14887;
  wire [13:0] _GEN_14889 = 14'h3a29 == index ? 14'h122 : _GEN_14888;
  wire [13:0] _GEN_14890 = 14'h3a2a == index ? 14'h120 : _GEN_14889;
  wire [13:0] _GEN_14891 = 14'h3a2b == index ? 14'h11e : _GEN_14890;
  wire [13:0] _GEN_14892 = 14'h3a2c == index ? 14'h11c : _GEN_14891;
  wire [13:0] _GEN_14893 = 14'h3a2d == index ? 14'h11a : _GEN_14892;
  wire [13:0] _GEN_14894 = 14'h3a2e == index ? 14'h118 : _GEN_14893;
  wire [13:0] _GEN_14895 = 14'h3a2f == index ? 14'h116 : _GEN_14894;
  wire [13:0] _GEN_14896 = 14'h3a30 == index ? 14'h114 : _GEN_14895;
  wire [13:0] _GEN_14897 = 14'h3a31 == index ? 14'h112 : _GEN_14896;
  wire [13:0] _GEN_14898 = 14'h3a32 == index ? 14'h110 : _GEN_14897;
  wire [13:0] _GEN_14899 = 14'h3a33 == index ? 14'h10e : _GEN_14898;
  wire [13:0] _GEN_14900 = 14'h3a34 == index ? 14'h10c : _GEN_14899;
  wire [13:0] _GEN_14901 = 14'h3a35 == index ? 14'h10a : _GEN_14900;
  wire [13:0] _GEN_14902 = 14'h3a36 == index ? 14'h108 : _GEN_14901;
  wire [13:0] _GEN_14903 = 14'h3a37 == index ? 14'h106 : _GEN_14902;
  wire [13:0] _GEN_14904 = 14'h3a38 == index ? 14'h104 : _GEN_14903;
  wire [13:0] _GEN_14905 = 14'h3a39 == index ? 14'h102 : _GEN_14904;
  wire [13:0] _GEN_14906 = 14'h3a3a == index ? 14'h100 : _GEN_14905;
  wire [13:0] _GEN_14907 = 14'h3a3b == index ? 14'hb9 : _GEN_14906;
  wire [13:0] _GEN_14908 = 14'h3a3c == index ? 14'hb8 : _GEN_14907;
  wire [13:0] _GEN_14909 = 14'h3a3d == index ? 14'hb7 : _GEN_14908;
  wire [13:0] _GEN_14910 = 14'h3a3e == index ? 14'hb6 : _GEN_14909;
  wire [13:0] _GEN_14911 = 14'h3a3f == index ? 14'hb5 : _GEN_14910;
  wire [13:0] _GEN_14912 = 14'h3a40 == index ? 14'hb4 : _GEN_14911;
  wire [13:0] _GEN_14913 = 14'h3a41 == index ? 14'hb3 : _GEN_14912;
  wire [13:0] _GEN_14914 = 14'h3a42 == index ? 14'hb2 : _GEN_14913;
  wire [13:0] _GEN_14915 = 14'h3a43 == index ? 14'hb1 : _GEN_14914;
  wire [13:0] _GEN_14916 = 14'h3a44 == index ? 14'hb0 : _GEN_14915;
  wire [13:0] _GEN_14917 = 14'h3a45 == index ? 14'haf : _GEN_14916;
  wire [13:0] _GEN_14918 = 14'h3a46 == index ? 14'hae : _GEN_14917;
  wire [13:0] _GEN_14919 = 14'h3a47 == index ? 14'had : _GEN_14918;
  wire [13:0] _GEN_14920 = 14'h3a48 == index ? 14'hac : _GEN_14919;
  wire [13:0] _GEN_14921 = 14'h3a49 == index ? 14'hab : _GEN_14920;
  wire [13:0] _GEN_14922 = 14'h3a4a == index ? 14'haa : _GEN_14921;
  wire [13:0] _GEN_14923 = 14'h3a4b == index ? 14'ha9 : _GEN_14922;
  wire [13:0] _GEN_14924 = 14'h3a4c == index ? 14'ha8 : _GEN_14923;
  wire [13:0] _GEN_14925 = 14'h3a4d == index ? 14'ha7 : _GEN_14924;
  wire [13:0] _GEN_14926 = 14'h3a4e == index ? 14'ha6 : _GEN_14925;
  wire [13:0] _GEN_14927 = 14'h3a4f == index ? 14'ha5 : _GEN_14926;
  wire [13:0] _GEN_14928 = 14'h3a50 == index ? 14'ha4 : _GEN_14927;
  wire [13:0] _GEN_14929 = 14'h3a51 == index ? 14'ha3 : _GEN_14928;
  wire [13:0] _GEN_14930 = 14'h3a52 == index ? 14'ha2 : _GEN_14929;
  wire [13:0] _GEN_14931 = 14'h3a53 == index ? 14'ha1 : _GEN_14930;
  wire [13:0] _GEN_14932 = 14'h3a54 == index ? 14'ha0 : _GEN_14931;
  wire [13:0] _GEN_14933 = 14'h3a55 == index ? 14'h9f : _GEN_14932;
  wire [13:0] _GEN_14934 = 14'h3a56 == index ? 14'h9e : _GEN_14933;
  wire [13:0] _GEN_14935 = 14'h3a57 == index ? 14'h9d : _GEN_14934;
  wire [13:0] _GEN_14936 = 14'h3a58 == index ? 14'h9c : _GEN_14935;
  wire [13:0] _GEN_14937 = 14'h3a59 == index ? 14'h9b : _GEN_14936;
  wire [13:0] _GEN_14938 = 14'h3a5a == index ? 14'h9a : _GEN_14937;
  wire [13:0] _GEN_14939 = 14'h3a5b == index ? 14'h99 : _GEN_14938;
  wire [13:0] _GEN_14940 = 14'h3a5c == index ? 14'h98 : _GEN_14939;
  wire [13:0] _GEN_14941 = 14'h3a5d == index ? 14'h97 : _GEN_14940;
  wire [13:0] _GEN_14942 = 14'h3a5e == index ? 14'h96 : _GEN_14941;
  wire [13:0] _GEN_14943 = 14'h3a5f == index ? 14'h95 : _GEN_14942;
  wire [13:0] _GEN_14944 = 14'h3a60 == index ? 14'h94 : _GEN_14943;
  wire [13:0] _GEN_14945 = 14'h3a61 == index ? 14'h93 : _GEN_14944;
  wire [13:0] _GEN_14946 = 14'h3a62 == index ? 14'h92 : _GEN_14945;
  wire [13:0] _GEN_14947 = 14'h3a63 == index ? 14'h91 : _GEN_14946;
  wire [13:0] _GEN_14948 = 14'h3a64 == index ? 14'h90 : _GEN_14947;
  wire [13:0] _GEN_14949 = 14'h3a65 == index ? 14'h8f : _GEN_14948;
  wire [13:0] _GEN_14950 = 14'h3a66 == index ? 14'h8e : _GEN_14949;
  wire [13:0] _GEN_14951 = 14'h3a67 == index ? 14'h8d : _GEN_14950;
  wire [13:0] _GEN_14952 = 14'h3a68 == index ? 14'h8c : _GEN_14951;
  wire [13:0] _GEN_14953 = 14'h3a69 == index ? 14'h8b : _GEN_14952;
  wire [13:0] _GEN_14954 = 14'h3a6a == index ? 14'h8a : _GEN_14953;
  wire [13:0] _GEN_14955 = 14'h3a6b == index ? 14'h89 : _GEN_14954;
  wire [13:0] _GEN_14956 = 14'h3a6c == index ? 14'h88 : _GEN_14955;
  wire [13:0] _GEN_14957 = 14'h3a6d == index ? 14'h87 : _GEN_14956;
  wire [13:0] _GEN_14958 = 14'h3a6e == index ? 14'h86 : _GEN_14957;
  wire [13:0] _GEN_14959 = 14'h3a6f == index ? 14'h85 : _GEN_14958;
  wire [13:0] _GEN_14960 = 14'h3a70 == index ? 14'h84 : _GEN_14959;
  wire [13:0] _GEN_14961 = 14'h3a71 == index ? 14'h83 : _GEN_14960;
  wire [13:0] _GEN_14962 = 14'h3a72 == index ? 14'h82 : _GEN_14961;
  wire [13:0] _GEN_14963 = 14'h3a73 == index ? 14'h81 : _GEN_14962;
  wire [13:0] _GEN_14964 = 14'h3a74 == index ? 14'h80 : _GEN_14963;
  wire [13:0] _GEN_14965 = 14'h3a75 == index ? 14'h74 : _GEN_14964;
  wire [13:0] _GEN_14966 = 14'h3a76 == index ? 14'h74 : _GEN_14965;
  wire [13:0] _GEN_14967 = 14'h3a77 == index ? 14'h74 : _GEN_14966;
  wire [13:0] _GEN_14968 = 14'h3a78 == index ? 14'h74 : _GEN_14967;
  wire [13:0] _GEN_14969 = 14'h3a79 == index ? 14'h74 : _GEN_14968;
  wire [13:0] _GEN_14970 = 14'h3a7a == index ? 14'h74 : _GEN_14969;
  wire [13:0] _GEN_14971 = 14'h3a7b == index ? 14'h74 : _GEN_14970;
  wire [13:0] _GEN_14972 = 14'h3a7c == index ? 14'h74 : _GEN_14971;
  wire [13:0] _GEN_14973 = 14'h3a7d == index ? 14'h74 : _GEN_14972;
  wire [13:0] _GEN_14974 = 14'h3a7e == index ? 14'h74 : _GEN_14973;
  wire [13:0] _GEN_14975 = 14'h3a7f == index ? 14'h74 : _GEN_14974;
  wire [13:0] _GEN_14976 = 14'h3a80 == index ? 14'h0 : _GEN_14975;
  wire [13:0] _GEN_14977 = 14'h3a81 == index ? 14'h3a80 : _GEN_14976;
  wire [13:0] _GEN_14978 = 14'h3a82 == index ? 14'h1d01 : _GEN_14977;
  wire [13:0] _GEN_14979 = 14'h3a83 == index ? 14'h1380 : _GEN_14978;
  wire [13:0] _GEN_14980 = 14'h3a84 == index ? 14'he81 : _GEN_14979;
  wire [13:0] _GEN_14981 = 14'h3a85 == index ? 14'hb82 : _GEN_14980;
  wire [13:0] _GEN_14982 = 14'h3a86 == index ? 14'h983 : _GEN_14981;
  wire [13:0] _GEN_14983 = 14'h3a87 == index ? 14'h805 : _GEN_14982;
  wire [13:0] _GEN_14984 = 14'h3a88 == index ? 14'h705 : _GEN_14983;
  wire [13:0] _GEN_14985 = 14'h3a89 == index ? 14'h680 : _GEN_14984;
  wire [13:0] _GEN_14986 = 14'h3a8a == index ? 14'h587 : _GEN_14985;
  wire [13:0] _GEN_14987 = 14'h3a8b == index ? 14'h507 : _GEN_14986;
  wire [13:0] _GEN_14988 = 14'h3a8c == index ? 14'h489 : _GEN_14987;
  wire [13:0] _GEN_14989 = 14'h3a8d == index ? 14'h480 : _GEN_14988;
  wire [13:0] _GEN_14990 = 14'h3a8e == index ? 14'h405 : _GEN_14989;
  wire [13:0] _GEN_14991 = 14'h3a8f == index ? 14'h38c : _GEN_14990;
  wire [13:0] _GEN_14992 = 14'h3a90 == index ? 14'h385 : _GEN_14991;
  wire [13:0] _GEN_14993 = 14'h3a91 == index ? 14'h30f : _GEN_14992;
  wire [13:0] _GEN_14994 = 14'h3a92 == index ? 14'h309 : _GEN_14993;
  wire [13:0] _GEN_14995 = 14'h3a93 == index ? 14'h303 : _GEN_14994;
  wire [13:0] _GEN_14996 = 14'h3a94 == index ? 14'h291 : _GEN_14995;
  wire [13:0] _GEN_14997 = 14'h3a95 == index ? 14'h28c : _GEN_14996;
  wire [13:0] _GEN_14998 = 14'h3a96 == index ? 14'h287 : _GEN_14997;
  wire [13:0] _GEN_14999 = 14'h3a97 == index ? 14'h282 : _GEN_14998;
  wire [13:0] _GEN_15000 = 14'h3a98 == index ? 14'h215 : _GEN_14999;
  wire [13:0] _GEN_15001 = 14'h3a99 == index ? 14'h211 : _GEN_15000;
  wire [13:0] _GEN_15002 = 14'h3a9a == index ? 14'h20d : _GEN_15001;
  wire [13:0] _GEN_15003 = 14'h3a9b == index ? 14'h209 : _GEN_15002;
  wire [13:0] _GEN_15004 = 14'h3a9c == index ? 14'h205 : _GEN_15003;
  wire [13:0] _GEN_15005 = 14'h3a9d == index ? 14'h201 : _GEN_15004;
  wire [13:0] _GEN_15006 = 14'h3a9e == index ? 14'h19b : _GEN_15005;
  wire [13:0] _GEN_15007 = 14'h3a9f == index ? 14'h198 : _GEN_15006;
  wire [13:0] _GEN_15008 = 14'h3aa0 == index ? 14'h195 : _GEN_15007;
  wire [13:0] _GEN_15009 = 14'h3aa1 == index ? 14'h192 : _GEN_15008;
  wire [13:0] _GEN_15010 = 14'h3aa2 == index ? 14'h18f : _GEN_15009;
  wire [13:0] _GEN_15011 = 14'h3aa3 == index ? 14'h18c : _GEN_15010;
  wire [13:0] _GEN_15012 = 14'h3aa4 == index ? 14'h189 : _GEN_15011;
  wire [13:0] _GEN_15013 = 14'h3aa5 == index ? 14'h186 : _GEN_15012;
  wire [13:0] _GEN_15014 = 14'h3aa6 == index ? 14'h183 : _GEN_15013;
  wire [13:0] _GEN_15015 = 14'h3aa7 == index ? 14'h180 : _GEN_15014;
  wire [13:0] _GEN_15016 = 14'h3aa8 == index ? 14'h125 : _GEN_15015;
  wire [13:0] _GEN_15017 = 14'h3aa9 == index ? 14'h123 : _GEN_15016;
  wire [13:0] _GEN_15018 = 14'h3aaa == index ? 14'h121 : _GEN_15017;
  wire [13:0] _GEN_15019 = 14'h3aab == index ? 14'h11f : _GEN_15018;
  wire [13:0] _GEN_15020 = 14'h3aac == index ? 14'h11d : _GEN_15019;
  wire [13:0] _GEN_15021 = 14'h3aad == index ? 14'h11b : _GEN_15020;
  wire [13:0] _GEN_15022 = 14'h3aae == index ? 14'h119 : _GEN_15021;
  wire [13:0] _GEN_15023 = 14'h3aaf == index ? 14'h117 : _GEN_15022;
  wire [13:0] _GEN_15024 = 14'h3ab0 == index ? 14'h115 : _GEN_15023;
  wire [13:0] _GEN_15025 = 14'h3ab1 == index ? 14'h113 : _GEN_15024;
  wire [13:0] _GEN_15026 = 14'h3ab2 == index ? 14'h111 : _GEN_15025;
  wire [13:0] _GEN_15027 = 14'h3ab3 == index ? 14'h10f : _GEN_15026;
  wire [13:0] _GEN_15028 = 14'h3ab4 == index ? 14'h10d : _GEN_15027;
  wire [13:0] _GEN_15029 = 14'h3ab5 == index ? 14'h10b : _GEN_15028;
  wire [13:0] _GEN_15030 = 14'h3ab6 == index ? 14'h109 : _GEN_15029;
  wire [13:0] _GEN_15031 = 14'h3ab7 == index ? 14'h107 : _GEN_15030;
  wire [13:0] _GEN_15032 = 14'h3ab8 == index ? 14'h105 : _GEN_15031;
  wire [13:0] _GEN_15033 = 14'h3ab9 == index ? 14'h103 : _GEN_15032;
  wire [13:0] _GEN_15034 = 14'h3aba == index ? 14'h101 : _GEN_15033;
  wire [13:0] _GEN_15035 = 14'h3abb == index ? 14'hba : _GEN_15034;
  wire [13:0] _GEN_15036 = 14'h3abc == index ? 14'hb9 : _GEN_15035;
  wire [13:0] _GEN_15037 = 14'h3abd == index ? 14'hb8 : _GEN_15036;
  wire [13:0] _GEN_15038 = 14'h3abe == index ? 14'hb7 : _GEN_15037;
  wire [13:0] _GEN_15039 = 14'h3abf == index ? 14'hb6 : _GEN_15038;
  wire [13:0] _GEN_15040 = 14'h3ac0 == index ? 14'hb5 : _GEN_15039;
  wire [13:0] _GEN_15041 = 14'h3ac1 == index ? 14'hb4 : _GEN_15040;
  wire [13:0] _GEN_15042 = 14'h3ac2 == index ? 14'hb3 : _GEN_15041;
  wire [13:0] _GEN_15043 = 14'h3ac3 == index ? 14'hb2 : _GEN_15042;
  wire [13:0] _GEN_15044 = 14'h3ac4 == index ? 14'hb1 : _GEN_15043;
  wire [13:0] _GEN_15045 = 14'h3ac5 == index ? 14'hb0 : _GEN_15044;
  wire [13:0] _GEN_15046 = 14'h3ac6 == index ? 14'haf : _GEN_15045;
  wire [13:0] _GEN_15047 = 14'h3ac7 == index ? 14'hae : _GEN_15046;
  wire [13:0] _GEN_15048 = 14'h3ac8 == index ? 14'had : _GEN_15047;
  wire [13:0] _GEN_15049 = 14'h3ac9 == index ? 14'hac : _GEN_15048;
  wire [13:0] _GEN_15050 = 14'h3aca == index ? 14'hab : _GEN_15049;
  wire [13:0] _GEN_15051 = 14'h3acb == index ? 14'haa : _GEN_15050;
  wire [13:0] _GEN_15052 = 14'h3acc == index ? 14'ha9 : _GEN_15051;
  wire [13:0] _GEN_15053 = 14'h3acd == index ? 14'ha8 : _GEN_15052;
  wire [13:0] _GEN_15054 = 14'h3ace == index ? 14'ha7 : _GEN_15053;
  wire [13:0] _GEN_15055 = 14'h3acf == index ? 14'ha6 : _GEN_15054;
  wire [13:0] _GEN_15056 = 14'h3ad0 == index ? 14'ha5 : _GEN_15055;
  wire [13:0] _GEN_15057 = 14'h3ad1 == index ? 14'ha4 : _GEN_15056;
  wire [13:0] _GEN_15058 = 14'h3ad2 == index ? 14'ha3 : _GEN_15057;
  wire [13:0] _GEN_15059 = 14'h3ad3 == index ? 14'ha2 : _GEN_15058;
  wire [13:0] _GEN_15060 = 14'h3ad4 == index ? 14'ha1 : _GEN_15059;
  wire [13:0] _GEN_15061 = 14'h3ad5 == index ? 14'ha0 : _GEN_15060;
  wire [13:0] _GEN_15062 = 14'h3ad6 == index ? 14'h9f : _GEN_15061;
  wire [13:0] _GEN_15063 = 14'h3ad7 == index ? 14'h9e : _GEN_15062;
  wire [13:0] _GEN_15064 = 14'h3ad8 == index ? 14'h9d : _GEN_15063;
  wire [13:0] _GEN_15065 = 14'h3ad9 == index ? 14'h9c : _GEN_15064;
  wire [13:0] _GEN_15066 = 14'h3ada == index ? 14'h9b : _GEN_15065;
  wire [13:0] _GEN_15067 = 14'h3adb == index ? 14'h9a : _GEN_15066;
  wire [13:0] _GEN_15068 = 14'h3adc == index ? 14'h99 : _GEN_15067;
  wire [13:0] _GEN_15069 = 14'h3add == index ? 14'h98 : _GEN_15068;
  wire [13:0] _GEN_15070 = 14'h3ade == index ? 14'h97 : _GEN_15069;
  wire [13:0] _GEN_15071 = 14'h3adf == index ? 14'h96 : _GEN_15070;
  wire [13:0] _GEN_15072 = 14'h3ae0 == index ? 14'h95 : _GEN_15071;
  wire [13:0] _GEN_15073 = 14'h3ae1 == index ? 14'h94 : _GEN_15072;
  wire [13:0] _GEN_15074 = 14'h3ae2 == index ? 14'h93 : _GEN_15073;
  wire [13:0] _GEN_15075 = 14'h3ae3 == index ? 14'h92 : _GEN_15074;
  wire [13:0] _GEN_15076 = 14'h3ae4 == index ? 14'h91 : _GEN_15075;
  wire [13:0] _GEN_15077 = 14'h3ae5 == index ? 14'h90 : _GEN_15076;
  wire [13:0] _GEN_15078 = 14'h3ae6 == index ? 14'h8f : _GEN_15077;
  wire [13:0] _GEN_15079 = 14'h3ae7 == index ? 14'h8e : _GEN_15078;
  wire [13:0] _GEN_15080 = 14'h3ae8 == index ? 14'h8d : _GEN_15079;
  wire [13:0] _GEN_15081 = 14'h3ae9 == index ? 14'h8c : _GEN_15080;
  wire [13:0] _GEN_15082 = 14'h3aea == index ? 14'h8b : _GEN_15081;
  wire [13:0] _GEN_15083 = 14'h3aeb == index ? 14'h8a : _GEN_15082;
  wire [13:0] _GEN_15084 = 14'h3aec == index ? 14'h89 : _GEN_15083;
  wire [13:0] _GEN_15085 = 14'h3aed == index ? 14'h88 : _GEN_15084;
  wire [13:0] _GEN_15086 = 14'h3aee == index ? 14'h87 : _GEN_15085;
  wire [13:0] _GEN_15087 = 14'h3aef == index ? 14'h86 : _GEN_15086;
  wire [13:0] _GEN_15088 = 14'h3af0 == index ? 14'h85 : _GEN_15087;
  wire [13:0] _GEN_15089 = 14'h3af1 == index ? 14'h84 : _GEN_15088;
  wire [13:0] _GEN_15090 = 14'h3af2 == index ? 14'h83 : _GEN_15089;
  wire [13:0] _GEN_15091 = 14'h3af3 == index ? 14'h82 : _GEN_15090;
  wire [13:0] _GEN_15092 = 14'h3af4 == index ? 14'h81 : _GEN_15091;
  wire [13:0] _GEN_15093 = 14'h3af5 == index ? 14'h80 : _GEN_15092;
  wire [13:0] _GEN_15094 = 14'h3af6 == index ? 14'h75 : _GEN_15093;
  wire [13:0] _GEN_15095 = 14'h3af7 == index ? 14'h75 : _GEN_15094;
  wire [13:0] _GEN_15096 = 14'h3af8 == index ? 14'h75 : _GEN_15095;
  wire [13:0] _GEN_15097 = 14'h3af9 == index ? 14'h75 : _GEN_15096;
  wire [13:0] _GEN_15098 = 14'h3afa == index ? 14'h75 : _GEN_15097;
  wire [13:0] _GEN_15099 = 14'h3afb == index ? 14'h75 : _GEN_15098;
  wire [13:0] _GEN_15100 = 14'h3afc == index ? 14'h75 : _GEN_15099;
  wire [13:0] _GEN_15101 = 14'h3afd == index ? 14'h75 : _GEN_15100;
  wire [13:0] _GEN_15102 = 14'h3afe == index ? 14'h75 : _GEN_15101;
  wire [13:0] _GEN_15103 = 14'h3aff == index ? 14'h75 : _GEN_15102;
  wire [13:0] _GEN_15104 = 14'h3b00 == index ? 14'h0 : _GEN_15103;
  wire [13:0] _GEN_15105 = 14'h3b01 == index ? 14'h3b00 : _GEN_15104;
  wire [13:0] _GEN_15106 = 14'h3b02 == index ? 14'h1d80 : _GEN_15105;
  wire [13:0] _GEN_15107 = 14'h3b03 == index ? 14'h1381 : _GEN_15106;
  wire [13:0] _GEN_15108 = 14'h3b04 == index ? 14'he82 : _GEN_15107;
  wire [13:0] _GEN_15109 = 14'h3b05 == index ? 14'hb83 : _GEN_15108;
  wire [13:0] _GEN_15110 = 14'h3b06 == index ? 14'h984 : _GEN_15109;
  wire [13:0] _GEN_15111 = 14'h3b07 == index ? 14'h806 : _GEN_15110;
  wire [13:0] _GEN_15112 = 14'h3b08 == index ? 14'h706 : _GEN_15111;
  wire [13:0] _GEN_15113 = 14'h3b09 == index ? 14'h681 : _GEN_15112;
  wire [13:0] _GEN_15114 = 14'h3b0a == index ? 14'h588 : _GEN_15113;
  wire [13:0] _GEN_15115 = 14'h3b0b == index ? 14'h508 : _GEN_15114;
  wire [13:0] _GEN_15116 = 14'h3b0c == index ? 14'h48a : _GEN_15115;
  wire [13:0] _GEN_15117 = 14'h3b0d == index ? 14'h481 : _GEN_15116;
  wire [13:0] _GEN_15118 = 14'h3b0e == index ? 14'h406 : _GEN_15117;
  wire [13:0] _GEN_15119 = 14'h3b0f == index ? 14'h38d : _GEN_15118;
  wire [13:0] _GEN_15120 = 14'h3b10 == index ? 14'h386 : _GEN_15119;
  wire [13:0] _GEN_15121 = 14'h3b11 == index ? 14'h310 : _GEN_15120;
  wire [13:0] _GEN_15122 = 14'h3b12 == index ? 14'h30a : _GEN_15121;
  wire [13:0] _GEN_15123 = 14'h3b13 == index ? 14'h304 : _GEN_15122;
  wire [13:0] _GEN_15124 = 14'h3b14 == index ? 14'h292 : _GEN_15123;
  wire [13:0] _GEN_15125 = 14'h3b15 == index ? 14'h28d : _GEN_15124;
  wire [13:0] _GEN_15126 = 14'h3b16 == index ? 14'h288 : _GEN_15125;
  wire [13:0] _GEN_15127 = 14'h3b17 == index ? 14'h283 : _GEN_15126;
  wire [13:0] _GEN_15128 = 14'h3b18 == index ? 14'h216 : _GEN_15127;
  wire [13:0] _GEN_15129 = 14'h3b19 == index ? 14'h212 : _GEN_15128;
  wire [13:0] _GEN_15130 = 14'h3b1a == index ? 14'h20e : _GEN_15129;
  wire [13:0] _GEN_15131 = 14'h3b1b == index ? 14'h20a : _GEN_15130;
  wire [13:0] _GEN_15132 = 14'h3b1c == index ? 14'h206 : _GEN_15131;
  wire [13:0] _GEN_15133 = 14'h3b1d == index ? 14'h202 : _GEN_15132;
  wire [13:0] _GEN_15134 = 14'h3b1e == index ? 14'h19c : _GEN_15133;
  wire [13:0] _GEN_15135 = 14'h3b1f == index ? 14'h199 : _GEN_15134;
  wire [13:0] _GEN_15136 = 14'h3b20 == index ? 14'h196 : _GEN_15135;
  wire [13:0] _GEN_15137 = 14'h3b21 == index ? 14'h193 : _GEN_15136;
  wire [13:0] _GEN_15138 = 14'h3b22 == index ? 14'h190 : _GEN_15137;
  wire [13:0] _GEN_15139 = 14'h3b23 == index ? 14'h18d : _GEN_15138;
  wire [13:0] _GEN_15140 = 14'h3b24 == index ? 14'h18a : _GEN_15139;
  wire [13:0] _GEN_15141 = 14'h3b25 == index ? 14'h187 : _GEN_15140;
  wire [13:0] _GEN_15142 = 14'h3b26 == index ? 14'h184 : _GEN_15141;
  wire [13:0] _GEN_15143 = 14'h3b27 == index ? 14'h181 : _GEN_15142;
  wire [13:0] _GEN_15144 = 14'h3b28 == index ? 14'h126 : _GEN_15143;
  wire [13:0] _GEN_15145 = 14'h3b29 == index ? 14'h124 : _GEN_15144;
  wire [13:0] _GEN_15146 = 14'h3b2a == index ? 14'h122 : _GEN_15145;
  wire [13:0] _GEN_15147 = 14'h3b2b == index ? 14'h120 : _GEN_15146;
  wire [13:0] _GEN_15148 = 14'h3b2c == index ? 14'h11e : _GEN_15147;
  wire [13:0] _GEN_15149 = 14'h3b2d == index ? 14'h11c : _GEN_15148;
  wire [13:0] _GEN_15150 = 14'h3b2e == index ? 14'h11a : _GEN_15149;
  wire [13:0] _GEN_15151 = 14'h3b2f == index ? 14'h118 : _GEN_15150;
  wire [13:0] _GEN_15152 = 14'h3b30 == index ? 14'h116 : _GEN_15151;
  wire [13:0] _GEN_15153 = 14'h3b31 == index ? 14'h114 : _GEN_15152;
  wire [13:0] _GEN_15154 = 14'h3b32 == index ? 14'h112 : _GEN_15153;
  wire [13:0] _GEN_15155 = 14'h3b33 == index ? 14'h110 : _GEN_15154;
  wire [13:0] _GEN_15156 = 14'h3b34 == index ? 14'h10e : _GEN_15155;
  wire [13:0] _GEN_15157 = 14'h3b35 == index ? 14'h10c : _GEN_15156;
  wire [13:0] _GEN_15158 = 14'h3b36 == index ? 14'h10a : _GEN_15157;
  wire [13:0] _GEN_15159 = 14'h3b37 == index ? 14'h108 : _GEN_15158;
  wire [13:0] _GEN_15160 = 14'h3b38 == index ? 14'h106 : _GEN_15159;
  wire [13:0] _GEN_15161 = 14'h3b39 == index ? 14'h104 : _GEN_15160;
  wire [13:0] _GEN_15162 = 14'h3b3a == index ? 14'h102 : _GEN_15161;
  wire [13:0] _GEN_15163 = 14'h3b3b == index ? 14'h100 : _GEN_15162;
  wire [13:0] _GEN_15164 = 14'h3b3c == index ? 14'hba : _GEN_15163;
  wire [13:0] _GEN_15165 = 14'h3b3d == index ? 14'hb9 : _GEN_15164;
  wire [13:0] _GEN_15166 = 14'h3b3e == index ? 14'hb8 : _GEN_15165;
  wire [13:0] _GEN_15167 = 14'h3b3f == index ? 14'hb7 : _GEN_15166;
  wire [13:0] _GEN_15168 = 14'h3b40 == index ? 14'hb6 : _GEN_15167;
  wire [13:0] _GEN_15169 = 14'h3b41 == index ? 14'hb5 : _GEN_15168;
  wire [13:0] _GEN_15170 = 14'h3b42 == index ? 14'hb4 : _GEN_15169;
  wire [13:0] _GEN_15171 = 14'h3b43 == index ? 14'hb3 : _GEN_15170;
  wire [13:0] _GEN_15172 = 14'h3b44 == index ? 14'hb2 : _GEN_15171;
  wire [13:0] _GEN_15173 = 14'h3b45 == index ? 14'hb1 : _GEN_15172;
  wire [13:0] _GEN_15174 = 14'h3b46 == index ? 14'hb0 : _GEN_15173;
  wire [13:0] _GEN_15175 = 14'h3b47 == index ? 14'haf : _GEN_15174;
  wire [13:0] _GEN_15176 = 14'h3b48 == index ? 14'hae : _GEN_15175;
  wire [13:0] _GEN_15177 = 14'h3b49 == index ? 14'had : _GEN_15176;
  wire [13:0] _GEN_15178 = 14'h3b4a == index ? 14'hac : _GEN_15177;
  wire [13:0] _GEN_15179 = 14'h3b4b == index ? 14'hab : _GEN_15178;
  wire [13:0] _GEN_15180 = 14'h3b4c == index ? 14'haa : _GEN_15179;
  wire [13:0] _GEN_15181 = 14'h3b4d == index ? 14'ha9 : _GEN_15180;
  wire [13:0] _GEN_15182 = 14'h3b4e == index ? 14'ha8 : _GEN_15181;
  wire [13:0] _GEN_15183 = 14'h3b4f == index ? 14'ha7 : _GEN_15182;
  wire [13:0] _GEN_15184 = 14'h3b50 == index ? 14'ha6 : _GEN_15183;
  wire [13:0] _GEN_15185 = 14'h3b51 == index ? 14'ha5 : _GEN_15184;
  wire [13:0] _GEN_15186 = 14'h3b52 == index ? 14'ha4 : _GEN_15185;
  wire [13:0] _GEN_15187 = 14'h3b53 == index ? 14'ha3 : _GEN_15186;
  wire [13:0] _GEN_15188 = 14'h3b54 == index ? 14'ha2 : _GEN_15187;
  wire [13:0] _GEN_15189 = 14'h3b55 == index ? 14'ha1 : _GEN_15188;
  wire [13:0] _GEN_15190 = 14'h3b56 == index ? 14'ha0 : _GEN_15189;
  wire [13:0] _GEN_15191 = 14'h3b57 == index ? 14'h9f : _GEN_15190;
  wire [13:0] _GEN_15192 = 14'h3b58 == index ? 14'h9e : _GEN_15191;
  wire [13:0] _GEN_15193 = 14'h3b59 == index ? 14'h9d : _GEN_15192;
  wire [13:0] _GEN_15194 = 14'h3b5a == index ? 14'h9c : _GEN_15193;
  wire [13:0] _GEN_15195 = 14'h3b5b == index ? 14'h9b : _GEN_15194;
  wire [13:0] _GEN_15196 = 14'h3b5c == index ? 14'h9a : _GEN_15195;
  wire [13:0] _GEN_15197 = 14'h3b5d == index ? 14'h99 : _GEN_15196;
  wire [13:0] _GEN_15198 = 14'h3b5e == index ? 14'h98 : _GEN_15197;
  wire [13:0] _GEN_15199 = 14'h3b5f == index ? 14'h97 : _GEN_15198;
  wire [13:0] _GEN_15200 = 14'h3b60 == index ? 14'h96 : _GEN_15199;
  wire [13:0] _GEN_15201 = 14'h3b61 == index ? 14'h95 : _GEN_15200;
  wire [13:0] _GEN_15202 = 14'h3b62 == index ? 14'h94 : _GEN_15201;
  wire [13:0] _GEN_15203 = 14'h3b63 == index ? 14'h93 : _GEN_15202;
  wire [13:0] _GEN_15204 = 14'h3b64 == index ? 14'h92 : _GEN_15203;
  wire [13:0] _GEN_15205 = 14'h3b65 == index ? 14'h91 : _GEN_15204;
  wire [13:0] _GEN_15206 = 14'h3b66 == index ? 14'h90 : _GEN_15205;
  wire [13:0] _GEN_15207 = 14'h3b67 == index ? 14'h8f : _GEN_15206;
  wire [13:0] _GEN_15208 = 14'h3b68 == index ? 14'h8e : _GEN_15207;
  wire [13:0] _GEN_15209 = 14'h3b69 == index ? 14'h8d : _GEN_15208;
  wire [13:0] _GEN_15210 = 14'h3b6a == index ? 14'h8c : _GEN_15209;
  wire [13:0] _GEN_15211 = 14'h3b6b == index ? 14'h8b : _GEN_15210;
  wire [13:0] _GEN_15212 = 14'h3b6c == index ? 14'h8a : _GEN_15211;
  wire [13:0] _GEN_15213 = 14'h3b6d == index ? 14'h89 : _GEN_15212;
  wire [13:0] _GEN_15214 = 14'h3b6e == index ? 14'h88 : _GEN_15213;
  wire [13:0] _GEN_15215 = 14'h3b6f == index ? 14'h87 : _GEN_15214;
  wire [13:0] _GEN_15216 = 14'h3b70 == index ? 14'h86 : _GEN_15215;
  wire [13:0] _GEN_15217 = 14'h3b71 == index ? 14'h85 : _GEN_15216;
  wire [13:0] _GEN_15218 = 14'h3b72 == index ? 14'h84 : _GEN_15217;
  wire [13:0] _GEN_15219 = 14'h3b73 == index ? 14'h83 : _GEN_15218;
  wire [13:0] _GEN_15220 = 14'h3b74 == index ? 14'h82 : _GEN_15219;
  wire [13:0] _GEN_15221 = 14'h3b75 == index ? 14'h81 : _GEN_15220;
  wire [13:0] _GEN_15222 = 14'h3b76 == index ? 14'h80 : _GEN_15221;
  wire [13:0] _GEN_15223 = 14'h3b77 == index ? 14'h76 : _GEN_15222;
  wire [13:0] _GEN_15224 = 14'h3b78 == index ? 14'h76 : _GEN_15223;
  wire [13:0] _GEN_15225 = 14'h3b79 == index ? 14'h76 : _GEN_15224;
  wire [13:0] _GEN_15226 = 14'h3b7a == index ? 14'h76 : _GEN_15225;
  wire [13:0] _GEN_15227 = 14'h3b7b == index ? 14'h76 : _GEN_15226;
  wire [13:0] _GEN_15228 = 14'h3b7c == index ? 14'h76 : _GEN_15227;
  wire [13:0] _GEN_15229 = 14'h3b7d == index ? 14'h76 : _GEN_15228;
  wire [13:0] _GEN_15230 = 14'h3b7e == index ? 14'h76 : _GEN_15229;
  wire [13:0] _GEN_15231 = 14'h3b7f == index ? 14'h76 : _GEN_15230;
  wire [13:0] _GEN_15232 = 14'h3b80 == index ? 14'h0 : _GEN_15231;
  wire [13:0] _GEN_15233 = 14'h3b81 == index ? 14'h3b80 : _GEN_15232;
  wire [13:0] _GEN_15234 = 14'h3b82 == index ? 14'h1d81 : _GEN_15233;
  wire [13:0] _GEN_15235 = 14'h3b83 == index ? 14'h1382 : _GEN_15234;
  wire [13:0] _GEN_15236 = 14'h3b84 == index ? 14'he83 : _GEN_15235;
  wire [13:0] _GEN_15237 = 14'h3b85 == index ? 14'hb84 : _GEN_15236;
  wire [13:0] _GEN_15238 = 14'h3b86 == index ? 14'h985 : _GEN_15237;
  wire [13:0] _GEN_15239 = 14'h3b87 == index ? 14'h880 : _GEN_15238;
  wire [13:0] _GEN_15240 = 14'h3b88 == index ? 14'h707 : _GEN_15239;
  wire [13:0] _GEN_15241 = 14'h3b89 == index ? 14'h682 : _GEN_15240;
  wire [13:0] _GEN_15242 = 14'h3b8a == index ? 14'h589 : _GEN_15241;
  wire [13:0] _GEN_15243 = 14'h3b8b == index ? 14'h509 : _GEN_15242;
  wire [13:0] _GEN_15244 = 14'h3b8c == index ? 14'h48b : _GEN_15243;
  wire [13:0] _GEN_15245 = 14'h3b8d == index ? 14'h482 : _GEN_15244;
  wire [13:0] _GEN_15246 = 14'h3b8e == index ? 14'h407 : _GEN_15245;
  wire [13:0] _GEN_15247 = 14'h3b8f == index ? 14'h38e : _GEN_15246;
  wire [13:0] _GEN_15248 = 14'h3b90 == index ? 14'h387 : _GEN_15247;
  wire [13:0] _GEN_15249 = 14'h3b91 == index ? 14'h380 : _GEN_15248;
  wire [13:0] _GEN_15250 = 14'h3b92 == index ? 14'h30b : _GEN_15249;
  wire [13:0] _GEN_15251 = 14'h3b93 == index ? 14'h305 : _GEN_15250;
  wire [13:0] _GEN_15252 = 14'h3b94 == index ? 14'h293 : _GEN_15251;
  wire [13:0] _GEN_15253 = 14'h3b95 == index ? 14'h28e : _GEN_15252;
  wire [13:0] _GEN_15254 = 14'h3b96 == index ? 14'h289 : _GEN_15253;
  wire [13:0] _GEN_15255 = 14'h3b97 == index ? 14'h284 : _GEN_15254;
  wire [13:0] _GEN_15256 = 14'h3b98 == index ? 14'h217 : _GEN_15255;
  wire [13:0] _GEN_15257 = 14'h3b99 == index ? 14'h213 : _GEN_15256;
  wire [13:0] _GEN_15258 = 14'h3b9a == index ? 14'h20f : _GEN_15257;
  wire [13:0] _GEN_15259 = 14'h3b9b == index ? 14'h20b : _GEN_15258;
  wire [13:0] _GEN_15260 = 14'h3b9c == index ? 14'h207 : _GEN_15259;
  wire [13:0] _GEN_15261 = 14'h3b9d == index ? 14'h203 : _GEN_15260;
  wire [13:0] _GEN_15262 = 14'h3b9e == index ? 14'h19d : _GEN_15261;
  wire [13:0] _GEN_15263 = 14'h3b9f == index ? 14'h19a : _GEN_15262;
  wire [13:0] _GEN_15264 = 14'h3ba0 == index ? 14'h197 : _GEN_15263;
  wire [13:0] _GEN_15265 = 14'h3ba1 == index ? 14'h194 : _GEN_15264;
  wire [13:0] _GEN_15266 = 14'h3ba2 == index ? 14'h191 : _GEN_15265;
  wire [13:0] _GEN_15267 = 14'h3ba3 == index ? 14'h18e : _GEN_15266;
  wire [13:0] _GEN_15268 = 14'h3ba4 == index ? 14'h18b : _GEN_15267;
  wire [13:0] _GEN_15269 = 14'h3ba5 == index ? 14'h188 : _GEN_15268;
  wire [13:0] _GEN_15270 = 14'h3ba6 == index ? 14'h185 : _GEN_15269;
  wire [13:0] _GEN_15271 = 14'h3ba7 == index ? 14'h182 : _GEN_15270;
  wire [13:0] _GEN_15272 = 14'h3ba8 == index ? 14'h127 : _GEN_15271;
  wire [13:0] _GEN_15273 = 14'h3ba9 == index ? 14'h125 : _GEN_15272;
  wire [13:0] _GEN_15274 = 14'h3baa == index ? 14'h123 : _GEN_15273;
  wire [13:0] _GEN_15275 = 14'h3bab == index ? 14'h121 : _GEN_15274;
  wire [13:0] _GEN_15276 = 14'h3bac == index ? 14'h11f : _GEN_15275;
  wire [13:0] _GEN_15277 = 14'h3bad == index ? 14'h11d : _GEN_15276;
  wire [13:0] _GEN_15278 = 14'h3bae == index ? 14'h11b : _GEN_15277;
  wire [13:0] _GEN_15279 = 14'h3baf == index ? 14'h119 : _GEN_15278;
  wire [13:0] _GEN_15280 = 14'h3bb0 == index ? 14'h117 : _GEN_15279;
  wire [13:0] _GEN_15281 = 14'h3bb1 == index ? 14'h115 : _GEN_15280;
  wire [13:0] _GEN_15282 = 14'h3bb2 == index ? 14'h113 : _GEN_15281;
  wire [13:0] _GEN_15283 = 14'h3bb3 == index ? 14'h111 : _GEN_15282;
  wire [13:0] _GEN_15284 = 14'h3bb4 == index ? 14'h10f : _GEN_15283;
  wire [13:0] _GEN_15285 = 14'h3bb5 == index ? 14'h10d : _GEN_15284;
  wire [13:0] _GEN_15286 = 14'h3bb6 == index ? 14'h10b : _GEN_15285;
  wire [13:0] _GEN_15287 = 14'h3bb7 == index ? 14'h109 : _GEN_15286;
  wire [13:0] _GEN_15288 = 14'h3bb8 == index ? 14'h107 : _GEN_15287;
  wire [13:0] _GEN_15289 = 14'h3bb9 == index ? 14'h105 : _GEN_15288;
  wire [13:0] _GEN_15290 = 14'h3bba == index ? 14'h103 : _GEN_15289;
  wire [13:0] _GEN_15291 = 14'h3bbb == index ? 14'h101 : _GEN_15290;
  wire [13:0] _GEN_15292 = 14'h3bbc == index ? 14'hbb : _GEN_15291;
  wire [13:0] _GEN_15293 = 14'h3bbd == index ? 14'hba : _GEN_15292;
  wire [13:0] _GEN_15294 = 14'h3bbe == index ? 14'hb9 : _GEN_15293;
  wire [13:0] _GEN_15295 = 14'h3bbf == index ? 14'hb8 : _GEN_15294;
  wire [13:0] _GEN_15296 = 14'h3bc0 == index ? 14'hb7 : _GEN_15295;
  wire [13:0] _GEN_15297 = 14'h3bc1 == index ? 14'hb6 : _GEN_15296;
  wire [13:0] _GEN_15298 = 14'h3bc2 == index ? 14'hb5 : _GEN_15297;
  wire [13:0] _GEN_15299 = 14'h3bc3 == index ? 14'hb4 : _GEN_15298;
  wire [13:0] _GEN_15300 = 14'h3bc4 == index ? 14'hb3 : _GEN_15299;
  wire [13:0] _GEN_15301 = 14'h3bc5 == index ? 14'hb2 : _GEN_15300;
  wire [13:0] _GEN_15302 = 14'h3bc6 == index ? 14'hb1 : _GEN_15301;
  wire [13:0] _GEN_15303 = 14'h3bc7 == index ? 14'hb0 : _GEN_15302;
  wire [13:0] _GEN_15304 = 14'h3bc8 == index ? 14'haf : _GEN_15303;
  wire [13:0] _GEN_15305 = 14'h3bc9 == index ? 14'hae : _GEN_15304;
  wire [13:0] _GEN_15306 = 14'h3bca == index ? 14'had : _GEN_15305;
  wire [13:0] _GEN_15307 = 14'h3bcb == index ? 14'hac : _GEN_15306;
  wire [13:0] _GEN_15308 = 14'h3bcc == index ? 14'hab : _GEN_15307;
  wire [13:0] _GEN_15309 = 14'h3bcd == index ? 14'haa : _GEN_15308;
  wire [13:0] _GEN_15310 = 14'h3bce == index ? 14'ha9 : _GEN_15309;
  wire [13:0] _GEN_15311 = 14'h3bcf == index ? 14'ha8 : _GEN_15310;
  wire [13:0] _GEN_15312 = 14'h3bd0 == index ? 14'ha7 : _GEN_15311;
  wire [13:0] _GEN_15313 = 14'h3bd1 == index ? 14'ha6 : _GEN_15312;
  wire [13:0] _GEN_15314 = 14'h3bd2 == index ? 14'ha5 : _GEN_15313;
  wire [13:0] _GEN_15315 = 14'h3bd3 == index ? 14'ha4 : _GEN_15314;
  wire [13:0] _GEN_15316 = 14'h3bd4 == index ? 14'ha3 : _GEN_15315;
  wire [13:0] _GEN_15317 = 14'h3bd5 == index ? 14'ha2 : _GEN_15316;
  wire [13:0] _GEN_15318 = 14'h3bd6 == index ? 14'ha1 : _GEN_15317;
  wire [13:0] _GEN_15319 = 14'h3bd7 == index ? 14'ha0 : _GEN_15318;
  wire [13:0] _GEN_15320 = 14'h3bd8 == index ? 14'h9f : _GEN_15319;
  wire [13:0] _GEN_15321 = 14'h3bd9 == index ? 14'h9e : _GEN_15320;
  wire [13:0] _GEN_15322 = 14'h3bda == index ? 14'h9d : _GEN_15321;
  wire [13:0] _GEN_15323 = 14'h3bdb == index ? 14'h9c : _GEN_15322;
  wire [13:0] _GEN_15324 = 14'h3bdc == index ? 14'h9b : _GEN_15323;
  wire [13:0] _GEN_15325 = 14'h3bdd == index ? 14'h9a : _GEN_15324;
  wire [13:0] _GEN_15326 = 14'h3bde == index ? 14'h99 : _GEN_15325;
  wire [13:0] _GEN_15327 = 14'h3bdf == index ? 14'h98 : _GEN_15326;
  wire [13:0] _GEN_15328 = 14'h3be0 == index ? 14'h97 : _GEN_15327;
  wire [13:0] _GEN_15329 = 14'h3be1 == index ? 14'h96 : _GEN_15328;
  wire [13:0] _GEN_15330 = 14'h3be2 == index ? 14'h95 : _GEN_15329;
  wire [13:0] _GEN_15331 = 14'h3be3 == index ? 14'h94 : _GEN_15330;
  wire [13:0] _GEN_15332 = 14'h3be4 == index ? 14'h93 : _GEN_15331;
  wire [13:0] _GEN_15333 = 14'h3be5 == index ? 14'h92 : _GEN_15332;
  wire [13:0] _GEN_15334 = 14'h3be6 == index ? 14'h91 : _GEN_15333;
  wire [13:0] _GEN_15335 = 14'h3be7 == index ? 14'h90 : _GEN_15334;
  wire [13:0] _GEN_15336 = 14'h3be8 == index ? 14'h8f : _GEN_15335;
  wire [13:0] _GEN_15337 = 14'h3be9 == index ? 14'h8e : _GEN_15336;
  wire [13:0] _GEN_15338 = 14'h3bea == index ? 14'h8d : _GEN_15337;
  wire [13:0] _GEN_15339 = 14'h3beb == index ? 14'h8c : _GEN_15338;
  wire [13:0] _GEN_15340 = 14'h3bec == index ? 14'h8b : _GEN_15339;
  wire [13:0] _GEN_15341 = 14'h3bed == index ? 14'h8a : _GEN_15340;
  wire [13:0] _GEN_15342 = 14'h3bee == index ? 14'h89 : _GEN_15341;
  wire [13:0] _GEN_15343 = 14'h3bef == index ? 14'h88 : _GEN_15342;
  wire [13:0] _GEN_15344 = 14'h3bf0 == index ? 14'h87 : _GEN_15343;
  wire [13:0] _GEN_15345 = 14'h3bf1 == index ? 14'h86 : _GEN_15344;
  wire [13:0] _GEN_15346 = 14'h3bf2 == index ? 14'h85 : _GEN_15345;
  wire [13:0] _GEN_15347 = 14'h3bf3 == index ? 14'h84 : _GEN_15346;
  wire [13:0] _GEN_15348 = 14'h3bf4 == index ? 14'h83 : _GEN_15347;
  wire [13:0] _GEN_15349 = 14'h3bf5 == index ? 14'h82 : _GEN_15348;
  wire [13:0] _GEN_15350 = 14'h3bf6 == index ? 14'h81 : _GEN_15349;
  wire [13:0] _GEN_15351 = 14'h3bf7 == index ? 14'h80 : _GEN_15350;
  wire [13:0] _GEN_15352 = 14'h3bf8 == index ? 14'h77 : _GEN_15351;
  wire [13:0] _GEN_15353 = 14'h3bf9 == index ? 14'h77 : _GEN_15352;
  wire [13:0] _GEN_15354 = 14'h3bfa == index ? 14'h77 : _GEN_15353;
  wire [13:0] _GEN_15355 = 14'h3bfb == index ? 14'h77 : _GEN_15354;
  wire [13:0] _GEN_15356 = 14'h3bfc == index ? 14'h77 : _GEN_15355;
  wire [13:0] _GEN_15357 = 14'h3bfd == index ? 14'h77 : _GEN_15356;
  wire [13:0] _GEN_15358 = 14'h3bfe == index ? 14'h77 : _GEN_15357;
  wire [13:0] _GEN_15359 = 14'h3bff == index ? 14'h77 : _GEN_15358;
  wire [13:0] _GEN_15360 = 14'h3c00 == index ? 14'h0 : _GEN_15359;
  wire [13:0] _GEN_15361 = 14'h3c01 == index ? 14'h3c00 : _GEN_15360;
  wire [13:0] _GEN_15362 = 14'h3c02 == index ? 14'h1e00 : _GEN_15361;
  wire [13:0] _GEN_15363 = 14'h3c03 == index ? 14'h1400 : _GEN_15362;
  wire [13:0] _GEN_15364 = 14'h3c04 == index ? 14'hf00 : _GEN_15363;
  wire [13:0] _GEN_15365 = 14'h3c05 == index ? 14'hc00 : _GEN_15364;
  wire [13:0] _GEN_15366 = 14'h3c06 == index ? 14'ha00 : _GEN_15365;
  wire [13:0] _GEN_15367 = 14'h3c07 == index ? 14'h881 : _GEN_15366;
  wire [13:0] _GEN_15368 = 14'h3c08 == index ? 14'h780 : _GEN_15367;
  wire [13:0] _GEN_15369 = 14'h3c09 == index ? 14'h683 : _GEN_15368;
  wire [13:0] _GEN_15370 = 14'h3c0a == index ? 14'h600 : _GEN_15369;
  wire [13:0] _GEN_15371 = 14'h3c0b == index ? 14'h50a : _GEN_15370;
  wire [13:0] _GEN_15372 = 14'h3c0c == index ? 14'h500 : _GEN_15371;
  wire [13:0] _GEN_15373 = 14'h3c0d == index ? 14'h483 : _GEN_15372;
  wire [13:0] _GEN_15374 = 14'h3c0e == index ? 14'h408 : _GEN_15373;
  wire [13:0] _GEN_15375 = 14'h3c0f == index ? 14'h400 : _GEN_15374;
  wire [13:0] _GEN_15376 = 14'h3c10 == index ? 14'h388 : _GEN_15375;
  wire [13:0] _GEN_15377 = 14'h3c11 == index ? 14'h381 : _GEN_15376;
  wire [13:0] _GEN_15378 = 14'h3c12 == index ? 14'h30c : _GEN_15377;
  wire [13:0] _GEN_15379 = 14'h3c13 == index ? 14'h306 : _GEN_15378;
  wire [13:0] _GEN_15380 = 14'h3c14 == index ? 14'h300 : _GEN_15379;
  wire [13:0] _GEN_15381 = 14'h3c15 == index ? 14'h28f : _GEN_15380;
  wire [13:0] _GEN_15382 = 14'h3c16 == index ? 14'h28a : _GEN_15381;
  wire [13:0] _GEN_15383 = 14'h3c17 == index ? 14'h285 : _GEN_15382;
  wire [13:0] _GEN_15384 = 14'h3c18 == index ? 14'h280 : _GEN_15383;
  wire [13:0] _GEN_15385 = 14'h3c19 == index ? 14'h214 : _GEN_15384;
  wire [13:0] _GEN_15386 = 14'h3c1a == index ? 14'h210 : _GEN_15385;
  wire [13:0] _GEN_15387 = 14'h3c1b == index ? 14'h20c : _GEN_15386;
  wire [13:0] _GEN_15388 = 14'h3c1c == index ? 14'h208 : _GEN_15387;
  wire [13:0] _GEN_15389 = 14'h3c1d == index ? 14'h204 : _GEN_15388;
  wire [13:0] _GEN_15390 = 14'h3c1e == index ? 14'h200 : _GEN_15389;
  wire [13:0] _GEN_15391 = 14'h3c1f == index ? 14'h19b : _GEN_15390;
  wire [13:0] _GEN_15392 = 14'h3c20 == index ? 14'h198 : _GEN_15391;
  wire [13:0] _GEN_15393 = 14'h3c21 == index ? 14'h195 : _GEN_15392;
  wire [13:0] _GEN_15394 = 14'h3c22 == index ? 14'h192 : _GEN_15393;
  wire [13:0] _GEN_15395 = 14'h3c23 == index ? 14'h18f : _GEN_15394;
  wire [13:0] _GEN_15396 = 14'h3c24 == index ? 14'h18c : _GEN_15395;
  wire [13:0] _GEN_15397 = 14'h3c25 == index ? 14'h189 : _GEN_15396;
  wire [13:0] _GEN_15398 = 14'h3c26 == index ? 14'h186 : _GEN_15397;
  wire [13:0] _GEN_15399 = 14'h3c27 == index ? 14'h183 : _GEN_15398;
  wire [13:0] _GEN_15400 = 14'h3c28 == index ? 14'h180 : _GEN_15399;
  wire [13:0] _GEN_15401 = 14'h3c29 == index ? 14'h126 : _GEN_15400;
  wire [13:0] _GEN_15402 = 14'h3c2a == index ? 14'h124 : _GEN_15401;
  wire [13:0] _GEN_15403 = 14'h3c2b == index ? 14'h122 : _GEN_15402;
  wire [13:0] _GEN_15404 = 14'h3c2c == index ? 14'h120 : _GEN_15403;
  wire [13:0] _GEN_15405 = 14'h3c2d == index ? 14'h11e : _GEN_15404;
  wire [13:0] _GEN_15406 = 14'h3c2e == index ? 14'h11c : _GEN_15405;
  wire [13:0] _GEN_15407 = 14'h3c2f == index ? 14'h11a : _GEN_15406;
  wire [13:0] _GEN_15408 = 14'h3c30 == index ? 14'h118 : _GEN_15407;
  wire [13:0] _GEN_15409 = 14'h3c31 == index ? 14'h116 : _GEN_15408;
  wire [13:0] _GEN_15410 = 14'h3c32 == index ? 14'h114 : _GEN_15409;
  wire [13:0] _GEN_15411 = 14'h3c33 == index ? 14'h112 : _GEN_15410;
  wire [13:0] _GEN_15412 = 14'h3c34 == index ? 14'h110 : _GEN_15411;
  wire [13:0] _GEN_15413 = 14'h3c35 == index ? 14'h10e : _GEN_15412;
  wire [13:0] _GEN_15414 = 14'h3c36 == index ? 14'h10c : _GEN_15413;
  wire [13:0] _GEN_15415 = 14'h3c37 == index ? 14'h10a : _GEN_15414;
  wire [13:0] _GEN_15416 = 14'h3c38 == index ? 14'h108 : _GEN_15415;
  wire [13:0] _GEN_15417 = 14'h3c39 == index ? 14'h106 : _GEN_15416;
  wire [13:0] _GEN_15418 = 14'h3c3a == index ? 14'h104 : _GEN_15417;
  wire [13:0] _GEN_15419 = 14'h3c3b == index ? 14'h102 : _GEN_15418;
  wire [13:0] _GEN_15420 = 14'h3c3c == index ? 14'h100 : _GEN_15419;
  wire [13:0] _GEN_15421 = 14'h3c3d == index ? 14'hbb : _GEN_15420;
  wire [13:0] _GEN_15422 = 14'h3c3e == index ? 14'hba : _GEN_15421;
  wire [13:0] _GEN_15423 = 14'h3c3f == index ? 14'hb9 : _GEN_15422;
  wire [13:0] _GEN_15424 = 14'h3c40 == index ? 14'hb8 : _GEN_15423;
  wire [13:0] _GEN_15425 = 14'h3c41 == index ? 14'hb7 : _GEN_15424;
  wire [13:0] _GEN_15426 = 14'h3c42 == index ? 14'hb6 : _GEN_15425;
  wire [13:0] _GEN_15427 = 14'h3c43 == index ? 14'hb5 : _GEN_15426;
  wire [13:0] _GEN_15428 = 14'h3c44 == index ? 14'hb4 : _GEN_15427;
  wire [13:0] _GEN_15429 = 14'h3c45 == index ? 14'hb3 : _GEN_15428;
  wire [13:0] _GEN_15430 = 14'h3c46 == index ? 14'hb2 : _GEN_15429;
  wire [13:0] _GEN_15431 = 14'h3c47 == index ? 14'hb1 : _GEN_15430;
  wire [13:0] _GEN_15432 = 14'h3c48 == index ? 14'hb0 : _GEN_15431;
  wire [13:0] _GEN_15433 = 14'h3c49 == index ? 14'haf : _GEN_15432;
  wire [13:0] _GEN_15434 = 14'h3c4a == index ? 14'hae : _GEN_15433;
  wire [13:0] _GEN_15435 = 14'h3c4b == index ? 14'had : _GEN_15434;
  wire [13:0] _GEN_15436 = 14'h3c4c == index ? 14'hac : _GEN_15435;
  wire [13:0] _GEN_15437 = 14'h3c4d == index ? 14'hab : _GEN_15436;
  wire [13:0] _GEN_15438 = 14'h3c4e == index ? 14'haa : _GEN_15437;
  wire [13:0] _GEN_15439 = 14'h3c4f == index ? 14'ha9 : _GEN_15438;
  wire [13:0] _GEN_15440 = 14'h3c50 == index ? 14'ha8 : _GEN_15439;
  wire [13:0] _GEN_15441 = 14'h3c51 == index ? 14'ha7 : _GEN_15440;
  wire [13:0] _GEN_15442 = 14'h3c52 == index ? 14'ha6 : _GEN_15441;
  wire [13:0] _GEN_15443 = 14'h3c53 == index ? 14'ha5 : _GEN_15442;
  wire [13:0] _GEN_15444 = 14'h3c54 == index ? 14'ha4 : _GEN_15443;
  wire [13:0] _GEN_15445 = 14'h3c55 == index ? 14'ha3 : _GEN_15444;
  wire [13:0] _GEN_15446 = 14'h3c56 == index ? 14'ha2 : _GEN_15445;
  wire [13:0] _GEN_15447 = 14'h3c57 == index ? 14'ha1 : _GEN_15446;
  wire [13:0] _GEN_15448 = 14'h3c58 == index ? 14'ha0 : _GEN_15447;
  wire [13:0] _GEN_15449 = 14'h3c59 == index ? 14'h9f : _GEN_15448;
  wire [13:0] _GEN_15450 = 14'h3c5a == index ? 14'h9e : _GEN_15449;
  wire [13:0] _GEN_15451 = 14'h3c5b == index ? 14'h9d : _GEN_15450;
  wire [13:0] _GEN_15452 = 14'h3c5c == index ? 14'h9c : _GEN_15451;
  wire [13:0] _GEN_15453 = 14'h3c5d == index ? 14'h9b : _GEN_15452;
  wire [13:0] _GEN_15454 = 14'h3c5e == index ? 14'h9a : _GEN_15453;
  wire [13:0] _GEN_15455 = 14'h3c5f == index ? 14'h99 : _GEN_15454;
  wire [13:0] _GEN_15456 = 14'h3c60 == index ? 14'h98 : _GEN_15455;
  wire [13:0] _GEN_15457 = 14'h3c61 == index ? 14'h97 : _GEN_15456;
  wire [13:0] _GEN_15458 = 14'h3c62 == index ? 14'h96 : _GEN_15457;
  wire [13:0] _GEN_15459 = 14'h3c63 == index ? 14'h95 : _GEN_15458;
  wire [13:0] _GEN_15460 = 14'h3c64 == index ? 14'h94 : _GEN_15459;
  wire [13:0] _GEN_15461 = 14'h3c65 == index ? 14'h93 : _GEN_15460;
  wire [13:0] _GEN_15462 = 14'h3c66 == index ? 14'h92 : _GEN_15461;
  wire [13:0] _GEN_15463 = 14'h3c67 == index ? 14'h91 : _GEN_15462;
  wire [13:0] _GEN_15464 = 14'h3c68 == index ? 14'h90 : _GEN_15463;
  wire [13:0] _GEN_15465 = 14'h3c69 == index ? 14'h8f : _GEN_15464;
  wire [13:0] _GEN_15466 = 14'h3c6a == index ? 14'h8e : _GEN_15465;
  wire [13:0] _GEN_15467 = 14'h3c6b == index ? 14'h8d : _GEN_15466;
  wire [13:0] _GEN_15468 = 14'h3c6c == index ? 14'h8c : _GEN_15467;
  wire [13:0] _GEN_15469 = 14'h3c6d == index ? 14'h8b : _GEN_15468;
  wire [13:0] _GEN_15470 = 14'h3c6e == index ? 14'h8a : _GEN_15469;
  wire [13:0] _GEN_15471 = 14'h3c6f == index ? 14'h89 : _GEN_15470;
  wire [13:0] _GEN_15472 = 14'h3c70 == index ? 14'h88 : _GEN_15471;
  wire [13:0] _GEN_15473 = 14'h3c71 == index ? 14'h87 : _GEN_15472;
  wire [13:0] _GEN_15474 = 14'h3c72 == index ? 14'h86 : _GEN_15473;
  wire [13:0] _GEN_15475 = 14'h3c73 == index ? 14'h85 : _GEN_15474;
  wire [13:0] _GEN_15476 = 14'h3c74 == index ? 14'h84 : _GEN_15475;
  wire [13:0] _GEN_15477 = 14'h3c75 == index ? 14'h83 : _GEN_15476;
  wire [13:0] _GEN_15478 = 14'h3c76 == index ? 14'h82 : _GEN_15477;
  wire [13:0] _GEN_15479 = 14'h3c77 == index ? 14'h81 : _GEN_15478;
  wire [13:0] _GEN_15480 = 14'h3c78 == index ? 14'h80 : _GEN_15479;
  wire [13:0] _GEN_15481 = 14'h3c79 == index ? 14'h78 : _GEN_15480;
  wire [13:0] _GEN_15482 = 14'h3c7a == index ? 14'h78 : _GEN_15481;
  wire [13:0] _GEN_15483 = 14'h3c7b == index ? 14'h78 : _GEN_15482;
  wire [13:0] _GEN_15484 = 14'h3c7c == index ? 14'h78 : _GEN_15483;
  wire [13:0] _GEN_15485 = 14'h3c7d == index ? 14'h78 : _GEN_15484;
  wire [13:0] _GEN_15486 = 14'h3c7e == index ? 14'h78 : _GEN_15485;
  wire [13:0] _GEN_15487 = 14'h3c7f == index ? 14'h78 : _GEN_15486;
  wire [13:0] _GEN_15488 = 14'h3c80 == index ? 14'h0 : _GEN_15487;
  wire [13:0] _GEN_15489 = 14'h3c81 == index ? 14'h3c80 : _GEN_15488;
  wire [13:0] _GEN_15490 = 14'h3c82 == index ? 14'h1e01 : _GEN_15489;
  wire [13:0] _GEN_15491 = 14'h3c83 == index ? 14'h1401 : _GEN_15490;
  wire [13:0] _GEN_15492 = 14'h3c84 == index ? 14'hf01 : _GEN_15491;
  wire [13:0] _GEN_15493 = 14'h3c85 == index ? 14'hc01 : _GEN_15492;
  wire [13:0] _GEN_15494 = 14'h3c86 == index ? 14'ha01 : _GEN_15493;
  wire [13:0] _GEN_15495 = 14'h3c87 == index ? 14'h882 : _GEN_15494;
  wire [13:0] _GEN_15496 = 14'h3c88 == index ? 14'h781 : _GEN_15495;
  wire [13:0] _GEN_15497 = 14'h3c89 == index ? 14'h684 : _GEN_15496;
  wire [13:0] _GEN_15498 = 14'h3c8a == index ? 14'h601 : _GEN_15497;
  wire [13:0] _GEN_15499 = 14'h3c8b == index ? 14'h580 : _GEN_15498;
  wire [13:0] _GEN_15500 = 14'h3c8c == index ? 14'h501 : _GEN_15499;
  wire [13:0] _GEN_15501 = 14'h3c8d == index ? 14'h484 : _GEN_15500;
  wire [13:0] _GEN_15502 = 14'h3c8e == index ? 14'h409 : _GEN_15501;
  wire [13:0] _GEN_15503 = 14'h3c8f == index ? 14'h401 : _GEN_15502;
  wire [13:0] _GEN_15504 = 14'h3c90 == index ? 14'h389 : _GEN_15503;
  wire [13:0] _GEN_15505 = 14'h3c91 == index ? 14'h382 : _GEN_15504;
  wire [13:0] _GEN_15506 = 14'h3c92 == index ? 14'h30d : _GEN_15505;
  wire [13:0] _GEN_15507 = 14'h3c93 == index ? 14'h307 : _GEN_15506;
  wire [13:0] _GEN_15508 = 14'h3c94 == index ? 14'h301 : _GEN_15507;
  wire [13:0] _GEN_15509 = 14'h3c95 == index ? 14'h290 : _GEN_15508;
  wire [13:0] _GEN_15510 = 14'h3c96 == index ? 14'h28b : _GEN_15509;
  wire [13:0] _GEN_15511 = 14'h3c97 == index ? 14'h286 : _GEN_15510;
  wire [13:0] _GEN_15512 = 14'h3c98 == index ? 14'h281 : _GEN_15511;
  wire [13:0] _GEN_15513 = 14'h3c99 == index ? 14'h215 : _GEN_15512;
  wire [13:0] _GEN_15514 = 14'h3c9a == index ? 14'h211 : _GEN_15513;
  wire [13:0] _GEN_15515 = 14'h3c9b == index ? 14'h20d : _GEN_15514;
  wire [13:0] _GEN_15516 = 14'h3c9c == index ? 14'h209 : _GEN_15515;
  wire [13:0] _GEN_15517 = 14'h3c9d == index ? 14'h205 : _GEN_15516;
  wire [13:0] _GEN_15518 = 14'h3c9e == index ? 14'h201 : _GEN_15517;
  wire [13:0] _GEN_15519 = 14'h3c9f == index ? 14'h19c : _GEN_15518;
  wire [13:0] _GEN_15520 = 14'h3ca0 == index ? 14'h199 : _GEN_15519;
  wire [13:0] _GEN_15521 = 14'h3ca1 == index ? 14'h196 : _GEN_15520;
  wire [13:0] _GEN_15522 = 14'h3ca2 == index ? 14'h193 : _GEN_15521;
  wire [13:0] _GEN_15523 = 14'h3ca3 == index ? 14'h190 : _GEN_15522;
  wire [13:0] _GEN_15524 = 14'h3ca4 == index ? 14'h18d : _GEN_15523;
  wire [13:0] _GEN_15525 = 14'h3ca5 == index ? 14'h18a : _GEN_15524;
  wire [13:0] _GEN_15526 = 14'h3ca6 == index ? 14'h187 : _GEN_15525;
  wire [13:0] _GEN_15527 = 14'h3ca7 == index ? 14'h184 : _GEN_15526;
  wire [13:0] _GEN_15528 = 14'h3ca8 == index ? 14'h181 : _GEN_15527;
  wire [13:0] _GEN_15529 = 14'h3ca9 == index ? 14'h127 : _GEN_15528;
  wire [13:0] _GEN_15530 = 14'h3caa == index ? 14'h125 : _GEN_15529;
  wire [13:0] _GEN_15531 = 14'h3cab == index ? 14'h123 : _GEN_15530;
  wire [13:0] _GEN_15532 = 14'h3cac == index ? 14'h121 : _GEN_15531;
  wire [13:0] _GEN_15533 = 14'h3cad == index ? 14'h11f : _GEN_15532;
  wire [13:0] _GEN_15534 = 14'h3cae == index ? 14'h11d : _GEN_15533;
  wire [13:0] _GEN_15535 = 14'h3caf == index ? 14'h11b : _GEN_15534;
  wire [13:0] _GEN_15536 = 14'h3cb0 == index ? 14'h119 : _GEN_15535;
  wire [13:0] _GEN_15537 = 14'h3cb1 == index ? 14'h117 : _GEN_15536;
  wire [13:0] _GEN_15538 = 14'h3cb2 == index ? 14'h115 : _GEN_15537;
  wire [13:0] _GEN_15539 = 14'h3cb3 == index ? 14'h113 : _GEN_15538;
  wire [13:0] _GEN_15540 = 14'h3cb4 == index ? 14'h111 : _GEN_15539;
  wire [13:0] _GEN_15541 = 14'h3cb5 == index ? 14'h10f : _GEN_15540;
  wire [13:0] _GEN_15542 = 14'h3cb6 == index ? 14'h10d : _GEN_15541;
  wire [13:0] _GEN_15543 = 14'h3cb7 == index ? 14'h10b : _GEN_15542;
  wire [13:0] _GEN_15544 = 14'h3cb8 == index ? 14'h109 : _GEN_15543;
  wire [13:0] _GEN_15545 = 14'h3cb9 == index ? 14'h107 : _GEN_15544;
  wire [13:0] _GEN_15546 = 14'h3cba == index ? 14'h105 : _GEN_15545;
  wire [13:0] _GEN_15547 = 14'h3cbb == index ? 14'h103 : _GEN_15546;
  wire [13:0] _GEN_15548 = 14'h3cbc == index ? 14'h101 : _GEN_15547;
  wire [13:0] _GEN_15549 = 14'h3cbd == index ? 14'hbc : _GEN_15548;
  wire [13:0] _GEN_15550 = 14'h3cbe == index ? 14'hbb : _GEN_15549;
  wire [13:0] _GEN_15551 = 14'h3cbf == index ? 14'hba : _GEN_15550;
  wire [13:0] _GEN_15552 = 14'h3cc0 == index ? 14'hb9 : _GEN_15551;
  wire [13:0] _GEN_15553 = 14'h3cc1 == index ? 14'hb8 : _GEN_15552;
  wire [13:0] _GEN_15554 = 14'h3cc2 == index ? 14'hb7 : _GEN_15553;
  wire [13:0] _GEN_15555 = 14'h3cc3 == index ? 14'hb6 : _GEN_15554;
  wire [13:0] _GEN_15556 = 14'h3cc4 == index ? 14'hb5 : _GEN_15555;
  wire [13:0] _GEN_15557 = 14'h3cc5 == index ? 14'hb4 : _GEN_15556;
  wire [13:0] _GEN_15558 = 14'h3cc6 == index ? 14'hb3 : _GEN_15557;
  wire [13:0] _GEN_15559 = 14'h3cc7 == index ? 14'hb2 : _GEN_15558;
  wire [13:0] _GEN_15560 = 14'h3cc8 == index ? 14'hb1 : _GEN_15559;
  wire [13:0] _GEN_15561 = 14'h3cc9 == index ? 14'hb0 : _GEN_15560;
  wire [13:0] _GEN_15562 = 14'h3cca == index ? 14'haf : _GEN_15561;
  wire [13:0] _GEN_15563 = 14'h3ccb == index ? 14'hae : _GEN_15562;
  wire [13:0] _GEN_15564 = 14'h3ccc == index ? 14'had : _GEN_15563;
  wire [13:0] _GEN_15565 = 14'h3ccd == index ? 14'hac : _GEN_15564;
  wire [13:0] _GEN_15566 = 14'h3cce == index ? 14'hab : _GEN_15565;
  wire [13:0] _GEN_15567 = 14'h3ccf == index ? 14'haa : _GEN_15566;
  wire [13:0] _GEN_15568 = 14'h3cd0 == index ? 14'ha9 : _GEN_15567;
  wire [13:0] _GEN_15569 = 14'h3cd1 == index ? 14'ha8 : _GEN_15568;
  wire [13:0] _GEN_15570 = 14'h3cd2 == index ? 14'ha7 : _GEN_15569;
  wire [13:0] _GEN_15571 = 14'h3cd3 == index ? 14'ha6 : _GEN_15570;
  wire [13:0] _GEN_15572 = 14'h3cd4 == index ? 14'ha5 : _GEN_15571;
  wire [13:0] _GEN_15573 = 14'h3cd5 == index ? 14'ha4 : _GEN_15572;
  wire [13:0] _GEN_15574 = 14'h3cd6 == index ? 14'ha3 : _GEN_15573;
  wire [13:0] _GEN_15575 = 14'h3cd7 == index ? 14'ha2 : _GEN_15574;
  wire [13:0] _GEN_15576 = 14'h3cd8 == index ? 14'ha1 : _GEN_15575;
  wire [13:0] _GEN_15577 = 14'h3cd9 == index ? 14'ha0 : _GEN_15576;
  wire [13:0] _GEN_15578 = 14'h3cda == index ? 14'h9f : _GEN_15577;
  wire [13:0] _GEN_15579 = 14'h3cdb == index ? 14'h9e : _GEN_15578;
  wire [13:0] _GEN_15580 = 14'h3cdc == index ? 14'h9d : _GEN_15579;
  wire [13:0] _GEN_15581 = 14'h3cdd == index ? 14'h9c : _GEN_15580;
  wire [13:0] _GEN_15582 = 14'h3cde == index ? 14'h9b : _GEN_15581;
  wire [13:0] _GEN_15583 = 14'h3cdf == index ? 14'h9a : _GEN_15582;
  wire [13:0] _GEN_15584 = 14'h3ce0 == index ? 14'h99 : _GEN_15583;
  wire [13:0] _GEN_15585 = 14'h3ce1 == index ? 14'h98 : _GEN_15584;
  wire [13:0] _GEN_15586 = 14'h3ce2 == index ? 14'h97 : _GEN_15585;
  wire [13:0] _GEN_15587 = 14'h3ce3 == index ? 14'h96 : _GEN_15586;
  wire [13:0] _GEN_15588 = 14'h3ce4 == index ? 14'h95 : _GEN_15587;
  wire [13:0] _GEN_15589 = 14'h3ce5 == index ? 14'h94 : _GEN_15588;
  wire [13:0] _GEN_15590 = 14'h3ce6 == index ? 14'h93 : _GEN_15589;
  wire [13:0] _GEN_15591 = 14'h3ce7 == index ? 14'h92 : _GEN_15590;
  wire [13:0] _GEN_15592 = 14'h3ce8 == index ? 14'h91 : _GEN_15591;
  wire [13:0] _GEN_15593 = 14'h3ce9 == index ? 14'h90 : _GEN_15592;
  wire [13:0] _GEN_15594 = 14'h3cea == index ? 14'h8f : _GEN_15593;
  wire [13:0] _GEN_15595 = 14'h3ceb == index ? 14'h8e : _GEN_15594;
  wire [13:0] _GEN_15596 = 14'h3cec == index ? 14'h8d : _GEN_15595;
  wire [13:0] _GEN_15597 = 14'h3ced == index ? 14'h8c : _GEN_15596;
  wire [13:0] _GEN_15598 = 14'h3cee == index ? 14'h8b : _GEN_15597;
  wire [13:0] _GEN_15599 = 14'h3cef == index ? 14'h8a : _GEN_15598;
  wire [13:0] _GEN_15600 = 14'h3cf0 == index ? 14'h89 : _GEN_15599;
  wire [13:0] _GEN_15601 = 14'h3cf1 == index ? 14'h88 : _GEN_15600;
  wire [13:0] _GEN_15602 = 14'h3cf2 == index ? 14'h87 : _GEN_15601;
  wire [13:0] _GEN_15603 = 14'h3cf3 == index ? 14'h86 : _GEN_15602;
  wire [13:0] _GEN_15604 = 14'h3cf4 == index ? 14'h85 : _GEN_15603;
  wire [13:0] _GEN_15605 = 14'h3cf5 == index ? 14'h84 : _GEN_15604;
  wire [13:0] _GEN_15606 = 14'h3cf6 == index ? 14'h83 : _GEN_15605;
  wire [13:0] _GEN_15607 = 14'h3cf7 == index ? 14'h82 : _GEN_15606;
  wire [13:0] _GEN_15608 = 14'h3cf8 == index ? 14'h81 : _GEN_15607;
  wire [13:0] _GEN_15609 = 14'h3cf9 == index ? 14'h80 : _GEN_15608;
  wire [13:0] _GEN_15610 = 14'h3cfa == index ? 14'h79 : _GEN_15609;
  wire [13:0] _GEN_15611 = 14'h3cfb == index ? 14'h79 : _GEN_15610;
  wire [13:0] _GEN_15612 = 14'h3cfc == index ? 14'h79 : _GEN_15611;
  wire [13:0] _GEN_15613 = 14'h3cfd == index ? 14'h79 : _GEN_15612;
  wire [13:0] _GEN_15614 = 14'h3cfe == index ? 14'h79 : _GEN_15613;
  wire [13:0] _GEN_15615 = 14'h3cff == index ? 14'h79 : _GEN_15614;
  wire [13:0] _GEN_15616 = 14'h3d00 == index ? 14'h0 : _GEN_15615;
  wire [13:0] _GEN_15617 = 14'h3d01 == index ? 14'h3d00 : _GEN_15616;
  wire [13:0] _GEN_15618 = 14'h3d02 == index ? 14'h1e80 : _GEN_15617;
  wire [13:0] _GEN_15619 = 14'h3d03 == index ? 14'h1402 : _GEN_15618;
  wire [13:0] _GEN_15620 = 14'h3d04 == index ? 14'hf02 : _GEN_15619;
  wire [13:0] _GEN_15621 = 14'h3d05 == index ? 14'hc02 : _GEN_15620;
  wire [13:0] _GEN_15622 = 14'h3d06 == index ? 14'ha02 : _GEN_15621;
  wire [13:0] _GEN_15623 = 14'h3d07 == index ? 14'h883 : _GEN_15622;
  wire [13:0] _GEN_15624 = 14'h3d08 == index ? 14'h782 : _GEN_15623;
  wire [13:0] _GEN_15625 = 14'h3d09 == index ? 14'h685 : _GEN_15624;
  wire [13:0] _GEN_15626 = 14'h3d0a == index ? 14'h602 : _GEN_15625;
  wire [13:0] _GEN_15627 = 14'h3d0b == index ? 14'h581 : _GEN_15626;
  wire [13:0] _GEN_15628 = 14'h3d0c == index ? 14'h502 : _GEN_15627;
  wire [13:0] _GEN_15629 = 14'h3d0d == index ? 14'h485 : _GEN_15628;
  wire [13:0] _GEN_15630 = 14'h3d0e == index ? 14'h40a : _GEN_15629;
  wire [13:0] _GEN_15631 = 14'h3d0f == index ? 14'h402 : _GEN_15630;
  wire [13:0] _GEN_15632 = 14'h3d10 == index ? 14'h38a : _GEN_15631;
  wire [13:0] _GEN_15633 = 14'h3d11 == index ? 14'h383 : _GEN_15632;
  wire [13:0] _GEN_15634 = 14'h3d12 == index ? 14'h30e : _GEN_15633;
  wire [13:0] _GEN_15635 = 14'h3d13 == index ? 14'h308 : _GEN_15634;
  wire [13:0] _GEN_15636 = 14'h3d14 == index ? 14'h302 : _GEN_15635;
  wire [13:0] _GEN_15637 = 14'h3d15 == index ? 14'h291 : _GEN_15636;
  wire [13:0] _GEN_15638 = 14'h3d16 == index ? 14'h28c : _GEN_15637;
  wire [13:0] _GEN_15639 = 14'h3d17 == index ? 14'h287 : _GEN_15638;
  wire [13:0] _GEN_15640 = 14'h3d18 == index ? 14'h282 : _GEN_15639;
  wire [13:0] _GEN_15641 = 14'h3d19 == index ? 14'h216 : _GEN_15640;
  wire [13:0] _GEN_15642 = 14'h3d1a == index ? 14'h212 : _GEN_15641;
  wire [13:0] _GEN_15643 = 14'h3d1b == index ? 14'h20e : _GEN_15642;
  wire [13:0] _GEN_15644 = 14'h3d1c == index ? 14'h20a : _GEN_15643;
  wire [13:0] _GEN_15645 = 14'h3d1d == index ? 14'h206 : _GEN_15644;
  wire [13:0] _GEN_15646 = 14'h3d1e == index ? 14'h202 : _GEN_15645;
  wire [13:0] _GEN_15647 = 14'h3d1f == index ? 14'h19d : _GEN_15646;
  wire [13:0] _GEN_15648 = 14'h3d20 == index ? 14'h19a : _GEN_15647;
  wire [13:0] _GEN_15649 = 14'h3d21 == index ? 14'h197 : _GEN_15648;
  wire [13:0] _GEN_15650 = 14'h3d22 == index ? 14'h194 : _GEN_15649;
  wire [13:0] _GEN_15651 = 14'h3d23 == index ? 14'h191 : _GEN_15650;
  wire [13:0] _GEN_15652 = 14'h3d24 == index ? 14'h18e : _GEN_15651;
  wire [13:0] _GEN_15653 = 14'h3d25 == index ? 14'h18b : _GEN_15652;
  wire [13:0] _GEN_15654 = 14'h3d26 == index ? 14'h188 : _GEN_15653;
  wire [13:0] _GEN_15655 = 14'h3d27 == index ? 14'h185 : _GEN_15654;
  wire [13:0] _GEN_15656 = 14'h3d28 == index ? 14'h182 : _GEN_15655;
  wire [13:0] _GEN_15657 = 14'h3d29 == index ? 14'h128 : _GEN_15656;
  wire [13:0] _GEN_15658 = 14'h3d2a == index ? 14'h126 : _GEN_15657;
  wire [13:0] _GEN_15659 = 14'h3d2b == index ? 14'h124 : _GEN_15658;
  wire [13:0] _GEN_15660 = 14'h3d2c == index ? 14'h122 : _GEN_15659;
  wire [13:0] _GEN_15661 = 14'h3d2d == index ? 14'h120 : _GEN_15660;
  wire [13:0] _GEN_15662 = 14'h3d2e == index ? 14'h11e : _GEN_15661;
  wire [13:0] _GEN_15663 = 14'h3d2f == index ? 14'h11c : _GEN_15662;
  wire [13:0] _GEN_15664 = 14'h3d30 == index ? 14'h11a : _GEN_15663;
  wire [13:0] _GEN_15665 = 14'h3d31 == index ? 14'h118 : _GEN_15664;
  wire [13:0] _GEN_15666 = 14'h3d32 == index ? 14'h116 : _GEN_15665;
  wire [13:0] _GEN_15667 = 14'h3d33 == index ? 14'h114 : _GEN_15666;
  wire [13:0] _GEN_15668 = 14'h3d34 == index ? 14'h112 : _GEN_15667;
  wire [13:0] _GEN_15669 = 14'h3d35 == index ? 14'h110 : _GEN_15668;
  wire [13:0] _GEN_15670 = 14'h3d36 == index ? 14'h10e : _GEN_15669;
  wire [13:0] _GEN_15671 = 14'h3d37 == index ? 14'h10c : _GEN_15670;
  wire [13:0] _GEN_15672 = 14'h3d38 == index ? 14'h10a : _GEN_15671;
  wire [13:0] _GEN_15673 = 14'h3d39 == index ? 14'h108 : _GEN_15672;
  wire [13:0] _GEN_15674 = 14'h3d3a == index ? 14'h106 : _GEN_15673;
  wire [13:0] _GEN_15675 = 14'h3d3b == index ? 14'h104 : _GEN_15674;
  wire [13:0] _GEN_15676 = 14'h3d3c == index ? 14'h102 : _GEN_15675;
  wire [13:0] _GEN_15677 = 14'h3d3d == index ? 14'h100 : _GEN_15676;
  wire [13:0] _GEN_15678 = 14'h3d3e == index ? 14'hbc : _GEN_15677;
  wire [13:0] _GEN_15679 = 14'h3d3f == index ? 14'hbb : _GEN_15678;
  wire [13:0] _GEN_15680 = 14'h3d40 == index ? 14'hba : _GEN_15679;
  wire [13:0] _GEN_15681 = 14'h3d41 == index ? 14'hb9 : _GEN_15680;
  wire [13:0] _GEN_15682 = 14'h3d42 == index ? 14'hb8 : _GEN_15681;
  wire [13:0] _GEN_15683 = 14'h3d43 == index ? 14'hb7 : _GEN_15682;
  wire [13:0] _GEN_15684 = 14'h3d44 == index ? 14'hb6 : _GEN_15683;
  wire [13:0] _GEN_15685 = 14'h3d45 == index ? 14'hb5 : _GEN_15684;
  wire [13:0] _GEN_15686 = 14'h3d46 == index ? 14'hb4 : _GEN_15685;
  wire [13:0] _GEN_15687 = 14'h3d47 == index ? 14'hb3 : _GEN_15686;
  wire [13:0] _GEN_15688 = 14'h3d48 == index ? 14'hb2 : _GEN_15687;
  wire [13:0] _GEN_15689 = 14'h3d49 == index ? 14'hb1 : _GEN_15688;
  wire [13:0] _GEN_15690 = 14'h3d4a == index ? 14'hb0 : _GEN_15689;
  wire [13:0] _GEN_15691 = 14'h3d4b == index ? 14'haf : _GEN_15690;
  wire [13:0] _GEN_15692 = 14'h3d4c == index ? 14'hae : _GEN_15691;
  wire [13:0] _GEN_15693 = 14'h3d4d == index ? 14'had : _GEN_15692;
  wire [13:0] _GEN_15694 = 14'h3d4e == index ? 14'hac : _GEN_15693;
  wire [13:0] _GEN_15695 = 14'h3d4f == index ? 14'hab : _GEN_15694;
  wire [13:0] _GEN_15696 = 14'h3d50 == index ? 14'haa : _GEN_15695;
  wire [13:0] _GEN_15697 = 14'h3d51 == index ? 14'ha9 : _GEN_15696;
  wire [13:0] _GEN_15698 = 14'h3d52 == index ? 14'ha8 : _GEN_15697;
  wire [13:0] _GEN_15699 = 14'h3d53 == index ? 14'ha7 : _GEN_15698;
  wire [13:0] _GEN_15700 = 14'h3d54 == index ? 14'ha6 : _GEN_15699;
  wire [13:0] _GEN_15701 = 14'h3d55 == index ? 14'ha5 : _GEN_15700;
  wire [13:0] _GEN_15702 = 14'h3d56 == index ? 14'ha4 : _GEN_15701;
  wire [13:0] _GEN_15703 = 14'h3d57 == index ? 14'ha3 : _GEN_15702;
  wire [13:0] _GEN_15704 = 14'h3d58 == index ? 14'ha2 : _GEN_15703;
  wire [13:0] _GEN_15705 = 14'h3d59 == index ? 14'ha1 : _GEN_15704;
  wire [13:0] _GEN_15706 = 14'h3d5a == index ? 14'ha0 : _GEN_15705;
  wire [13:0] _GEN_15707 = 14'h3d5b == index ? 14'h9f : _GEN_15706;
  wire [13:0] _GEN_15708 = 14'h3d5c == index ? 14'h9e : _GEN_15707;
  wire [13:0] _GEN_15709 = 14'h3d5d == index ? 14'h9d : _GEN_15708;
  wire [13:0] _GEN_15710 = 14'h3d5e == index ? 14'h9c : _GEN_15709;
  wire [13:0] _GEN_15711 = 14'h3d5f == index ? 14'h9b : _GEN_15710;
  wire [13:0] _GEN_15712 = 14'h3d60 == index ? 14'h9a : _GEN_15711;
  wire [13:0] _GEN_15713 = 14'h3d61 == index ? 14'h99 : _GEN_15712;
  wire [13:0] _GEN_15714 = 14'h3d62 == index ? 14'h98 : _GEN_15713;
  wire [13:0] _GEN_15715 = 14'h3d63 == index ? 14'h97 : _GEN_15714;
  wire [13:0] _GEN_15716 = 14'h3d64 == index ? 14'h96 : _GEN_15715;
  wire [13:0] _GEN_15717 = 14'h3d65 == index ? 14'h95 : _GEN_15716;
  wire [13:0] _GEN_15718 = 14'h3d66 == index ? 14'h94 : _GEN_15717;
  wire [13:0] _GEN_15719 = 14'h3d67 == index ? 14'h93 : _GEN_15718;
  wire [13:0] _GEN_15720 = 14'h3d68 == index ? 14'h92 : _GEN_15719;
  wire [13:0] _GEN_15721 = 14'h3d69 == index ? 14'h91 : _GEN_15720;
  wire [13:0] _GEN_15722 = 14'h3d6a == index ? 14'h90 : _GEN_15721;
  wire [13:0] _GEN_15723 = 14'h3d6b == index ? 14'h8f : _GEN_15722;
  wire [13:0] _GEN_15724 = 14'h3d6c == index ? 14'h8e : _GEN_15723;
  wire [13:0] _GEN_15725 = 14'h3d6d == index ? 14'h8d : _GEN_15724;
  wire [13:0] _GEN_15726 = 14'h3d6e == index ? 14'h8c : _GEN_15725;
  wire [13:0] _GEN_15727 = 14'h3d6f == index ? 14'h8b : _GEN_15726;
  wire [13:0] _GEN_15728 = 14'h3d70 == index ? 14'h8a : _GEN_15727;
  wire [13:0] _GEN_15729 = 14'h3d71 == index ? 14'h89 : _GEN_15728;
  wire [13:0] _GEN_15730 = 14'h3d72 == index ? 14'h88 : _GEN_15729;
  wire [13:0] _GEN_15731 = 14'h3d73 == index ? 14'h87 : _GEN_15730;
  wire [13:0] _GEN_15732 = 14'h3d74 == index ? 14'h86 : _GEN_15731;
  wire [13:0] _GEN_15733 = 14'h3d75 == index ? 14'h85 : _GEN_15732;
  wire [13:0] _GEN_15734 = 14'h3d76 == index ? 14'h84 : _GEN_15733;
  wire [13:0] _GEN_15735 = 14'h3d77 == index ? 14'h83 : _GEN_15734;
  wire [13:0] _GEN_15736 = 14'h3d78 == index ? 14'h82 : _GEN_15735;
  wire [13:0] _GEN_15737 = 14'h3d79 == index ? 14'h81 : _GEN_15736;
  wire [13:0] _GEN_15738 = 14'h3d7a == index ? 14'h80 : _GEN_15737;
  wire [13:0] _GEN_15739 = 14'h3d7b == index ? 14'h7a : _GEN_15738;
  wire [13:0] _GEN_15740 = 14'h3d7c == index ? 14'h7a : _GEN_15739;
  wire [13:0] _GEN_15741 = 14'h3d7d == index ? 14'h7a : _GEN_15740;
  wire [13:0] _GEN_15742 = 14'h3d7e == index ? 14'h7a : _GEN_15741;
  wire [13:0] _GEN_15743 = 14'h3d7f == index ? 14'h7a : _GEN_15742;
  wire [13:0] _GEN_15744 = 14'h3d80 == index ? 14'h0 : _GEN_15743;
  wire [13:0] _GEN_15745 = 14'h3d81 == index ? 14'h3d80 : _GEN_15744;
  wire [13:0] _GEN_15746 = 14'h3d82 == index ? 14'h1e81 : _GEN_15745;
  wire [13:0] _GEN_15747 = 14'h3d83 == index ? 14'h1480 : _GEN_15746;
  wire [13:0] _GEN_15748 = 14'h3d84 == index ? 14'hf03 : _GEN_15747;
  wire [13:0] _GEN_15749 = 14'h3d85 == index ? 14'hc03 : _GEN_15748;
  wire [13:0] _GEN_15750 = 14'h3d86 == index ? 14'ha03 : _GEN_15749;
  wire [13:0] _GEN_15751 = 14'h3d87 == index ? 14'h884 : _GEN_15750;
  wire [13:0] _GEN_15752 = 14'h3d88 == index ? 14'h783 : _GEN_15751;
  wire [13:0] _GEN_15753 = 14'h3d89 == index ? 14'h686 : _GEN_15752;
  wire [13:0] _GEN_15754 = 14'h3d8a == index ? 14'h603 : _GEN_15753;
  wire [13:0] _GEN_15755 = 14'h3d8b == index ? 14'h582 : _GEN_15754;
  wire [13:0] _GEN_15756 = 14'h3d8c == index ? 14'h503 : _GEN_15755;
  wire [13:0] _GEN_15757 = 14'h3d8d == index ? 14'h486 : _GEN_15756;
  wire [13:0] _GEN_15758 = 14'h3d8e == index ? 14'h40b : _GEN_15757;
  wire [13:0] _GEN_15759 = 14'h3d8f == index ? 14'h403 : _GEN_15758;
  wire [13:0] _GEN_15760 = 14'h3d90 == index ? 14'h38b : _GEN_15759;
  wire [13:0] _GEN_15761 = 14'h3d91 == index ? 14'h384 : _GEN_15760;
  wire [13:0] _GEN_15762 = 14'h3d92 == index ? 14'h30f : _GEN_15761;
  wire [13:0] _GEN_15763 = 14'h3d93 == index ? 14'h309 : _GEN_15762;
  wire [13:0] _GEN_15764 = 14'h3d94 == index ? 14'h303 : _GEN_15763;
  wire [13:0] _GEN_15765 = 14'h3d95 == index ? 14'h292 : _GEN_15764;
  wire [13:0] _GEN_15766 = 14'h3d96 == index ? 14'h28d : _GEN_15765;
  wire [13:0] _GEN_15767 = 14'h3d97 == index ? 14'h288 : _GEN_15766;
  wire [13:0] _GEN_15768 = 14'h3d98 == index ? 14'h283 : _GEN_15767;
  wire [13:0] _GEN_15769 = 14'h3d99 == index ? 14'h217 : _GEN_15768;
  wire [13:0] _GEN_15770 = 14'h3d9a == index ? 14'h213 : _GEN_15769;
  wire [13:0] _GEN_15771 = 14'h3d9b == index ? 14'h20f : _GEN_15770;
  wire [13:0] _GEN_15772 = 14'h3d9c == index ? 14'h20b : _GEN_15771;
  wire [13:0] _GEN_15773 = 14'h3d9d == index ? 14'h207 : _GEN_15772;
  wire [13:0] _GEN_15774 = 14'h3d9e == index ? 14'h203 : _GEN_15773;
  wire [13:0] _GEN_15775 = 14'h3d9f == index ? 14'h19e : _GEN_15774;
  wire [13:0] _GEN_15776 = 14'h3da0 == index ? 14'h19b : _GEN_15775;
  wire [13:0] _GEN_15777 = 14'h3da1 == index ? 14'h198 : _GEN_15776;
  wire [13:0] _GEN_15778 = 14'h3da2 == index ? 14'h195 : _GEN_15777;
  wire [13:0] _GEN_15779 = 14'h3da3 == index ? 14'h192 : _GEN_15778;
  wire [13:0] _GEN_15780 = 14'h3da4 == index ? 14'h18f : _GEN_15779;
  wire [13:0] _GEN_15781 = 14'h3da5 == index ? 14'h18c : _GEN_15780;
  wire [13:0] _GEN_15782 = 14'h3da6 == index ? 14'h189 : _GEN_15781;
  wire [13:0] _GEN_15783 = 14'h3da7 == index ? 14'h186 : _GEN_15782;
  wire [13:0] _GEN_15784 = 14'h3da8 == index ? 14'h183 : _GEN_15783;
  wire [13:0] _GEN_15785 = 14'h3da9 == index ? 14'h180 : _GEN_15784;
  wire [13:0] _GEN_15786 = 14'h3daa == index ? 14'h127 : _GEN_15785;
  wire [13:0] _GEN_15787 = 14'h3dab == index ? 14'h125 : _GEN_15786;
  wire [13:0] _GEN_15788 = 14'h3dac == index ? 14'h123 : _GEN_15787;
  wire [13:0] _GEN_15789 = 14'h3dad == index ? 14'h121 : _GEN_15788;
  wire [13:0] _GEN_15790 = 14'h3dae == index ? 14'h11f : _GEN_15789;
  wire [13:0] _GEN_15791 = 14'h3daf == index ? 14'h11d : _GEN_15790;
  wire [13:0] _GEN_15792 = 14'h3db0 == index ? 14'h11b : _GEN_15791;
  wire [13:0] _GEN_15793 = 14'h3db1 == index ? 14'h119 : _GEN_15792;
  wire [13:0] _GEN_15794 = 14'h3db2 == index ? 14'h117 : _GEN_15793;
  wire [13:0] _GEN_15795 = 14'h3db3 == index ? 14'h115 : _GEN_15794;
  wire [13:0] _GEN_15796 = 14'h3db4 == index ? 14'h113 : _GEN_15795;
  wire [13:0] _GEN_15797 = 14'h3db5 == index ? 14'h111 : _GEN_15796;
  wire [13:0] _GEN_15798 = 14'h3db6 == index ? 14'h10f : _GEN_15797;
  wire [13:0] _GEN_15799 = 14'h3db7 == index ? 14'h10d : _GEN_15798;
  wire [13:0] _GEN_15800 = 14'h3db8 == index ? 14'h10b : _GEN_15799;
  wire [13:0] _GEN_15801 = 14'h3db9 == index ? 14'h109 : _GEN_15800;
  wire [13:0] _GEN_15802 = 14'h3dba == index ? 14'h107 : _GEN_15801;
  wire [13:0] _GEN_15803 = 14'h3dbb == index ? 14'h105 : _GEN_15802;
  wire [13:0] _GEN_15804 = 14'h3dbc == index ? 14'h103 : _GEN_15803;
  wire [13:0] _GEN_15805 = 14'h3dbd == index ? 14'h101 : _GEN_15804;
  wire [13:0] _GEN_15806 = 14'h3dbe == index ? 14'hbd : _GEN_15805;
  wire [13:0] _GEN_15807 = 14'h3dbf == index ? 14'hbc : _GEN_15806;
  wire [13:0] _GEN_15808 = 14'h3dc0 == index ? 14'hbb : _GEN_15807;
  wire [13:0] _GEN_15809 = 14'h3dc1 == index ? 14'hba : _GEN_15808;
  wire [13:0] _GEN_15810 = 14'h3dc2 == index ? 14'hb9 : _GEN_15809;
  wire [13:0] _GEN_15811 = 14'h3dc3 == index ? 14'hb8 : _GEN_15810;
  wire [13:0] _GEN_15812 = 14'h3dc4 == index ? 14'hb7 : _GEN_15811;
  wire [13:0] _GEN_15813 = 14'h3dc5 == index ? 14'hb6 : _GEN_15812;
  wire [13:0] _GEN_15814 = 14'h3dc6 == index ? 14'hb5 : _GEN_15813;
  wire [13:0] _GEN_15815 = 14'h3dc7 == index ? 14'hb4 : _GEN_15814;
  wire [13:0] _GEN_15816 = 14'h3dc8 == index ? 14'hb3 : _GEN_15815;
  wire [13:0] _GEN_15817 = 14'h3dc9 == index ? 14'hb2 : _GEN_15816;
  wire [13:0] _GEN_15818 = 14'h3dca == index ? 14'hb1 : _GEN_15817;
  wire [13:0] _GEN_15819 = 14'h3dcb == index ? 14'hb0 : _GEN_15818;
  wire [13:0] _GEN_15820 = 14'h3dcc == index ? 14'haf : _GEN_15819;
  wire [13:0] _GEN_15821 = 14'h3dcd == index ? 14'hae : _GEN_15820;
  wire [13:0] _GEN_15822 = 14'h3dce == index ? 14'had : _GEN_15821;
  wire [13:0] _GEN_15823 = 14'h3dcf == index ? 14'hac : _GEN_15822;
  wire [13:0] _GEN_15824 = 14'h3dd0 == index ? 14'hab : _GEN_15823;
  wire [13:0] _GEN_15825 = 14'h3dd1 == index ? 14'haa : _GEN_15824;
  wire [13:0] _GEN_15826 = 14'h3dd2 == index ? 14'ha9 : _GEN_15825;
  wire [13:0] _GEN_15827 = 14'h3dd3 == index ? 14'ha8 : _GEN_15826;
  wire [13:0] _GEN_15828 = 14'h3dd4 == index ? 14'ha7 : _GEN_15827;
  wire [13:0] _GEN_15829 = 14'h3dd5 == index ? 14'ha6 : _GEN_15828;
  wire [13:0] _GEN_15830 = 14'h3dd6 == index ? 14'ha5 : _GEN_15829;
  wire [13:0] _GEN_15831 = 14'h3dd7 == index ? 14'ha4 : _GEN_15830;
  wire [13:0] _GEN_15832 = 14'h3dd8 == index ? 14'ha3 : _GEN_15831;
  wire [13:0] _GEN_15833 = 14'h3dd9 == index ? 14'ha2 : _GEN_15832;
  wire [13:0] _GEN_15834 = 14'h3dda == index ? 14'ha1 : _GEN_15833;
  wire [13:0] _GEN_15835 = 14'h3ddb == index ? 14'ha0 : _GEN_15834;
  wire [13:0] _GEN_15836 = 14'h3ddc == index ? 14'h9f : _GEN_15835;
  wire [13:0] _GEN_15837 = 14'h3ddd == index ? 14'h9e : _GEN_15836;
  wire [13:0] _GEN_15838 = 14'h3dde == index ? 14'h9d : _GEN_15837;
  wire [13:0] _GEN_15839 = 14'h3ddf == index ? 14'h9c : _GEN_15838;
  wire [13:0] _GEN_15840 = 14'h3de0 == index ? 14'h9b : _GEN_15839;
  wire [13:0] _GEN_15841 = 14'h3de1 == index ? 14'h9a : _GEN_15840;
  wire [13:0] _GEN_15842 = 14'h3de2 == index ? 14'h99 : _GEN_15841;
  wire [13:0] _GEN_15843 = 14'h3de3 == index ? 14'h98 : _GEN_15842;
  wire [13:0] _GEN_15844 = 14'h3de4 == index ? 14'h97 : _GEN_15843;
  wire [13:0] _GEN_15845 = 14'h3de5 == index ? 14'h96 : _GEN_15844;
  wire [13:0] _GEN_15846 = 14'h3de6 == index ? 14'h95 : _GEN_15845;
  wire [13:0] _GEN_15847 = 14'h3de7 == index ? 14'h94 : _GEN_15846;
  wire [13:0] _GEN_15848 = 14'h3de8 == index ? 14'h93 : _GEN_15847;
  wire [13:0] _GEN_15849 = 14'h3de9 == index ? 14'h92 : _GEN_15848;
  wire [13:0] _GEN_15850 = 14'h3dea == index ? 14'h91 : _GEN_15849;
  wire [13:0] _GEN_15851 = 14'h3deb == index ? 14'h90 : _GEN_15850;
  wire [13:0] _GEN_15852 = 14'h3dec == index ? 14'h8f : _GEN_15851;
  wire [13:0] _GEN_15853 = 14'h3ded == index ? 14'h8e : _GEN_15852;
  wire [13:0] _GEN_15854 = 14'h3dee == index ? 14'h8d : _GEN_15853;
  wire [13:0] _GEN_15855 = 14'h3def == index ? 14'h8c : _GEN_15854;
  wire [13:0] _GEN_15856 = 14'h3df0 == index ? 14'h8b : _GEN_15855;
  wire [13:0] _GEN_15857 = 14'h3df1 == index ? 14'h8a : _GEN_15856;
  wire [13:0] _GEN_15858 = 14'h3df2 == index ? 14'h89 : _GEN_15857;
  wire [13:0] _GEN_15859 = 14'h3df3 == index ? 14'h88 : _GEN_15858;
  wire [13:0] _GEN_15860 = 14'h3df4 == index ? 14'h87 : _GEN_15859;
  wire [13:0] _GEN_15861 = 14'h3df5 == index ? 14'h86 : _GEN_15860;
  wire [13:0] _GEN_15862 = 14'h3df6 == index ? 14'h85 : _GEN_15861;
  wire [13:0] _GEN_15863 = 14'h3df7 == index ? 14'h84 : _GEN_15862;
  wire [13:0] _GEN_15864 = 14'h3df8 == index ? 14'h83 : _GEN_15863;
  wire [13:0] _GEN_15865 = 14'h3df9 == index ? 14'h82 : _GEN_15864;
  wire [13:0] _GEN_15866 = 14'h3dfa == index ? 14'h81 : _GEN_15865;
  wire [13:0] _GEN_15867 = 14'h3dfb == index ? 14'h80 : _GEN_15866;
  wire [13:0] _GEN_15868 = 14'h3dfc == index ? 14'h7b : _GEN_15867;
  wire [13:0] _GEN_15869 = 14'h3dfd == index ? 14'h7b : _GEN_15868;
  wire [13:0] _GEN_15870 = 14'h3dfe == index ? 14'h7b : _GEN_15869;
  wire [13:0] _GEN_15871 = 14'h3dff == index ? 14'h7b : _GEN_15870;
  wire [13:0] _GEN_15872 = 14'h3e00 == index ? 14'h0 : _GEN_15871;
  wire [13:0] _GEN_15873 = 14'h3e01 == index ? 14'h3e00 : _GEN_15872;
  wire [13:0] _GEN_15874 = 14'h3e02 == index ? 14'h1f00 : _GEN_15873;
  wire [13:0] _GEN_15875 = 14'h3e03 == index ? 14'h1481 : _GEN_15874;
  wire [13:0] _GEN_15876 = 14'h3e04 == index ? 14'hf80 : _GEN_15875;
  wire [13:0] _GEN_15877 = 14'h3e05 == index ? 14'hc04 : _GEN_15876;
  wire [13:0] _GEN_15878 = 14'h3e06 == index ? 14'ha04 : _GEN_15877;
  wire [13:0] _GEN_15879 = 14'h3e07 == index ? 14'h885 : _GEN_15878;
  wire [13:0] _GEN_15880 = 14'h3e08 == index ? 14'h784 : _GEN_15879;
  wire [13:0] _GEN_15881 = 14'h3e09 == index ? 14'h687 : _GEN_15880;
  wire [13:0] _GEN_15882 = 14'h3e0a == index ? 14'h604 : _GEN_15881;
  wire [13:0] _GEN_15883 = 14'h3e0b == index ? 14'h583 : _GEN_15882;
  wire [13:0] _GEN_15884 = 14'h3e0c == index ? 14'h504 : _GEN_15883;
  wire [13:0] _GEN_15885 = 14'h3e0d == index ? 14'h487 : _GEN_15884;
  wire [13:0] _GEN_15886 = 14'h3e0e == index ? 14'h40c : _GEN_15885;
  wire [13:0] _GEN_15887 = 14'h3e0f == index ? 14'h404 : _GEN_15886;
  wire [13:0] _GEN_15888 = 14'h3e10 == index ? 14'h38c : _GEN_15887;
  wire [13:0] _GEN_15889 = 14'h3e11 == index ? 14'h385 : _GEN_15888;
  wire [13:0] _GEN_15890 = 14'h3e12 == index ? 14'h310 : _GEN_15889;
  wire [13:0] _GEN_15891 = 14'h3e13 == index ? 14'h30a : _GEN_15890;
  wire [13:0] _GEN_15892 = 14'h3e14 == index ? 14'h304 : _GEN_15891;
  wire [13:0] _GEN_15893 = 14'h3e15 == index ? 14'h293 : _GEN_15892;
  wire [13:0] _GEN_15894 = 14'h3e16 == index ? 14'h28e : _GEN_15893;
  wire [13:0] _GEN_15895 = 14'h3e17 == index ? 14'h289 : _GEN_15894;
  wire [13:0] _GEN_15896 = 14'h3e18 == index ? 14'h284 : _GEN_15895;
  wire [13:0] _GEN_15897 = 14'h3e19 == index ? 14'h218 : _GEN_15896;
  wire [13:0] _GEN_15898 = 14'h3e1a == index ? 14'h214 : _GEN_15897;
  wire [13:0] _GEN_15899 = 14'h3e1b == index ? 14'h210 : _GEN_15898;
  wire [13:0] _GEN_15900 = 14'h3e1c == index ? 14'h20c : _GEN_15899;
  wire [13:0] _GEN_15901 = 14'h3e1d == index ? 14'h208 : _GEN_15900;
  wire [13:0] _GEN_15902 = 14'h3e1e == index ? 14'h204 : _GEN_15901;
  wire [13:0] _GEN_15903 = 14'h3e1f == index ? 14'h200 : _GEN_15902;
  wire [13:0] _GEN_15904 = 14'h3e20 == index ? 14'h19c : _GEN_15903;
  wire [13:0] _GEN_15905 = 14'h3e21 == index ? 14'h199 : _GEN_15904;
  wire [13:0] _GEN_15906 = 14'h3e22 == index ? 14'h196 : _GEN_15905;
  wire [13:0] _GEN_15907 = 14'h3e23 == index ? 14'h193 : _GEN_15906;
  wire [13:0] _GEN_15908 = 14'h3e24 == index ? 14'h190 : _GEN_15907;
  wire [13:0] _GEN_15909 = 14'h3e25 == index ? 14'h18d : _GEN_15908;
  wire [13:0] _GEN_15910 = 14'h3e26 == index ? 14'h18a : _GEN_15909;
  wire [13:0] _GEN_15911 = 14'h3e27 == index ? 14'h187 : _GEN_15910;
  wire [13:0] _GEN_15912 = 14'h3e28 == index ? 14'h184 : _GEN_15911;
  wire [13:0] _GEN_15913 = 14'h3e29 == index ? 14'h181 : _GEN_15912;
  wire [13:0] _GEN_15914 = 14'h3e2a == index ? 14'h128 : _GEN_15913;
  wire [13:0] _GEN_15915 = 14'h3e2b == index ? 14'h126 : _GEN_15914;
  wire [13:0] _GEN_15916 = 14'h3e2c == index ? 14'h124 : _GEN_15915;
  wire [13:0] _GEN_15917 = 14'h3e2d == index ? 14'h122 : _GEN_15916;
  wire [13:0] _GEN_15918 = 14'h3e2e == index ? 14'h120 : _GEN_15917;
  wire [13:0] _GEN_15919 = 14'h3e2f == index ? 14'h11e : _GEN_15918;
  wire [13:0] _GEN_15920 = 14'h3e30 == index ? 14'h11c : _GEN_15919;
  wire [13:0] _GEN_15921 = 14'h3e31 == index ? 14'h11a : _GEN_15920;
  wire [13:0] _GEN_15922 = 14'h3e32 == index ? 14'h118 : _GEN_15921;
  wire [13:0] _GEN_15923 = 14'h3e33 == index ? 14'h116 : _GEN_15922;
  wire [13:0] _GEN_15924 = 14'h3e34 == index ? 14'h114 : _GEN_15923;
  wire [13:0] _GEN_15925 = 14'h3e35 == index ? 14'h112 : _GEN_15924;
  wire [13:0] _GEN_15926 = 14'h3e36 == index ? 14'h110 : _GEN_15925;
  wire [13:0] _GEN_15927 = 14'h3e37 == index ? 14'h10e : _GEN_15926;
  wire [13:0] _GEN_15928 = 14'h3e38 == index ? 14'h10c : _GEN_15927;
  wire [13:0] _GEN_15929 = 14'h3e39 == index ? 14'h10a : _GEN_15928;
  wire [13:0] _GEN_15930 = 14'h3e3a == index ? 14'h108 : _GEN_15929;
  wire [13:0] _GEN_15931 = 14'h3e3b == index ? 14'h106 : _GEN_15930;
  wire [13:0] _GEN_15932 = 14'h3e3c == index ? 14'h104 : _GEN_15931;
  wire [13:0] _GEN_15933 = 14'h3e3d == index ? 14'h102 : _GEN_15932;
  wire [13:0] _GEN_15934 = 14'h3e3e == index ? 14'h100 : _GEN_15933;
  wire [13:0] _GEN_15935 = 14'h3e3f == index ? 14'hbd : _GEN_15934;
  wire [13:0] _GEN_15936 = 14'h3e40 == index ? 14'hbc : _GEN_15935;
  wire [13:0] _GEN_15937 = 14'h3e41 == index ? 14'hbb : _GEN_15936;
  wire [13:0] _GEN_15938 = 14'h3e42 == index ? 14'hba : _GEN_15937;
  wire [13:0] _GEN_15939 = 14'h3e43 == index ? 14'hb9 : _GEN_15938;
  wire [13:0] _GEN_15940 = 14'h3e44 == index ? 14'hb8 : _GEN_15939;
  wire [13:0] _GEN_15941 = 14'h3e45 == index ? 14'hb7 : _GEN_15940;
  wire [13:0] _GEN_15942 = 14'h3e46 == index ? 14'hb6 : _GEN_15941;
  wire [13:0] _GEN_15943 = 14'h3e47 == index ? 14'hb5 : _GEN_15942;
  wire [13:0] _GEN_15944 = 14'h3e48 == index ? 14'hb4 : _GEN_15943;
  wire [13:0] _GEN_15945 = 14'h3e49 == index ? 14'hb3 : _GEN_15944;
  wire [13:0] _GEN_15946 = 14'h3e4a == index ? 14'hb2 : _GEN_15945;
  wire [13:0] _GEN_15947 = 14'h3e4b == index ? 14'hb1 : _GEN_15946;
  wire [13:0] _GEN_15948 = 14'h3e4c == index ? 14'hb0 : _GEN_15947;
  wire [13:0] _GEN_15949 = 14'h3e4d == index ? 14'haf : _GEN_15948;
  wire [13:0] _GEN_15950 = 14'h3e4e == index ? 14'hae : _GEN_15949;
  wire [13:0] _GEN_15951 = 14'h3e4f == index ? 14'had : _GEN_15950;
  wire [13:0] _GEN_15952 = 14'h3e50 == index ? 14'hac : _GEN_15951;
  wire [13:0] _GEN_15953 = 14'h3e51 == index ? 14'hab : _GEN_15952;
  wire [13:0] _GEN_15954 = 14'h3e52 == index ? 14'haa : _GEN_15953;
  wire [13:0] _GEN_15955 = 14'h3e53 == index ? 14'ha9 : _GEN_15954;
  wire [13:0] _GEN_15956 = 14'h3e54 == index ? 14'ha8 : _GEN_15955;
  wire [13:0] _GEN_15957 = 14'h3e55 == index ? 14'ha7 : _GEN_15956;
  wire [13:0] _GEN_15958 = 14'h3e56 == index ? 14'ha6 : _GEN_15957;
  wire [13:0] _GEN_15959 = 14'h3e57 == index ? 14'ha5 : _GEN_15958;
  wire [13:0] _GEN_15960 = 14'h3e58 == index ? 14'ha4 : _GEN_15959;
  wire [13:0] _GEN_15961 = 14'h3e59 == index ? 14'ha3 : _GEN_15960;
  wire [13:0] _GEN_15962 = 14'h3e5a == index ? 14'ha2 : _GEN_15961;
  wire [13:0] _GEN_15963 = 14'h3e5b == index ? 14'ha1 : _GEN_15962;
  wire [13:0] _GEN_15964 = 14'h3e5c == index ? 14'ha0 : _GEN_15963;
  wire [13:0] _GEN_15965 = 14'h3e5d == index ? 14'h9f : _GEN_15964;
  wire [13:0] _GEN_15966 = 14'h3e5e == index ? 14'h9e : _GEN_15965;
  wire [13:0] _GEN_15967 = 14'h3e5f == index ? 14'h9d : _GEN_15966;
  wire [13:0] _GEN_15968 = 14'h3e60 == index ? 14'h9c : _GEN_15967;
  wire [13:0] _GEN_15969 = 14'h3e61 == index ? 14'h9b : _GEN_15968;
  wire [13:0] _GEN_15970 = 14'h3e62 == index ? 14'h9a : _GEN_15969;
  wire [13:0] _GEN_15971 = 14'h3e63 == index ? 14'h99 : _GEN_15970;
  wire [13:0] _GEN_15972 = 14'h3e64 == index ? 14'h98 : _GEN_15971;
  wire [13:0] _GEN_15973 = 14'h3e65 == index ? 14'h97 : _GEN_15972;
  wire [13:0] _GEN_15974 = 14'h3e66 == index ? 14'h96 : _GEN_15973;
  wire [13:0] _GEN_15975 = 14'h3e67 == index ? 14'h95 : _GEN_15974;
  wire [13:0] _GEN_15976 = 14'h3e68 == index ? 14'h94 : _GEN_15975;
  wire [13:0] _GEN_15977 = 14'h3e69 == index ? 14'h93 : _GEN_15976;
  wire [13:0] _GEN_15978 = 14'h3e6a == index ? 14'h92 : _GEN_15977;
  wire [13:0] _GEN_15979 = 14'h3e6b == index ? 14'h91 : _GEN_15978;
  wire [13:0] _GEN_15980 = 14'h3e6c == index ? 14'h90 : _GEN_15979;
  wire [13:0] _GEN_15981 = 14'h3e6d == index ? 14'h8f : _GEN_15980;
  wire [13:0] _GEN_15982 = 14'h3e6e == index ? 14'h8e : _GEN_15981;
  wire [13:0] _GEN_15983 = 14'h3e6f == index ? 14'h8d : _GEN_15982;
  wire [13:0] _GEN_15984 = 14'h3e70 == index ? 14'h8c : _GEN_15983;
  wire [13:0] _GEN_15985 = 14'h3e71 == index ? 14'h8b : _GEN_15984;
  wire [13:0] _GEN_15986 = 14'h3e72 == index ? 14'h8a : _GEN_15985;
  wire [13:0] _GEN_15987 = 14'h3e73 == index ? 14'h89 : _GEN_15986;
  wire [13:0] _GEN_15988 = 14'h3e74 == index ? 14'h88 : _GEN_15987;
  wire [13:0] _GEN_15989 = 14'h3e75 == index ? 14'h87 : _GEN_15988;
  wire [13:0] _GEN_15990 = 14'h3e76 == index ? 14'h86 : _GEN_15989;
  wire [13:0] _GEN_15991 = 14'h3e77 == index ? 14'h85 : _GEN_15990;
  wire [13:0] _GEN_15992 = 14'h3e78 == index ? 14'h84 : _GEN_15991;
  wire [13:0] _GEN_15993 = 14'h3e79 == index ? 14'h83 : _GEN_15992;
  wire [13:0] _GEN_15994 = 14'h3e7a == index ? 14'h82 : _GEN_15993;
  wire [13:0] _GEN_15995 = 14'h3e7b == index ? 14'h81 : _GEN_15994;
  wire [13:0] _GEN_15996 = 14'h3e7c == index ? 14'h80 : _GEN_15995;
  wire [13:0] _GEN_15997 = 14'h3e7d == index ? 14'h7c : _GEN_15996;
  wire [13:0] _GEN_15998 = 14'h3e7e == index ? 14'h7c : _GEN_15997;
  wire [13:0] _GEN_15999 = 14'h3e7f == index ? 14'h7c : _GEN_15998;
  wire [13:0] _GEN_16000 = 14'h3e80 == index ? 14'h0 : _GEN_15999;
  wire [13:0] _GEN_16001 = 14'h3e81 == index ? 14'h3e80 : _GEN_16000;
  wire [13:0] _GEN_16002 = 14'h3e82 == index ? 14'h1f01 : _GEN_16001;
  wire [13:0] _GEN_16003 = 14'h3e83 == index ? 14'h1482 : _GEN_16002;
  wire [13:0] _GEN_16004 = 14'h3e84 == index ? 14'hf81 : _GEN_16003;
  wire [13:0] _GEN_16005 = 14'h3e85 == index ? 14'hc80 : _GEN_16004;
  wire [13:0] _GEN_16006 = 14'h3e86 == index ? 14'ha05 : _GEN_16005;
  wire [13:0] _GEN_16007 = 14'h3e87 == index ? 14'h886 : _GEN_16006;
  wire [13:0] _GEN_16008 = 14'h3e88 == index ? 14'h785 : _GEN_16007;
  wire [13:0] _GEN_16009 = 14'h3e89 == index ? 14'h688 : _GEN_16008;
  wire [13:0] _GEN_16010 = 14'h3e8a == index ? 14'h605 : _GEN_16009;
  wire [13:0] _GEN_16011 = 14'h3e8b == index ? 14'h584 : _GEN_16010;
  wire [13:0] _GEN_16012 = 14'h3e8c == index ? 14'h505 : _GEN_16011;
  wire [13:0] _GEN_16013 = 14'h3e8d == index ? 14'h488 : _GEN_16012;
  wire [13:0] _GEN_16014 = 14'h3e8e == index ? 14'h40d : _GEN_16013;
  wire [13:0] _GEN_16015 = 14'h3e8f == index ? 14'h405 : _GEN_16014;
  wire [13:0] _GEN_16016 = 14'h3e90 == index ? 14'h38d : _GEN_16015;
  wire [13:0] _GEN_16017 = 14'h3e91 == index ? 14'h386 : _GEN_16016;
  wire [13:0] _GEN_16018 = 14'h3e92 == index ? 14'h311 : _GEN_16017;
  wire [13:0] _GEN_16019 = 14'h3e93 == index ? 14'h30b : _GEN_16018;
  wire [13:0] _GEN_16020 = 14'h3e94 == index ? 14'h305 : _GEN_16019;
  wire [13:0] _GEN_16021 = 14'h3e95 == index ? 14'h294 : _GEN_16020;
  wire [13:0] _GEN_16022 = 14'h3e96 == index ? 14'h28f : _GEN_16021;
  wire [13:0] _GEN_16023 = 14'h3e97 == index ? 14'h28a : _GEN_16022;
  wire [13:0] _GEN_16024 = 14'h3e98 == index ? 14'h285 : _GEN_16023;
  wire [13:0] _GEN_16025 = 14'h3e99 == index ? 14'h280 : _GEN_16024;
  wire [13:0] _GEN_16026 = 14'h3e9a == index ? 14'h215 : _GEN_16025;
  wire [13:0] _GEN_16027 = 14'h3e9b == index ? 14'h211 : _GEN_16026;
  wire [13:0] _GEN_16028 = 14'h3e9c == index ? 14'h20d : _GEN_16027;
  wire [13:0] _GEN_16029 = 14'h3e9d == index ? 14'h209 : _GEN_16028;
  wire [13:0] _GEN_16030 = 14'h3e9e == index ? 14'h205 : _GEN_16029;
  wire [13:0] _GEN_16031 = 14'h3e9f == index ? 14'h201 : _GEN_16030;
  wire [13:0] _GEN_16032 = 14'h3ea0 == index ? 14'h19d : _GEN_16031;
  wire [13:0] _GEN_16033 = 14'h3ea1 == index ? 14'h19a : _GEN_16032;
  wire [13:0] _GEN_16034 = 14'h3ea2 == index ? 14'h197 : _GEN_16033;
  wire [13:0] _GEN_16035 = 14'h3ea3 == index ? 14'h194 : _GEN_16034;
  wire [13:0] _GEN_16036 = 14'h3ea4 == index ? 14'h191 : _GEN_16035;
  wire [13:0] _GEN_16037 = 14'h3ea5 == index ? 14'h18e : _GEN_16036;
  wire [13:0] _GEN_16038 = 14'h3ea6 == index ? 14'h18b : _GEN_16037;
  wire [13:0] _GEN_16039 = 14'h3ea7 == index ? 14'h188 : _GEN_16038;
  wire [13:0] _GEN_16040 = 14'h3ea8 == index ? 14'h185 : _GEN_16039;
  wire [13:0] _GEN_16041 = 14'h3ea9 == index ? 14'h182 : _GEN_16040;
  wire [13:0] _GEN_16042 = 14'h3eaa == index ? 14'h129 : _GEN_16041;
  wire [13:0] _GEN_16043 = 14'h3eab == index ? 14'h127 : _GEN_16042;
  wire [13:0] _GEN_16044 = 14'h3eac == index ? 14'h125 : _GEN_16043;
  wire [13:0] _GEN_16045 = 14'h3ead == index ? 14'h123 : _GEN_16044;
  wire [13:0] _GEN_16046 = 14'h3eae == index ? 14'h121 : _GEN_16045;
  wire [13:0] _GEN_16047 = 14'h3eaf == index ? 14'h11f : _GEN_16046;
  wire [13:0] _GEN_16048 = 14'h3eb0 == index ? 14'h11d : _GEN_16047;
  wire [13:0] _GEN_16049 = 14'h3eb1 == index ? 14'h11b : _GEN_16048;
  wire [13:0] _GEN_16050 = 14'h3eb2 == index ? 14'h119 : _GEN_16049;
  wire [13:0] _GEN_16051 = 14'h3eb3 == index ? 14'h117 : _GEN_16050;
  wire [13:0] _GEN_16052 = 14'h3eb4 == index ? 14'h115 : _GEN_16051;
  wire [13:0] _GEN_16053 = 14'h3eb5 == index ? 14'h113 : _GEN_16052;
  wire [13:0] _GEN_16054 = 14'h3eb6 == index ? 14'h111 : _GEN_16053;
  wire [13:0] _GEN_16055 = 14'h3eb7 == index ? 14'h10f : _GEN_16054;
  wire [13:0] _GEN_16056 = 14'h3eb8 == index ? 14'h10d : _GEN_16055;
  wire [13:0] _GEN_16057 = 14'h3eb9 == index ? 14'h10b : _GEN_16056;
  wire [13:0] _GEN_16058 = 14'h3eba == index ? 14'h109 : _GEN_16057;
  wire [13:0] _GEN_16059 = 14'h3ebb == index ? 14'h107 : _GEN_16058;
  wire [13:0] _GEN_16060 = 14'h3ebc == index ? 14'h105 : _GEN_16059;
  wire [13:0] _GEN_16061 = 14'h3ebd == index ? 14'h103 : _GEN_16060;
  wire [13:0] _GEN_16062 = 14'h3ebe == index ? 14'h101 : _GEN_16061;
  wire [13:0] _GEN_16063 = 14'h3ebf == index ? 14'hbe : _GEN_16062;
  wire [13:0] _GEN_16064 = 14'h3ec0 == index ? 14'hbd : _GEN_16063;
  wire [13:0] _GEN_16065 = 14'h3ec1 == index ? 14'hbc : _GEN_16064;
  wire [13:0] _GEN_16066 = 14'h3ec2 == index ? 14'hbb : _GEN_16065;
  wire [13:0] _GEN_16067 = 14'h3ec3 == index ? 14'hba : _GEN_16066;
  wire [13:0] _GEN_16068 = 14'h3ec4 == index ? 14'hb9 : _GEN_16067;
  wire [13:0] _GEN_16069 = 14'h3ec5 == index ? 14'hb8 : _GEN_16068;
  wire [13:0] _GEN_16070 = 14'h3ec6 == index ? 14'hb7 : _GEN_16069;
  wire [13:0] _GEN_16071 = 14'h3ec7 == index ? 14'hb6 : _GEN_16070;
  wire [13:0] _GEN_16072 = 14'h3ec8 == index ? 14'hb5 : _GEN_16071;
  wire [13:0] _GEN_16073 = 14'h3ec9 == index ? 14'hb4 : _GEN_16072;
  wire [13:0] _GEN_16074 = 14'h3eca == index ? 14'hb3 : _GEN_16073;
  wire [13:0] _GEN_16075 = 14'h3ecb == index ? 14'hb2 : _GEN_16074;
  wire [13:0] _GEN_16076 = 14'h3ecc == index ? 14'hb1 : _GEN_16075;
  wire [13:0] _GEN_16077 = 14'h3ecd == index ? 14'hb0 : _GEN_16076;
  wire [13:0] _GEN_16078 = 14'h3ece == index ? 14'haf : _GEN_16077;
  wire [13:0] _GEN_16079 = 14'h3ecf == index ? 14'hae : _GEN_16078;
  wire [13:0] _GEN_16080 = 14'h3ed0 == index ? 14'had : _GEN_16079;
  wire [13:0] _GEN_16081 = 14'h3ed1 == index ? 14'hac : _GEN_16080;
  wire [13:0] _GEN_16082 = 14'h3ed2 == index ? 14'hab : _GEN_16081;
  wire [13:0] _GEN_16083 = 14'h3ed3 == index ? 14'haa : _GEN_16082;
  wire [13:0] _GEN_16084 = 14'h3ed4 == index ? 14'ha9 : _GEN_16083;
  wire [13:0] _GEN_16085 = 14'h3ed5 == index ? 14'ha8 : _GEN_16084;
  wire [13:0] _GEN_16086 = 14'h3ed6 == index ? 14'ha7 : _GEN_16085;
  wire [13:0] _GEN_16087 = 14'h3ed7 == index ? 14'ha6 : _GEN_16086;
  wire [13:0] _GEN_16088 = 14'h3ed8 == index ? 14'ha5 : _GEN_16087;
  wire [13:0] _GEN_16089 = 14'h3ed9 == index ? 14'ha4 : _GEN_16088;
  wire [13:0] _GEN_16090 = 14'h3eda == index ? 14'ha3 : _GEN_16089;
  wire [13:0] _GEN_16091 = 14'h3edb == index ? 14'ha2 : _GEN_16090;
  wire [13:0] _GEN_16092 = 14'h3edc == index ? 14'ha1 : _GEN_16091;
  wire [13:0] _GEN_16093 = 14'h3edd == index ? 14'ha0 : _GEN_16092;
  wire [13:0] _GEN_16094 = 14'h3ede == index ? 14'h9f : _GEN_16093;
  wire [13:0] _GEN_16095 = 14'h3edf == index ? 14'h9e : _GEN_16094;
  wire [13:0] _GEN_16096 = 14'h3ee0 == index ? 14'h9d : _GEN_16095;
  wire [13:0] _GEN_16097 = 14'h3ee1 == index ? 14'h9c : _GEN_16096;
  wire [13:0] _GEN_16098 = 14'h3ee2 == index ? 14'h9b : _GEN_16097;
  wire [13:0] _GEN_16099 = 14'h3ee3 == index ? 14'h9a : _GEN_16098;
  wire [13:0] _GEN_16100 = 14'h3ee4 == index ? 14'h99 : _GEN_16099;
  wire [13:0] _GEN_16101 = 14'h3ee5 == index ? 14'h98 : _GEN_16100;
  wire [13:0] _GEN_16102 = 14'h3ee6 == index ? 14'h97 : _GEN_16101;
  wire [13:0] _GEN_16103 = 14'h3ee7 == index ? 14'h96 : _GEN_16102;
  wire [13:0] _GEN_16104 = 14'h3ee8 == index ? 14'h95 : _GEN_16103;
  wire [13:0] _GEN_16105 = 14'h3ee9 == index ? 14'h94 : _GEN_16104;
  wire [13:0] _GEN_16106 = 14'h3eea == index ? 14'h93 : _GEN_16105;
  wire [13:0] _GEN_16107 = 14'h3eeb == index ? 14'h92 : _GEN_16106;
  wire [13:0] _GEN_16108 = 14'h3eec == index ? 14'h91 : _GEN_16107;
  wire [13:0] _GEN_16109 = 14'h3eed == index ? 14'h90 : _GEN_16108;
  wire [13:0] _GEN_16110 = 14'h3eee == index ? 14'h8f : _GEN_16109;
  wire [13:0] _GEN_16111 = 14'h3eef == index ? 14'h8e : _GEN_16110;
  wire [13:0] _GEN_16112 = 14'h3ef0 == index ? 14'h8d : _GEN_16111;
  wire [13:0] _GEN_16113 = 14'h3ef1 == index ? 14'h8c : _GEN_16112;
  wire [13:0] _GEN_16114 = 14'h3ef2 == index ? 14'h8b : _GEN_16113;
  wire [13:0] _GEN_16115 = 14'h3ef3 == index ? 14'h8a : _GEN_16114;
  wire [13:0] _GEN_16116 = 14'h3ef4 == index ? 14'h89 : _GEN_16115;
  wire [13:0] _GEN_16117 = 14'h3ef5 == index ? 14'h88 : _GEN_16116;
  wire [13:0] _GEN_16118 = 14'h3ef6 == index ? 14'h87 : _GEN_16117;
  wire [13:0] _GEN_16119 = 14'h3ef7 == index ? 14'h86 : _GEN_16118;
  wire [13:0] _GEN_16120 = 14'h3ef8 == index ? 14'h85 : _GEN_16119;
  wire [13:0] _GEN_16121 = 14'h3ef9 == index ? 14'h84 : _GEN_16120;
  wire [13:0] _GEN_16122 = 14'h3efa == index ? 14'h83 : _GEN_16121;
  wire [13:0] _GEN_16123 = 14'h3efb == index ? 14'h82 : _GEN_16122;
  wire [13:0] _GEN_16124 = 14'h3efc == index ? 14'h81 : _GEN_16123;
  wire [13:0] _GEN_16125 = 14'h3efd == index ? 14'h80 : _GEN_16124;
  wire [13:0] _GEN_16126 = 14'h3efe == index ? 14'h7d : _GEN_16125;
  wire [13:0] _GEN_16127 = 14'h3eff == index ? 14'h7d : _GEN_16126;
  wire [13:0] _GEN_16128 = 14'h3f00 == index ? 14'h0 : _GEN_16127;
  wire [13:0] _GEN_16129 = 14'h3f01 == index ? 14'h3f00 : _GEN_16128;
  wire [13:0] _GEN_16130 = 14'h3f02 == index ? 14'h1f80 : _GEN_16129;
  wire [13:0] _GEN_16131 = 14'h3f03 == index ? 14'h1500 : _GEN_16130;
  wire [13:0] _GEN_16132 = 14'h3f04 == index ? 14'hf82 : _GEN_16131;
  wire [13:0] _GEN_16133 = 14'h3f05 == index ? 14'hc81 : _GEN_16132;
  wire [13:0] _GEN_16134 = 14'h3f06 == index ? 14'ha80 : _GEN_16133;
  wire [13:0] _GEN_16135 = 14'h3f07 == index ? 14'h900 : _GEN_16134;
  wire [13:0] _GEN_16136 = 14'h3f08 == index ? 14'h786 : _GEN_16135;
  wire [13:0] _GEN_16137 = 14'h3f09 == index ? 14'h700 : _GEN_16136;
  wire [13:0] _GEN_16138 = 14'h3f0a == index ? 14'h606 : _GEN_16137;
  wire [13:0] _GEN_16139 = 14'h3f0b == index ? 14'h585 : _GEN_16138;
  wire [13:0] _GEN_16140 = 14'h3f0c == index ? 14'h506 : _GEN_16139;
  wire [13:0] _GEN_16141 = 14'h3f0d == index ? 14'h489 : _GEN_16140;
  wire [13:0] _GEN_16142 = 14'h3f0e == index ? 14'h480 : _GEN_16141;
  wire [13:0] _GEN_16143 = 14'h3f0f == index ? 14'h406 : _GEN_16142;
  wire [13:0] _GEN_16144 = 14'h3f10 == index ? 14'h38e : _GEN_16143;
  wire [13:0] _GEN_16145 = 14'h3f11 == index ? 14'h387 : _GEN_16144;
  wire [13:0] _GEN_16146 = 14'h3f12 == index ? 14'h380 : _GEN_16145;
  wire [13:0] _GEN_16147 = 14'h3f13 == index ? 14'h30c : _GEN_16146;
  wire [13:0] _GEN_16148 = 14'h3f14 == index ? 14'h306 : _GEN_16147;
  wire [13:0] _GEN_16149 = 14'h3f15 == index ? 14'h300 : _GEN_16148;
  wire [13:0] _GEN_16150 = 14'h3f16 == index ? 14'h290 : _GEN_16149;
  wire [13:0] _GEN_16151 = 14'h3f17 == index ? 14'h28b : _GEN_16150;
  wire [13:0] _GEN_16152 = 14'h3f18 == index ? 14'h286 : _GEN_16151;
  wire [13:0] _GEN_16153 = 14'h3f19 == index ? 14'h281 : _GEN_16152;
  wire [13:0] _GEN_16154 = 14'h3f1a == index ? 14'h216 : _GEN_16153;
  wire [13:0] _GEN_16155 = 14'h3f1b == index ? 14'h212 : _GEN_16154;
  wire [13:0] _GEN_16156 = 14'h3f1c == index ? 14'h20e : _GEN_16155;
  wire [13:0] _GEN_16157 = 14'h3f1d == index ? 14'h20a : _GEN_16156;
  wire [13:0] _GEN_16158 = 14'h3f1e == index ? 14'h206 : _GEN_16157;
  wire [13:0] _GEN_16159 = 14'h3f1f == index ? 14'h202 : _GEN_16158;
  wire [13:0] _GEN_16160 = 14'h3f20 == index ? 14'h19e : _GEN_16159;
  wire [13:0] _GEN_16161 = 14'h3f21 == index ? 14'h19b : _GEN_16160;
  wire [13:0] _GEN_16162 = 14'h3f22 == index ? 14'h198 : _GEN_16161;
  wire [13:0] _GEN_16163 = 14'h3f23 == index ? 14'h195 : _GEN_16162;
  wire [13:0] _GEN_16164 = 14'h3f24 == index ? 14'h192 : _GEN_16163;
  wire [13:0] _GEN_16165 = 14'h3f25 == index ? 14'h18f : _GEN_16164;
  wire [13:0] _GEN_16166 = 14'h3f26 == index ? 14'h18c : _GEN_16165;
  wire [13:0] _GEN_16167 = 14'h3f27 == index ? 14'h189 : _GEN_16166;
  wire [13:0] _GEN_16168 = 14'h3f28 == index ? 14'h186 : _GEN_16167;
  wire [13:0] _GEN_16169 = 14'h3f29 == index ? 14'h183 : _GEN_16168;
  wire [13:0] _GEN_16170 = 14'h3f2a == index ? 14'h180 : _GEN_16169;
  wire [13:0] _GEN_16171 = 14'h3f2b == index ? 14'h128 : _GEN_16170;
  wire [13:0] _GEN_16172 = 14'h3f2c == index ? 14'h126 : _GEN_16171;
  wire [13:0] _GEN_16173 = 14'h3f2d == index ? 14'h124 : _GEN_16172;
  wire [13:0] _GEN_16174 = 14'h3f2e == index ? 14'h122 : _GEN_16173;
  wire [13:0] _GEN_16175 = 14'h3f2f == index ? 14'h120 : _GEN_16174;
  wire [13:0] _GEN_16176 = 14'h3f30 == index ? 14'h11e : _GEN_16175;
  wire [13:0] _GEN_16177 = 14'h3f31 == index ? 14'h11c : _GEN_16176;
  wire [13:0] _GEN_16178 = 14'h3f32 == index ? 14'h11a : _GEN_16177;
  wire [13:0] _GEN_16179 = 14'h3f33 == index ? 14'h118 : _GEN_16178;
  wire [13:0] _GEN_16180 = 14'h3f34 == index ? 14'h116 : _GEN_16179;
  wire [13:0] _GEN_16181 = 14'h3f35 == index ? 14'h114 : _GEN_16180;
  wire [13:0] _GEN_16182 = 14'h3f36 == index ? 14'h112 : _GEN_16181;
  wire [13:0] _GEN_16183 = 14'h3f37 == index ? 14'h110 : _GEN_16182;
  wire [13:0] _GEN_16184 = 14'h3f38 == index ? 14'h10e : _GEN_16183;
  wire [13:0] _GEN_16185 = 14'h3f39 == index ? 14'h10c : _GEN_16184;
  wire [13:0] _GEN_16186 = 14'h3f3a == index ? 14'h10a : _GEN_16185;
  wire [13:0] _GEN_16187 = 14'h3f3b == index ? 14'h108 : _GEN_16186;
  wire [13:0] _GEN_16188 = 14'h3f3c == index ? 14'h106 : _GEN_16187;
  wire [13:0] _GEN_16189 = 14'h3f3d == index ? 14'h104 : _GEN_16188;
  wire [13:0] _GEN_16190 = 14'h3f3e == index ? 14'h102 : _GEN_16189;
  wire [13:0] _GEN_16191 = 14'h3f3f == index ? 14'h100 : _GEN_16190;
  wire [13:0] _GEN_16192 = 14'h3f40 == index ? 14'hbe : _GEN_16191;
  wire [13:0] _GEN_16193 = 14'h3f41 == index ? 14'hbd : _GEN_16192;
  wire [13:0] _GEN_16194 = 14'h3f42 == index ? 14'hbc : _GEN_16193;
  wire [13:0] _GEN_16195 = 14'h3f43 == index ? 14'hbb : _GEN_16194;
  wire [13:0] _GEN_16196 = 14'h3f44 == index ? 14'hba : _GEN_16195;
  wire [13:0] _GEN_16197 = 14'h3f45 == index ? 14'hb9 : _GEN_16196;
  wire [13:0] _GEN_16198 = 14'h3f46 == index ? 14'hb8 : _GEN_16197;
  wire [13:0] _GEN_16199 = 14'h3f47 == index ? 14'hb7 : _GEN_16198;
  wire [13:0] _GEN_16200 = 14'h3f48 == index ? 14'hb6 : _GEN_16199;
  wire [13:0] _GEN_16201 = 14'h3f49 == index ? 14'hb5 : _GEN_16200;
  wire [13:0] _GEN_16202 = 14'h3f4a == index ? 14'hb4 : _GEN_16201;
  wire [13:0] _GEN_16203 = 14'h3f4b == index ? 14'hb3 : _GEN_16202;
  wire [13:0] _GEN_16204 = 14'h3f4c == index ? 14'hb2 : _GEN_16203;
  wire [13:0] _GEN_16205 = 14'h3f4d == index ? 14'hb1 : _GEN_16204;
  wire [13:0] _GEN_16206 = 14'h3f4e == index ? 14'hb0 : _GEN_16205;
  wire [13:0] _GEN_16207 = 14'h3f4f == index ? 14'haf : _GEN_16206;
  wire [13:0] _GEN_16208 = 14'h3f50 == index ? 14'hae : _GEN_16207;
  wire [13:0] _GEN_16209 = 14'h3f51 == index ? 14'had : _GEN_16208;
  wire [13:0] _GEN_16210 = 14'h3f52 == index ? 14'hac : _GEN_16209;
  wire [13:0] _GEN_16211 = 14'h3f53 == index ? 14'hab : _GEN_16210;
  wire [13:0] _GEN_16212 = 14'h3f54 == index ? 14'haa : _GEN_16211;
  wire [13:0] _GEN_16213 = 14'h3f55 == index ? 14'ha9 : _GEN_16212;
  wire [13:0] _GEN_16214 = 14'h3f56 == index ? 14'ha8 : _GEN_16213;
  wire [13:0] _GEN_16215 = 14'h3f57 == index ? 14'ha7 : _GEN_16214;
  wire [13:0] _GEN_16216 = 14'h3f58 == index ? 14'ha6 : _GEN_16215;
  wire [13:0] _GEN_16217 = 14'h3f59 == index ? 14'ha5 : _GEN_16216;
  wire [13:0] _GEN_16218 = 14'h3f5a == index ? 14'ha4 : _GEN_16217;
  wire [13:0] _GEN_16219 = 14'h3f5b == index ? 14'ha3 : _GEN_16218;
  wire [13:0] _GEN_16220 = 14'h3f5c == index ? 14'ha2 : _GEN_16219;
  wire [13:0] _GEN_16221 = 14'h3f5d == index ? 14'ha1 : _GEN_16220;
  wire [13:0] _GEN_16222 = 14'h3f5e == index ? 14'ha0 : _GEN_16221;
  wire [13:0] _GEN_16223 = 14'h3f5f == index ? 14'h9f : _GEN_16222;
  wire [13:0] _GEN_16224 = 14'h3f60 == index ? 14'h9e : _GEN_16223;
  wire [13:0] _GEN_16225 = 14'h3f61 == index ? 14'h9d : _GEN_16224;
  wire [13:0] _GEN_16226 = 14'h3f62 == index ? 14'h9c : _GEN_16225;
  wire [13:0] _GEN_16227 = 14'h3f63 == index ? 14'h9b : _GEN_16226;
  wire [13:0] _GEN_16228 = 14'h3f64 == index ? 14'h9a : _GEN_16227;
  wire [13:0] _GEN_16229 = 14'h3f65 == index ? 14'h99 : _GEN_16228;
  wire [13:0] _GEN_16230 = 14'h3f66 == index ? 14'h98 : _GEN_16229;
  wire [13:0] _GEN_16231 = 14'h3f67 == index ? 14'h97 : _GEN_16230;
  wire [13:0] _GEN_16232 = 14'h3f68 == index ? 14'h96 : _GEN_16231;
  wire [13:0] _GEN_16233 = 14'h3f69 == index ? 14'h95 : _GEN_16232;
  wire [13:0] _GEN_16234 = 14'h3f6a == index ? 14'h94 : _GEN_16233;
  wire [13:0] _GEN_16235 = 14'h3f6b == index ? 14'h93 : _GEN_16234;
  wire [13:0] _GEN_16236 = 14'h3f6c == index ? 14'h92 : _GEN_16235;
  wire [13:0] _GEN_16237 = 14'h3f6d == index ? 14'h91 : _GEN_16236;
  wire [13:0] _GEN_16238 = 14'h3f6e == index ? 14'h90 : _GEN_16237;
  wire [13:0] _GEN_16239 = 14'h3f6f == index ? 14'h8f : _GEN_16238;
  wire [13:0] _GEN_16240 = 14'h3f70 == index ? 14'h8e : _GEN_16239;
  wire [13:0] _GEN_16241 = 14'h3f71 == index ? 14'h8d : _GEN_16240;
  wire [13:0] _GEN_16242 = 14'h3f72 == index ? 14'h8c : _GEN_16241;
  wire [13:0] _GEN_16243 = 14'h3f73 == index ? 14'h8b : _GEN_16242;
  wire [13:0] _GEN_16244 = 14'h3f74 == index ? 14'h8a : _GEN_16243;
  wire [13:0] _GEN_16245 = 14'h3f75 == index ? 14'h89 : _GEN_16244;
  wire [13:0] _GEN_16246 = 14'h3f76 == index ? 14'h88 : _GEN_16245;
  wire [13:0] _GEN_16247 = 14'h3f77 == index ? 14'h87 : _GEN_16246;
  wire [13:0] _GEN_16248 = 14'h3f78 == index ? 14'h86 : _GEN_16247;
  wire [13:0] _GEN_16249 = 14'h3f79 == index ? 14'h85 : _GEN_16248;
  wire [13:0] _GEN_16250 = 14'h3f7a == index ? 14'h84 : _GEN_16249;
  wire [13:0] _GEN_16251 = 14'h3f7b == index ? 14'h83 : _GEN_16250;
  wire [13:0] _GEN_16252 = 14'h3f7c == index ? 14'h82 : _GEN_16251;
  wire [13:0] _GEN_16253 = 14'h3f7d == index ? 14'h81 : _GEN_16252;
  wire [13:0] _GEN_16254 = 14'h3f7e == index ? 14'h80 : _GEN_16253;
  wire [13:0] _GEN_16255 = 14'h3f7f == index ? 14'h7e : _GEN_16254;
  wire [13:0] _GEN_16256 = 14'h3f80 == index ? 14'h0 : _GEN_16255;
  wire [13:0] _GEN_16257 = 14'h3f81 == index ? 14'h3f80 : _GEN_16256;
  wire [13:0] _GEN_16258 = 14'h3f82 == index ? 14'h1f81 : _GEN_16257;
  wire [13:0] _GEN_16259 = 14'h3f83 == index ? 14'h1501 : _GEN_16258;
  wire [13:0] _GEN_16260 = 14'h3f84 == index ? 14'hf83 : _GEN_16259;
  wire [13:0] _GEN_16261 = 14'h3f85 == index ? 14'hc82 : _GEN_16260;
  wire [13:0] _GEN_16262 = 14'h3f86 == index ? 14'ha81 : _GEN_16261;
  wire [13:0] _GEN_16263 = 14'h3f87 == index ? 14'h901 : _GEN_16262;
  wire [13:0] _GEN_16264 = 14'h3f88 == index ? 14'h787 : _GEN_16263;
  wire [13:0] _GEN_16265 = 14'h3f89 == index ? 14'h701 : _GEN_16264;
  wire [13:0] _GEN_16266 = 14'h3f8a == index ? 14'h607 : _GEN_16265;
  wire [13:0] _GEN_16267 = 14'h3f8b == index ? 14'h586 : _GEN_16266;
  wire [13:0] _GEN_16268 = 14'h3f8c == index ? 14'h507 : _GEN_16267;
  wire [13:0] _GEN_16269 = 14'h3f8d == index ? 14'h48a : _GEN_16268;
  wire [13:0] _GEN_16270 = 14'h3f8e == index ? 14'h481 : _GEN_16269;
  wire [13:0] _GEN_16271 = 14'h3f8f == index ? 14'h407 : _GEN_16270;
  wire [13:0] _GEN_16272 = 14'h3f90 == index ? 14'h38f : _GEN_16271;
  wire [13:0] _GEN_16273 = 14'h3f91 == index ? 14'h388 : _GEN_16272;
  wire [13:0] _GEN_16274 = 14'h3f92 == index ? 14'h381 : _GEN_16273;
  wire [13:0] _GEN_16275 = 14'h3f93 == index ? 14'h30d : _GEN_16274;
  wire [13:0] _GEN_16276 = 14'h3f94 == index ? 14'h307 : _GEN_16275;
  wire [13:0] _GEN_16277 = 14'h3f95 == index ? 14'h301 : _GEN_16276;
  wire [13:0] _GEN_16278 = 14'h3f96 == index ? 14'h291 : _GEN_16277;
  wire [13:0] _GEN_16279 = 14'h3f97 == index ? 14'h28c : _GEN_16278;
  wire [13:0] _GEN_16280 = 14'h3f98 == index ? 14'h287 : _GEN_16279;
  wire [13:0] _GEN_16281 = 14'h3f99 == index ? 14'h282 : _GEN_16280;
  wire [13:0] _GEN_16282 = 14'h3f9a == index ? 14'h217 : _GEN_16281;
  wire [13:0] _GEN_16283 = 14'h3f9b == index ? 14'h213 : _GEN_16282;
  wire [13:0] _GEN_16284 = 14'h3f9c == index ? 14'h20f : _GEN_16283;
  wire [13:0] _GEN_16285 = 14'h3f9d == index ? 14'h20b : _GEN_16284;
  wire [13:0] _GEN_16286 = 14'h3f9e == index ? 14'h207 : _GEN_16285;
  wire [13:0] _GEN_16287 = 14'h3f9f == index ? 14'h203 : _GEN_16286;
  wire [13:0] _GEN_16288 = 14'h3fa0 == index ? 14'h19f : _GEN_16287;
  wire [13:0] _GEN_16289 = 14'h3fa1 == index ? 14'h19c : _GEN_16288;
  wire [13:0] _GEN_16290 = 14'h3fa2 == index ? 14'h199 : _GEN_16289;
  wire [13:0] _GEN_16291 = 14'h3fa3 == index ? 14'h196 : _GEN_16290;
  wire [13:0] _GEN_16292 = 14'h3fa4 == index ? 14'h193 : _GEN_16291;
  wire [13:0] _GEN_16293 = 14'h3fa5 == index ? 14'h190 : _GEN_16292;
  wire [13:0] _GEN_16294 = 14'h3fa6 == index ? 14'h18d : _GEN_16293;
  wire [13:0] _GEN_16295 = 14'h3fa7 == index ? 14'h18a : _GEN_16294;
  wire [13:0] _GEN_16296 = 14'h3fa8 == index ? 14'h187 : _GEN_16295;
  wire [13:0] _GEN_16297 = 14'h3fa9 == index ? 14'h184 : _GEN_16296;
  wire [13:0] _GEN_16298 = 14'h3faa == index ? 14'h181 : _GEN_16297;
  wire [13:0] _GEN_16299 = 14'h3fab == index ? 14'h129 : _GEN_16298;
  wire [13:0] _GEN_16300 = 14'h3fac == index ? 14'h127 : _GEN_16299;
  wire [13:0] _GEN_16301 = 14'h3fad == index ? 14'h125 : _GEN_16300;
  wire [13:0] _GEN_16302 = 14'h3fae == index ? 14'h123 : _GEN_16301;
  wire [13:0] _GEN_16303 = 14'h3faf == index ? 14'h121 : _GEN_16302;
  wire [13:0] _GEN_16304 = 14'h3fb0 == index ? 14'h11f : _GEN_16303;
  wire [13:0] _GEN_16305 = 14'h3fb1 == index ? 14'h11d : _GEN_16304;
  wire [13:0] _GEN_16306 = 14'h3fb2 == index ? 14'h11b : _GEN_16305;
  wire [13:0] _GEN_16307 = 14'h3fb3 == index ? 14'h119 : _GEN_16306;
  wire [13:0] _GEN_16308 = 14'h3fb4 == index ? 14'h117 : _GEN_16307;
  wire [13:0] _GEN_16309 = 14'h3fb5 == index ? 14'h115 : _GEN_16308;
  wire [13:0] _GEN_16310 = 14'h3fb6 == index ? 14'h113 : _GEN_16309;
  wire [13:0] _GEN_16311 = 14'h3fb7 == index ? 14'h111 : _GEN_16310;
  wire [13:0] _GEN_16312 = 14'h3fb8 == index ? 14'h10f : _GEN_16311;
  wire [13:0] _GEN_16313 = 14'h3fb9 == index ? 14'h10d : _GEN_16312;
  wire [13:0] _GEN_16314 = 14'h3fba == index ? 14'h10b : _GEN_16313;
  wire [13:0] _GEN_16315 = 14'h3fbb == index ? 14'h109 : _GEN_16314;
  wire [13:0] _GEN_16316 = 14'h3fbc == index ? 14'h107 : _GEN_16315;
  wire [13:0] _GEN_16317 = 14'h3fbd == index ? 14'h105 : _GEN_16316;
  wire [13:0] _GEN_16318 = 14'h3fbe == index ? 14'h103 : _GEN_16317;
  wire [13:0] _GEN_16319 = 14'h3fbf == index ? 14'h101 : _GEN_16318;
  wire [13:0] _GEN_16320 = 14'h3fc0 == index ? 14'hbf : _GEN_16319;
  wire [13:0] _GEN_16321 = 14'h3fc1 == index ? 14'hbe : _GEN_16320;
  wire [13:0] _GEN_16322 = 14'h3fc2 == index ? 14'hbd : _GEN_16321;
  wire [13:0] _GEN_16323 = 14'h3fc3 == index ? 14'hbc : _GEN_16322;
  wire [13:0] _GEN_16324 = 14'h3fc4 == index ? 14'hbb : _GEN_16323;
  wire [13:0] _GEN_16325 = 14'h3fc5 == index ? 14'hba : _GEN_16324;
  wire [13:0] _GEN_16326 = 14'h3fc6 == index ? 14'hb9 : _GEN_16325;
  wire [13:0] _GEN_16327 = 14'h3fc7 == index ? 14'hb8 : _GEN_16326;
  wire [13:0] _GEN_16328 = 14'h3fc8 == index ? 14'hb7 : _GEN_16327;
  wire [13:0] _GEN_16329 = 14'h3fc9 == index ? 14'hb6 : _GEN_16328;
  wire [13:0] _GEN_16330 = 14'h3fca == index ? 14'hb5 : _GEN_16329;
  wire [13:0] _GEN_16331 = 14'h3fcb == index ? 14'hb4 : _GEN_16330;
  wire [13:0] _GEN_16332 = 14'h3fcc == index ? 14'hb3 : _GEN_16331;
  wire [13:0] _GEN_16333 = 14'h3fcd == index ? 14'hb2 : _GEN_16332;
  wire [13:0] _GEN_16334 = 14'h3fce == index ? 14'hb1 : _GEN_16333;
  wire [13:0] _GEN_16335 = 14'h3fcf == index ? 14'hb0 : _GEN_16334;
  wire [13:0] _GEN_16336 = 14'h3fd0 == index ? 14'haf : _GEN_16335;
  wire [13:0] _GEN_16337 = 14'h3fd1 == index ? 14'hae : _GEN_16336;
  wire [13:0] _GEN_16338 = 14'h3fd2 == index ? 14'had : _GEN_16337;
  wire [13:0] _GEN_16339 = 14'h3fd3 == index ? 14'hac : _GEN_16338;
  wire [13:0] _GEN_16340 = 14'h3fd4 == index ? 14'hab : _GEN_16339;
  wire [13:0] _GEN_16341 = 14'h3fd5 == index ? 14'haa : _GEN_16340;
  wire [13:0] _GEN_16342 = 14'h3fd6 == index ? 14'ha9 : _GEN_16341;
  wire [13:0] _GEN_16343 = 14'h3fd7 == index ? 14'ha8 : _GEN_16342;
  wire [13:0] _GEN_16344 = 14'h3fd8 == index ? 14'ha7 : _GEN_16343;
  wire [13:0] _GEN_16345 = 14'h3fd9 == index ? 14'ha6 : _GEN_16344;
  wire [13:0] _GEN_16346 = 14'h3fda == index ? 14'ha5 : _GEN_16345;
  wire [13:0] _GEN_16347 = 14'h3fdb == index ? 14'ha4 : _GEN_16346;
  wire [13:0] _GEN_16348 = 14'h3fdc == index ? 14'ha3 : _GEN_16347;
  wire [13:0] _GEN_16349 = 14'h3fdd == index ? 14'ha2 : _GEN_16348;
  wire [13:0] _GEN_16350 = 14'h3fde == index ? 14'ha1 : _GEN_16349;
  wire [13:0] _GEN_16351 = 14'h3fdf == index ? 14'ha0 : _GEN_16350;
  wire [13:0] _GEN_16352 = 14'h3fe0 == index ? 14'h9f : _GEN_16351;
  wire [13:0] _GEN_16353 = 14'h3fe1 == index ? 14'h9e : _GEN_16352;
  wire [13:0] _GEN_16354 = 14'h3fe2 == index ? 14'h9d : _GEN_16353;
  wire [13:0] _GEN_16355 = 14'h3fe3 == index ? 14'h9c : _GEN_16354;
  wire [13:0] _GEN_16356 = 14'h3fe4 == index ? 14'h9b : _GEN_16355;
  wire [13:0] _GEN_16357 = 14'h3fe5 == index ? 14'h9a : _GEN_16356;
  wire [13:0] _GEN_16358 = 14'h3fe6 == index ? 14'h99 : _GEN_16357;
  wire [13:0] _GEN_16359 = 14'h3fe7 == index ? 14'h98 : _GEN_16358;
  wire [13:0] _GEN_16360 = 14'h3fe8 == index ? 14'h97 : _GEN_16359;
  wire [13:0] _GEN_16361 = 14'h3fe9 == index ? 14'h96 : _GEN_16360;
  wire [13:0] _GEN_16362 = 14'h3fea == index ? 14'h95 : _GEN_16361;
  wire [13:0] _GEN_16363 = 14'h3feb == index ? 14'h94 : _GEN_16362;
  wire [13:0] _GEN_16364 = 14'h3fec == index ? 14'h93 : _GEN_16363;
  wire [13:0] _GEN_16365 = 14'h3fed == index ? 14'h92 : _GEN_16364;
  wire [13:0] _GEN_16366 = 14'h3fee == index ? 14'h91 : _GEN_16365;
  wire [13:0] _GEN_16367 = 14'h3fef == index ? 14'h90 : _GEN_16366;
  wire [13:0] _GEN_16368 = 14'h3ff0 == index ? 14'h8f : _GEN_16367;
  wire [13:0] _GEN_16369 = 14'h3ff1 == index ? 14'h8e : _GEN_16368;
  wire [13:0] _GEN_16370 = 14'h3ff2 == index ? 14'h8d : _GEN_16369;
  wire [13:0] _GEN_16371 = 14'h3ff3 == index ? 14'h8c : _GEN_16370;
  wire [13:0] _GEN_16372 = 14'h3ff4 == index ? 14'h8b : _GEN_16371;
  wire [13:0] _GEN_16373 = 14'h3ff5 == index ? 14'h8a : _GEN_16372;
  wire [13:0] _GEN_16374 = 14'h3ff6 == index ? 14'h89 : _GEN_16373;
  wire [13:0] _GEN_16375 = 14'h3ff7 == index ? 14'h88 : _GEN_16374;
  wire [13:0] _GEN_16376 = 14'h3ff8 == index ? 14'h87 : _GEN_16375;
  wire [13:0] _GEN_16377 = 14'h3ff9 == index ? 14'h86 : _GEN_16376;
  wire [13:0] _GEN_16378 = 14'h3ffa == index ? 14'h85 : _GEN_16377;
  wire [13:0] _GEN_16379 = 14'h3ffb == index ? 14'h84 : _GEN_16378;
  wire [13:0] _GEN_16380 = 14'h3ffc == index ? 14'h83 : _GEN_16379;
  wire [13:0] _GEN_16381 = 14'h3ffd == index ? 14'h82 : _GEN_16380;
  wire [13:0] _GEN_16382 = 14'h3ffe == index ? 14'h81 : _GEN_16381;
  wire [13:0] _GEN_16383 = 14'h3fff == index ? 14'h80 : _GEN_16382;
  wire [63:0] divRes3 = io_in_isPow ? fastDivShift_io_out_s : {{57'd0}, _GEN_16383[13:7]};
  wire [63:0] _divRes2_T_1 = 64'h0 == io_in_op2_data ? 64'h0 : divRes3;
  wire [63:0] divRes2 = 64'h1 == io_in_op2_data ? io_in_op1_data : _divRes2_T_1;
  wire  _divRes_T = io_in_op1_data == io_in_op2_data;
  wire  _divRes_T_1 = io_in_op1_data < io_in_op2_data;
  wire [63:0] _divRes_T_3 = 64'h0 == io_in_op1_data ? 64'h0 : divRes2;
  wire [63:0] _divRes_T_4 = io_in_op1_data < io_in_op2_data ? 64'h0 : _divRes_T_3;
  wire [63:0] divRes = io_in_op1_data == io_in_op2_data ? 64'h1 : _divRes_T_4;
  wire [63:0] remRes3 = io_in_isPow ? fastDivShift_io_out_r : {{57'd0}, _GEN_16383[6:0]};
  wire [63:0] _remRes2_T_1 = 64'h0 == io_in_op2_data ? 64'h0 : remRes3;
  wire [63:0] remRes2 = 64'h1 == io_in_op2_data ? 64'h0 : _remRes2_T_1;
  wire [63:0] _remRes_T_3 = 64'h0 == io_in_op1_data ? 64'h0 : remRes2;
  wire [63:0] _remRes_T_4 = _divRes_T_1 ? io_in_op1_data : _remRes_T_3;
  wire [63:0] remRes = _divRes_T ? 64'h0 : _remRes_T_4;
  ysyx_040656_FastDivShift fastDivShift (
    .io_in_op1_data(fastDivShift_io_in_op1_data),
    .io_in_op2_data(fastDivShift_io_in_op2_data),
    .io_out_r(fastDivShift_io_out_r),
    .io_out_s(fastDivShift_io_out_s)
  );
  assign io_out_r = io_in_valid ? remRes : 64'h0;
  assign io_out_s = io_in_valid ? divRes : 64'h0;
  assign io_out_valid = io_in_valid;
  assign fastDivShift_io_in_op1_data = io_in_op1_data;
  assign fastDivShift_io_in_op2_data = io_in_op2_data;
endmodule
module ysyx_040656_DivCache(
  input         clock,
  input         reset,
  input  [63:0] io_in_op1_data,
  input  [63:0] io_in_op2_data,
  input  [63:0] io_in_s,
  input  [63:0] io_in_r,
  input         io_in_wen,
  input         io_in_valid,
  input         io_in_sign,
  input         io_in_isDiv,
  output        io_in_ready,
  output [63:0] io_out_s,
  output [63:0] io_out_r,
  output        io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif
  reg [129:0] key_0;
  reg [129:0] key_1;
  reg [129:0] key_2;
  reg [129:0] key_3;
  reg [129:0] key_4;
  reg [129:0] key_5;
  reg [63:0] value_0;
  reg [63:0] value_1;
  reg [63:0] value_2;
  reg [63:0] value_3;
  reg [63:0] value_4;
  reg [63:0] value_5;
  reg [2:0] cur;
  reg [63:0] hitValue;
  wire [129:0] _hit_0_T_2 = {io_in_op1_data,io_in_op2_data,io_in_sign,io_in_isDiv};
  wire  hit_0 = key_0 == _hit_0_T_2;
  wire [63:0] _GEN_0 = hit_0 ? value_0 : hitValue;
  wire  hit_1 = key_1 == _hit_0_T_2;
  wire [63:0] _GEN_1 = hit_1 ? value_1 : _GEN_0;
  wire  hit_2 = key_2 == _hit_0_T_2;
  wire [63:0] _GEN_2 = hit_2 ? value_2 : _GEN_1;
  wire  hit_3 = key_3 == _hit_0_T_2;
  wire  hit_4 = key_4 == _hit_0_T_2;
  wire  hit_5 = key_5 == _hit_0_T_2;
  wire [2:0] _cur_T_1 = cur + 3'h1;
  wire [5:0] _io_out_valid_T = {hit_5,hit_4,hit_3,hit_2,hit_1,hit_0};
  reg  io_out_valid_REG;
  reg  io_in_ready_REG;
  assign io_in_ready = ~io_in_valid | io_in_ready_REG;
  assign io_out_s = io_out_valid & io_in_isDiv ? hitValue : 64'h0;
  assign io_out_r = io_out_valid & ~io_in_isDiv ? hitValue : 64'h0;
  assign io_out_valid = io_out_valid_REG;
  always @(posedge clock) begin
    if (reset) begin
      key_0 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h0 == cur) begin
        key_0 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      key_1 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h1 == cur) begin
        key_1 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      key_2 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h2 == cur) begin
        key_2 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      key_3 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h3 == cur) begin
        key_3 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      key_4 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h4 == cur) begin
        key_4 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      key_5 <= 130'h0;
    end else if (io_in_wen) begin
      if (3'h5 == cur) begin
        key_5 <= _hit_0_T_2;
      end
    end
    if (reset) begin
      value_0 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h0 == cur) begin
        if (io_in_isDiv) begin
          value_0 <= io_in_s;
        end else begin
          value_0 <= io_in_r;
        end
      end
    end
    if (reset) begin
      value_1 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h1 == cur) begin
        if (io_in_isDiv) begin
          value_1 <= io_in_s;
        end else begin
          value_1 <= io_in_r;
        end
      end
    end
    if (reset) begin
      value_2 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h2 == cur) begin
        if (io_in_isDiv) begin
          value_2 <= io_in_s;
        end else begin
          value_2 <= io_in_r;
        end
      end
    end
    if (reset) begin
      value_3 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h3 == cur) begin
        if (io_in_isDiv) begin
          value_3 <= io_in_s;
        end else begin
          value_3 <= io_in_r;
        end
      end
    end
    if (reset) begin
      value_4 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h4 == cur) begin
        if (io_in_isDiv) begin
          value_4 <= io_in_s;
        end else begin
          value_4 <= io_in_r;
        end
      end
    end
    if (reset) begin
      value_5 <= 64'h0;
    end else if (io_in_wen) begin
      if (3'h5 == cur) begin
        if (io_in_isDiv) begin
          value_5 <= io_in_s;
        end else begin
          value_5 <= io_in_r;
        end
      end
    end
    if (reset) begin
      cur <= 3'h0;
    end else if (io_in_wen) begin
      if (cur < 3'h5) begin
        cur <= _cur_T_1;
      end else begin
        cur <= 3'h0;
      end
    end
    if (reset) begin
      hitValue <= 64'h0;
    end else if (hit_5) begin
      hitValue <= value_5;
    end else if (hit_4) begin
      hitValue <= value_4;
    end else if (hit_3) begin
      hitValue <= value_3;
    end else begin
      hitValue <= _GEN_2;
    end
    io_out_valid_REG <= |_io_out_valid_T & io_in_valid;
    io_in_ready_REG <= io_in_valid;
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  key_0 = _RAND_0[129:0];
  _RAND_1 = {5{`RANDOM}};
  key_1 = _RAND_1[129:0];
  _RAND_2 = {5{`RANDOM}};
  key_2 = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  key_3 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  key_4 = _RAND_4[129:0];
  _RAND_5 = {5{`RANDOM}};
  key_5 = _RAND_5[129:0];
  _RAND_6 = {2{`RANDOM}};
  value_0 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  value_1 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  value_2 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  value_3 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  value_4 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  value_5 = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  cur = _RAND_12[2:0];
  _RAND_13 = {2{`RANDOM}};
  hitValue = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  io_in_ready_REG = _RAND_15[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Mdu(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_op1_data,
  input  [63:0] io_in_bits_op2_data,
  input  [5:0]  io_in_bits_func,
  output        io_out_valid,
  output [63:0] io_out_bits
);
  wire  mul_clock;
  wire  mul_reset;
  wire  mul_io_in_valid;
  wire [63:0] mul_io_in_bits_op1;
  wire [63:0] mul_io_in_bits_op2;
  wire [5:0] mul_io_in_bits_func;
  wire  mul_io_out_valid;
  wire [127:0] mul_io_out_bits_dataout;
  wire  div_clock;
  wire  div_reset;
  wire  div_io_in_valid;
  wire  div_io_in_bits_sign;
  wire [63:0] div_io_in_bits_x;
  wire [63:0] div_io_in_bits_y;
  wire [5:0] div_io_in_bits_func;
  wire  div_io_out_valid;
  wire [63:0] div_io_out_bits_s;
  wire [63:0] div_io_out_bits_r;
  wire [63:0] fastDiv_io_in_op1_data;
  wire [63:0] fastDiv_io_in_op2_data;
  wire  fastDiv_io_in_valid;
  wire  fastDiv_io_in_isPow;
  wire [63:0] fastDiv_io_out_r;
  wire [63:0] fastDiv_io_out_s;
  wire  fastDiv_io_out_valid;
  wire  divCache_clock;
  wire  divCache_reset;
  wire [63:0] divCache_io_in_op1_data;
  wire [63:0] divCache_io_in_op2_data;
  wire [63:0] divCache_io_in_s;
  wire [63:0] divCache_io_in_r;
  wire  divCache_io_in_wen;
  wire  divCache_io_in_valid;
  wire  divCache_io_in_sign;
  wire  divCache_io_in_isDiv;
  wire  divCache_io_in_ready;
  wire [63:0] divCache_io_out_s;
  wire [63:0] divCache_io_out_r;
  wire  divCache_io_out_valid;
  wire  isDiv = 6'h27 == io_in_bits_func | (6'h26 == io_in_bits_func | (6'h22 == io_in_bits_func | 6'h21 ==
    io_in_bits_func));
  wire  isRem = 6'h24 == io_in_bits_func | (6'h23 == io_in_bits_func | (6'h29 == io_in_bits_func | 6'h28 ==
    io_in_bits_func));
  wire  isMul = 6'h1f == io_in_bits_func | (6'h20 == io_in_bits_func | (6'h1e == io_in_bits_func | (6'h25 ==
    io_in_bits_func | 6'h1d == io_in_bits_func)));
  wire  isW = 6'h29 == io_in_bits_func | (6'h28 == io_in_bits_func | (6'h27 == io_in_bits_func | (6'h27 ==
    io_in_bits_func | (6'h26 == io_in_bits_func | 6'h25 == io_in_bits_func))));
  wire  isMulH = 6'h1e == io_in_bits_func | (6'h20 == io_in_bits_func | 6'h1f == io_in_bits_func);
  wire  isSign = 6'h28 == io_in_bits_func | (6'h23 == io_in_bits_func | (6'h26 == io_in_bits_func | 6'h21 ==
    io_in_bits_func));
  wire [63:0] _isPow_T_1 = io_in_bits_op2_data - 64'h1;
  wire [63:0] _isPow_T_2 = io_in_bits_op2_data & _isPow_T_1;
  wire  _isPow_T_4 = io_in_bits_op2_data != 64'h0;
  wire  isPow = _isPow_T_2 == 64'h0 & io_in_bits_op2_data != 64'h0;
  wire  _isFast_T = isDiv | isRem;
  wire  _isFast_T_3 = io_in_bits_op1_data < 64'h80;
  wire  _isFast_T_6 = io_in_bits_op2_data < 64'h80;
  wire  _isFast_T_7 = _isFast_T_3 & _isFast_T_6;
  wire  _isFast_T_8 = io_in_bits_op2_data > 64'h0;
  wire  _isFast_T_9 = _isFast_T_7 & _isFast_T_8;
  wire  _isFast_T_13 = ~isSign & (io_in_bits_op1_data <= io_in_bits_op2_data | isPow);
  wire  _isFast_T_14 = _isFast_T_9 | _isFast_T_13;
  wire  isFast = (isDiv | isRem) & _isPow_T_4 & _isFast_T_14;
  wire [63:0] mulRes = isMulH ? mul_io_out_bits_dataout[127:64] : mul_io_out_bits_dataout[63:0];
  wire [31:0] _div_io_in_bits_x_T_6 = io_in_bits_op1_data[31] ? 32'hffffffff : 32'h0;
  wire [63:0] _div_io_in_bits_x_T_8 = {_div_io_in_bits_x_T_6,io_in_bits_op1_data[31:0]};
  wire [63:0] _div_io_in_bits_x_T_12 = {32'h0,io_in_bits_op1_data[31:0]};
  wire [63:0] _div_io_in_bits_x_T_14 = 6'h21 == io_in_bits_func ? io_in_bits_op1_data : 64'h0;
  wire [63:0] _div_io_in_bits_x_T_16 = 6'h22 == io_in_bits_func ? io_in_bits_op1_data : _div_io_in_bits_x_T_14;
  wire [63:0] _div_io_in_bits_x_T_18 = 6'h26 == io_in_bits_func ? _div_io_in_bits_x_T_8 : _div_io_in_bits_x_T_16;
  wire [63:0] _div_io_in_bits_x_T_20 = 6'h27 == io_in_bits_func ? _div_io_in_bits_x_T_12 : _div_io_in_bits_x_T_18;
  wire [31:0] _div_io_in_bits_y_T_6 = io_in_bits_op2_data[31] ? 32'hffffffff : 32'h0;
  wire [63:0] _div_io_in_bits_y_T_8 = {_div_io_in_bits_y_T_6,io_in_bits_op2_data[31:0]};
  wire [63:0] _div_io_in_bits_y_T_12 = {32'h0,io_in_bits_op2_data[31:0]};
  wire [63:0] _div_io_in_bits_y_T_14 = 6'h21 == io_in_bits_func ? io_in_bits_op2_data : 64'h0;
  wire [63:0] _div_io_in_bits_y_T_16 = 6'h22 == io_in_bits_func ? io_in_bits_op2_data : _div_io_in_bits_y_T_14;
  wire [63:0] _div_io_in_bits_y_T_18 = 6'h26 == io_in_bits_func ? _div_io_in_bits_y_T_8 : _div_io_in_bits_y_T_16;
  wire [63:0] _div_io_in_bits_y_T_20 = 6'h27 == io_in_bits_func ? _div_io_in_bits_y_T_12 : _div_io_in_bits_y_T_18;
  wire [63:0] _div_io_in_bits_x_T_35 = 6'h23 == io_in_bits_func ? io_in_bits_op1_data : 64'h0;
  wire [63:0] _div_io_in_bits_x_T_37 = 6'h24 == io_in_bits_func ? io_in_bits_op1_data : _div_io_in_bits_x_T_35;
  wire [63:0] _div_io_in_bits_x_T_39 = 6'h28 == io_in_bits_func ? _div_io_in_bits_x_T_8 : _div_io_in_bits_x_T_37;
  wire [63:0] _div_io_in_bits_x_T_41 = 6'h29 == io_in_bits_func ? _div_io_in_bits_x_T_12 : _div_io_in_bits_x_T_39;
  wire [63:0] _div_io_in_bits_y_T_35 = 6'h23 == io_in_bits_func ? io_in_bits_op2_data : 64'h0;
  wire [63:0] _div_io_in_bits_y_T_37 = 6'h24 == io_in_bits_func ? io_in_bits_op2_data : _div_io_in_bits_y_T_35;
  wire [63:0] _div_io_in_bits_y_T_39 = 6'h28 == io_in_bits_func ? _div_io_in_bits_y_T_8 : _div_io_in_bits_y_T_37;
  wire [63:0] _div_io_in_bits_y_T_41 = 6'h29 == io_in_bits_func ? _div_io_in_bits_y_T_12 : _div_io_in_bits_y_T_39;
  wire [63:0] _GEN_0 = isRem ? _div_io_in_bits_x_T_41 : 64'h0;
  wire [63:0] _GEN_1 = isRem ? _div_io_in_bits_y_T_41 : 64'h1;
  wire  _GEN_2 = isRem & isSign;
  wire  _divValid_T_2 = ~isFast;
  wire  divValid = io_in_valid & _isFast_T & ~isFast;
  wire [63:0] _divRes_T = divCache_io_out_valid ? divCache_io_out_s : div_io_out_bits_s;
  wire [63:0] divRes = isFast ? fastDiv_io_out_s : _divRes_T;
  wire [63:0] _RemRes_T = divCache_io_out_valid ? divCache_io_out_r : div_io_out_bits_r;
  wire [63:0] RemRes = isFast ? fastDiv_io_out_r : _RemRes_T;
  wire [63:0] _res_T = isMul ? mulRes : 64'h0;
  wire [63:0] _res_T_1 = isDiv ? divRes : _res_T;
  wire [63:0] res = isRem ? RemRes : _res_T_1;
  wire  _io_out_valid_T_2 = _isFast_T & _divValid_T_2;
  wire  _io_out_valid_T_3 = div_io_out_valid | divCache_io_out_valid;
  wire  _io_out_valid_T_5 = _io_out_valid_T_2 ? _io_out_valid_T_3 : isMul & mul_io_out_valid;
  wire  _io_out_valid_T_6 = isFast ? fastDiv_io_out_valid : _io_out_valid_T_5;
  wire  io_out_bits_signBit = res[31];
  wire [31:0] _io_out_bits_T_2 = io_out_bits_signBit ? 32'hffffffff : 32'h0;
  wire [63:0] _io_out_bits_T_3 = {_io_out_bits_T_2,res[31:0]};
  ysyx_040656_ExternalMul mul (
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_op1(mul_io_in_bits_op1),
    .io_in_bits_op2(mul_io_in_bits_op2),
    .io_in_bits_func(mul_io_in_bits_func),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits_dataout(mul_io_out_bits_dataout)
  );
  ysyx_040656_ExternalDiv div (
    .clock(div_clock),
    .reset(div_reset),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_sign(div_io_in_bits_sign),
    .io_in_bits_x(div_io_in_bits_x),
    .io_in_bits_y(div_io_in_bits_y),
    .io_in_bits_func(div_io_in_bits_func),
    .io_out_valid(div_io_out_valid),
    .io_out_bits_s(div_io_out_bits_s),
    .io_out_bits_r(div_io_out_bits_r)
  );
  ysyx_040656_FastDiv fastDiv (
    .io_in_op1_data(fastDiv_io_in_op1_data),
    .io_in_op2_data(fastDiv_io_in_op2_data),
    .io_in_valid(fastDiv_io_in_valid),
    .io_in_isPow(fastDiv_io_in_isPow),
    .io_out_r(fastDiv_io_out_r),
    .io_out_s(fastDiv_io_out_s),
    .io_out_valid(fastDiv_io_out_valid)
  );
  ysyx_040656_DivCache divCache (
    .clock(divCache_clock),
    .reset(divCache_reset),
    .io_in_op1_data(divCache_io_in_op1_data),
    .io_in_op2_data(divCache_io_in_op2_data),
    .io_in_s(divCache_io_in_s),
    .io_in_r(divCache_io_in_r),
    .io_in_wen(divCache_io_in_wen),
    .io_in_valid(divCache_io_in_valid),
    .io_in_sign(divCache_io_in_sign),
    .io_in_isDiv(divCache_io_in_isDiv),
    .io_in_ready(divCache_io_in_ready),
    .io_out_s(divCache_io_out_s),
    .io_out_r(divCache_io_out_r),
    .io_out_valid(divCache_io_out_valid)
  );
  assign io_out_valid = io_in_valid & _io_out_valid_T_6;
  assign io_out_bits = isW ? _io_out_bits_T_3 : res;
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & isMul;
  assign mul_io_in_bits_op1 = isMul ? io_in_bits_op1_data : 64'h0;
  assign mul_io_in_bits_op2 = isMul ? io_in_bits_op2_data : 64'h0;
  assign mul_io_in_bits_func = io_in_bits_func;
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = ~divCache_io_out_valid & divCache_io_in_ready & divValid;
  assign div_io_in_bits_sign = isDiv ? isSign : _GEN_2;
  assign div_io_in_bits_x = isDiv ? _div_io_in_bits_x_T_20 : _GEN_0;
  assign div_io_in_bits_y = isDiv ? _div_io_in_bits_y_T_20 : _GEN_1;
  assign div_io_in_bits_func = io_in_bits_func;
  assign fastDiv_io_in_op1_data = div_io_in_bits_x;
  assign fastDiv_io_in_op2_data = div_io_in_bits_y;
  assign fastDiv_io_in_valid = io_in_valid & isFast;
  assign fastDiv_io_in_isPow = _isPow_T_2 == 64'h0 & io_in_bits_op2_data != 64'h0;
  assign divCache_clock = clock;
  assign divCache_reset = reset;
  assign divCache_io_in_op1_data = div_io_in_bits_x;
  assign divCache_io_in_op2_data = div_io_in_bits_y;
  assign divCache_io_in_s = div_io_out_bits_s;
  assign divCache_io_in_r = div_io_out_bits_r;
  assign divCache_io_in_wen = div_io_out_valid;
  assign divCache_io_in_valid = io_in_valid & _isFast_T & ~isFast;
  assign divCache_io_in_sign = div_io_in_bits_sign;
  assign divCache_io_in_isDiv = 6'h27 == io_in_bits_func | (6'h26 == io_in_bits_func | (6'h22 == io_in_bits_func | 6'h21
     == io_in_bits_func));
endmodule
module ysyx_040656_Lsu(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [5:0]  io_in_bits_func,
  input  [63:0] io_in_bits_rs2_data,
  output        io_out_valid,
  output [63:0] io_out_bits_data,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [1:0]  io_dmem_req_bits_size,
  output [2:0]  io_dmem_req_bits_cmd,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [63:0] io_mmio_req_bits_wdata,
  output [1:0]  io_mmio_req_bits_size,
  output [2:0]  io_mmio_req_bits_cmd,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif
  wire [5:0] shift = {io_in_bits_addr[2:0], 3'h0};
  wire  addrAtMMIO_selVec_0 = io_in_bits_addr <= 32'h1ffffff;
  wire  addrAtMMIO_selVec_1 = io_in_bits_addr >= 32'h2000000 & io_in_bits_addr <= 32'h200ffff;
  wire  addrAtMMIO_selVec_2 = io_in_bits_addr >= 32'h2010000 & io_in_bits_addr <= 32'h7fffffff;
  wire  addrAtMMIO_selVec_3 = io_in_bits_addr >= 32'hfc000000;
  wire [3:0] _addrAtMMIO_hit_T = {addrAtMMIO_selVec_3,addrAtMMIO_selVec_2,addrAtMMIO_selVec_1,addrAtMMIO_selVec_0};
  wire  addrAtMMIO_hit = |_addrAtMMIO_hit_T;
  wire  addrAtMMIO = addrAtMMIO_hit & io_in_valid;
  reg [1:0] lsuStatus;
  wire [1:0] _size_T_17 = 6'h14 == io_in_bits_func ? 2'h2 : {{1'd0}, 6'h13 == io_in_bits_func};
  wire [1:0] _size_T_19 = 6'h15 == io_in_bits_func ? 2'h3 : _size_T_17;
  wire [1:0] _size_T_21 = 6'h16 == io_in_bits_func ? 2'h0 : _size_T_19;
  wire [1:0] _size_T_23 = 6'h17 == io_in_bits_func ? 2'h1 : _size_T_21;
  wire [1:0] _size_T_25 = 6'h18 == io_in_bits_func ? 2'h2 : _size_T_23;
  wire [1:0] _size_T_27 = 6'h19 == io_in_bits_func ? 2'h0 : _size_T_25;
  wire [1:0] _size_T_29 = 6'h1a == io_in_bits_func ? 2'h1 : _size_T_27;
  wire [1:0] _size_T_31 = 6'h1b == io_in_bits_func ? 2'h2 : _size_T_29;
  wire [1:0] size = 6'h1c == io_in_bits_func ? 2'h3 : _size_T_31;
  wire [63:0] _wdata_T_2 = {56'h0,io_in_bits_rs2_data[7:0]};
  wire [63:0] _wdata_T_5 = {48'h0,io_in_bits_rs2_data[15:0]};
  wire [63:0] _wdata_T_8 = {32'h0,io_in_bits_rs2_data[31:0]};
  wire [63:0] _wdata_T_10 = 2'h1 == size ? _wdata_T_5 : _wdata_T_2;
  wire [63:0] _wdata_T_12 = 2'h2 == size ? _wdata_T_8 : _wdata_T_10;
  wire [63:0] wdata = 2'h3 == size ? io_in_bits_rs2_data : _wdata_T_12;
  wire  isStore = 6'h1c == io_in_bits_func | (6'h1b == io_in_bits_func | (6'h1a == io_in_bits_func | 6'h19 ==
    io_in_bits_func));
  wire  _T_26 = io_mmio_resp_ready & io_mmio_resp_valid;
  wire  _T_28 = ~addrAtMMIO;
  wire  _T_29 = io_dmem_resp_ready & io_dmem_resp_valid;
  wire  _T_31 = addrAtMMIO & _T_26 | ~addrAtMMIO & _T_29;
  wire [63:0] _readBuffer_T = io_mmio_resp_bits_rdata >> shift;
  wire [63:0] _readBuffer_T_1 = addrAtMMIO ? _readBuffer_T : io_dmem_resp_bits_rdata;
  wire [63:0] _readBuffer_T_2 = isStore ? 64'hdeadc0de : _readBuffer_T_1;
  wire [63:0] _GEN_4 = addrAtMMIO & _T_26 | ~addrAtMMIO & _T_29 ? _readBuffer_T_2 : 64'h0;
  wire [63:0] _GEN_7 = 2'h2 == lsuStatus ? _GEN_4 : 64'h0;
  wire [63:0] _GEN_10 = 2'h1 == lsuStatus ? 64'h0 : _GEN_7;
  wire [63:0] readBuffer = 2'h0 == lsuStatus ? 64'h0 : _GEN_10;
  wire [55:0] _data_T_4 = readBuffer[7] ? 56'hffffffffffffff : 56'h0;
  wire [63:0] _data_T_6 = {_data_T_4,readBuffer[7:0]};
  wire [47:0] _data_T_10 = readBuffer[15] ? 48'hffffffffffff : 48'h0;
  wire [63:0] _data_T_12 = {_data_T_10,readBuffer[15:0]};
  wire [31:0] _data_T_16 = readBuffer[31] ? 32'hffffffff : 32'h0;
  wire [63:0] _data_T_18 = {_data_T_16,readBuffer[31:0]};
  wire [63:0] _data_T_23 = {56'h0,readBuffer[7:0]};
  wire [63:0] _data_T_27 = {48'h0,readBuffer[15:0]};
  wire [63:0] _data_T_31 = {32'h0,readBuffer[31:0]};
  wire [63:0] _data_T_33 = 6'h12 == io_in_bits_func ? _data_T_6 : readBuffer;
  wire [63:0] _data_T_35 = 6'h13 == io_in_bits_func ? _data_T_12 : _data_T_33;
  wire [63:0] _data_T_37 = 6'h14 == io_in_bits_func ? _data_T_18 : _data_T_35;
  wire [63:0] _data_T_39 = 6'h15 == io_in_bits_func ? readBuffer : _data_T_37;
  wire [63:0] _data_T_41 = 6'h16 == io_in_bits_func ? _data_T_23 : _data_T_39;
  wire [63:0] _data_T_43 = 6'h17 == io_in_bits_func ? _data_T_27 : _data_T_41;
  wire [63:0] _wdataOut_T_3 = {wdata[55:0],8'h0};
  wire [63:0] _wdataOut_T_6 = {wdata[47:0],16'h0};
  wire [63:0] _wdataOut_T_9 = {wdata[39:0],24'h0};
  wire [63:0] _wdataOut_T_12 = {wdata[31:0],32'h0};
  wire [63:0] _wdataOut_T_15 = {wdata[23:0],40'h0};
  wire [63:0] _wdataOut_T_18 = {wdata[15:0],48'h0};
  wire [63:0] _wdataOut_T_21 = {wdata[7:0],56'h0};
  wire [63:0] _wdataOut_T_23 = 3'h1 == io_in_bits_addr[2:0] ? _wdataOut_T_3 : wdata;
  wire [63:0] _wdataOut_T_25 = 3'h2 == io_in_bits_addr[2:0] ? _wdataOut_T_6 : _wdataOut_T_23;
  wire [63:0] _wdataOut_T_27 = 3'h3 == io_in_bits_addr[2:0] ? _wdataOut_T_9 : _wdataOut_T_25;
  wire [63:0] _wdataOut_T_29 = 3'h4 == io_in_bits_addr[2:0] ? _wdataOut_T_12 : _wdataOut_T_27;
  wire [63:0] _wdataOut_T_31 = 3'h5 == io_in_bits_addr[2:0] ? _wdataOut_T_15 : _wdataOut_T_29;
  wire [63:0] _wdataOut_T_33 = 3'h6 == io_in_bits_addr[2:0] ? _wdataOut_T_18 : _wdataOut_T_31;
  wire  _T_3 = lsuStatus == 2'h1 | lsuStatus == 2'h0 & io_in_valid;
  wire  _T_12 = io_mmio_req_ready & io_mmio_req_valid;
  wire  _T_15 = io_dmem_req_ready & io_dmem_req_valid;
  wire  _T_17 = addrAtMMIO & _T_12 | _T_28 & _T_15;
  wire [1:0] _GEN_3 = addrAtMMIO & _T_26 | ~addrAtMMIO & _T_29 ? 2'h0 : lsuStatus;
  wire  _GEN_11 = 2'h1 == lsuStatus ? 1'h0 : 2'h2 == lsuStatus & _T_31;
  assign io_out_valid = 2'h0 == lsuStatus ? 1'h0 : _GEN_11;
  assign io_out_bits_data = 6'h18 == io_in_bits_func ? _data_T_31 : _data_T_43;
  assign io_dmem_req_valid = (lsuStatus == 2'h1 | lsuStatus == 2'h0 & io_in_valid) & _T_28;
  assign io_dmem_req_bits_addr = io_in_bits_addr;
  assign io_dmem_req_bits_wdata = 3'h7 == io_in_bits_addr[2:0] ? _wdataOut_T_21 : _wdataOut_T_33;
  assign io_dmem_req_bits_size = 6'h1c == io_in_bits_func ? 2'h3 : _size_T_31;
  assign io_dmem_req_bits_cmd = {{2'd0}, isStore};
  assign io_dmem_resp_ready = 1'h1;
  assign io_mmio_req_valid = _T_3 & addrAtMMIO;
  assign io_mmio_req_bits_addr = io_in_bits_addr;
  assign io_mmio_req_bits_wdata = 3'h7 == io_in_bits_addr[2:0] ? _wdataOut_T_21 : _wdataOut_T_33;
  assign io_mmio_req_bits_size = 6'h1c == io_in_bits_func ? 2'h3 : _size_T_31;
  assign io_mmio_req_bits_cmd = {{2'd0}, isStore};
  assign io_mmio_resp_ready = 1'h1;
  always @(posedge clock) begin
    if (reset) begin
      lsuStatus <= 2'h0;
    end else if (2'h0 == lsuStatus) begin
      if (io_in_valid) begin
        if (addrAtMMIO & _T_12 | _T_28 & _T_15) begin
          lsuStatus <= 2'h2;
        end else begin
          lsuStatus <= 2'h1;
        end
      end
    end else if (2'h1 == lsuStatus) begin
      if (_T_17) begin
        lsuStatus <= 2'h2;
      end
    end else if (2'h2 == lsuStatus) begin
      lsuStatus <= _GEN_3;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lsuStatus = _RAND_0[1:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Csr(
  input         clock,
  input         reset,
  input         io_req_valid,
  input  [31:0] io_req_bits_pc,
  input  [5:0]  io_req_bits_cmd,
  input  [11:0] io_req_bits_addr,
  input  [63:0] io_req_bits_wdata,
  input  [4:0]  io_req_bits_rd,
  input         io_req_bits_valid,
  output [63:0] io_resp_bits_rdata,
  output        io_redirect_valid,
  output [31:0] io_redirect_target,
  output        io_en,
  output        io_raiseIntr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
`endif
  reg [1:0] mode;
  reg [63:0] reg_satp;
  reg [63:0] reg_sepc;
  reg [63:0] reg_sstatus;
  reg [63:0] reg_sedeleg;
  reg [63:0] reg_sideleg;
  reg [63:0] reg_sie;
  reg [63:0] reg_stvec;
  reg [63:0] reg_scounteren;
  reg [63:0] reg_sscratch;
  reg [63:0] reg_scause;
  reg [63:0] reg_stval;
  reg [63:0] reg_sip;
  reg [63:0] reg_mhartid;
  reg [63:0] reg_mstatus;
  reg [63:0] reg_misa;
  reg [63:0] reg_medeleg;
  reg [63:0] reg_mideleg;
  reg [63:0] reg_mie;
  reg [61:0] reg_mtvec_BASE;
  reg [1:0] reg_mtvec_MODE;
  reg [63:0] reg_mscratch;
  reg [63:0] reg_mepc;
  reg  reg_mcause_interrupt;
  reg [62:0] reg_mcause_exc_code;
  reg [63:0] reg_mtval;
  reg [51:0] reg_mip_reserved;
  reg  reg_mip_intr_e_m;
  reg  reg_mip_intr_e_h;
  reg  reg_mip_intr_e_s;
  reg  reg_mip_intr_e_u;
  reg  reg_mip_intr_t_m;
  reg  reg_mip_intr_t_h;
  reg  reg_mip_intr_t_s;
  reg  reg_mip_intr_t_u;
  reg  reg_mip_intr_s_m;
  reg  reg_mip_intr_s_h;
  reg  reg_mip_intr_s_s;
  reg  reg_mip_intr_s_u;
  reg  reg_mip_MEIP;
  reg  reg_mip_reserved_2;
  reg  reg_mip_SEIP;
  reg  reg_mip_UEIP;
  reg  reg_mip_MTIP;
  reg  reg_mip_reserved_3;
  reg  reg_mip_STIP;
  reg  reg_mip_UTIP;
  reg  reg_mip_MSIP;
  reg  reg_mip_reserved_4;
  reg  reg_mip_SSIP;
  reg  reg_mip_USIP;
  reg [63:0] reg_pmpcfg0;
  reg [63:0] reg_pmpcfg1;
  reg [63:0] reg_pmpcfg2;
  reg [63:0] reg_pmpcfg3;
  reg [63:0] reg_pmpaddr0;
  reg [63:0] mcycle;
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1;
  wire [5:0] mip2_lo_1 = {reg_mip_intr_t_s,reg_mip_intr_t_u,reg_mip_intr_s_m,reg_mip_intr_s_h,reg_mip_intr_s_s,
    reg_mip_intr_s_u};
  wire [11:0] _mip2_T_1 = {reg_mip_intr_e_m,reg_mip_intr_e_h,reg_mip_intr_e_s,reg_mip_intr_e_u,reg_mip_intr_t_m,
    reg_mip_intr_t_h,mip2_lo_1};
  wire  mip2_s_u = _mip2_T_1[0];
  wire  mip2_s_s = _mip2_T_1[1];
  wire  mip2_s_h = _mip2_T_1[2];
  wire  mip2_s_m = _mip2_T_1[3];
  wire  mip2_t_u = _mip2_T_1[4];
  wire  mip2_t_s = _mip2_T_1[5];
  wire  mip2_t_h = _mip2_T_1[6];
  wire  mip2_t_m = _mip2_T_1[7];
  wire  mip2_e_u = _mip2_T_1[8];
  wire  mip2_e_s = _mip2_T_1[9];
  wire  mip2_e_h = _mip2_T_1[10];
  wire  mip2_e_m = _mip2_T_1[11];
  wire  mstatusStruct_IE_u = reg_mstatus[0];
  wire  mstatusStruct_IE_s = reg_mstatus[1];
  wire  mstatusStruct_IE_h = reg_mstatus[2];
  wire  mstatusStruct_IE_m = reg_mstatus[3];
  wire  mstatusStruct_PIE_u = reg_mstatus[4];
  wire  mstatusStruct_PIE_s = reg_mstatus[5];
  wire  mstatusStruct_PIE_h = reg_mstatus[6];
  wire  mstatusStruct_PIE_m = reg_mstatus[7];
  wire  mstatusStruct_SPP = reg_mstatus[8];
  wire [1:0] mstatusStruct_reserved_2 = reg_mstatus[10:9];
  wire [1:0] mstatusStruct_MPP = reg_mstatus[12:11];
  wire [1:0] mstatusStruct_FS = reg_mstatus[14:13];
  wire [1:0] mstatusStruct_XS = reg_mstatus[16:15];
  wire  mstatusStruct_MPRV = reg_mstatus[17];
  wire  mstatusStruct_SUM = reg_mstatus[18];
  wire  mstatusStruct_MXR = reg_mstatus[19];
  wire  mstatusStruct_TVM = reg_mstatus[20];
  wire  mstatusStruct_TW = reg_mstatus[21];
  wire  mstatusStruct_TSR = reg_mstatus[22];
  wire [39:0] mstatusStruct_reserved = reg_mstatus[62:23];
  wire  mstatusStruct_SD = reg_mstatus[63];
  wire [63:0] _read_csr_data_T = {reg_mtvec_BASE,reg_mtvec_MODE};
  wire [63:0] _read_csr_data_T_1 = {reg_mcause_interrupt,reg_mcause_exc_code};
  wire [5:0] read_csr_data_lo_lo = {reg_mip_STIP,reg_mip_UTIP,reg_mip_MSIP,reg_mip_reserved_4,reg_mip_SSIP,reg_mip_USIP}
    ;
  wire [11:0] read_csr_data_lo = {reg_mip_MEIP,reg_mip_reserved_2,reg_mip_SEIP,reg_mip_UEIP,reg_mip_MTIP,
    reg_mip_reserved_3,read_csr_data_lo_lo};
  wire [75:0] _read_csr_data_T_2 = {reg_mip_reserved,reg_mip_intr_e_m,reg_mip_intr_e_h,reg_mip_intr_e_s,reg_mip_intr_e_u
    ,reg_mip_intr_t_m,reg_mip_intr_t_h,mip2_lo_1,read_csr_data_lo};
  wire [63:0] _read_csr_data_T_4 = 12'h180 == io_req_bits_addr ? reg_satp : 64'h0;
  wire [63:0] _read_csr_data_T_6 = 12'h141 == io_req_bits_addr ? reg_sepc : _read_csr_data_T_4;
  wire [63:0] _read_csr_data_T_8 = 12'h100 == io_req_bits_addr ? reg_sstatus : _read_csr_data_T_6;
  wire [63:0] _read_csr_data_T_10 = 12'h102 == io_req_bits_addr ? reg_sedeleg : _read_csr_data_T_8;
  wire [63:0] _read_csr_data_T_12 = 12'h103 == io_req_bits_addr ? reg_sideleg : _read_csr_data_T_10;
  wire [63:0] _read_csr_data_T_14 = 12'h104 == io_req_bits_addr ? reg_sie : _read_csr_data_T_12;
  wire [63:0] _read_csr_data_T_16 = 12'h105 == io_req_bits_addr ? reg_stvec : _read_csr_data_T_14;
  wire [63:0] _read_csr_data_T_18 = 12'h106 == io_req_bits_addr ? reg_scounteren : _read_csr_data_T_16;
  wire [63:0] _read_csr_data_T_20 = 12'h140 == io_req_bits_addr ? reg_sscratch : _read_csr_data_T_18;
  wire [63:0] _read_csr_data_T_22 = 12'h142 == io_req_bits_addr ? reg_scause : _read_csr_data_T_20;
  wire [63:0] _read_csr_data_T_24 = 12'h143 == io_req_bits_addr ? reg_stval : _read_csr_data_T_22;
  wire [63:0] _read_csr_data_T_26 = 12'h144 == io_req_bits_addr ? reg_sip : _read_csr_data_T_24;
  wire [102:0] _read_csr_data_T_28 = 12'hf12 == io_req_bits_addr ? 103'h7f7f7f7f7f7f7f7f7f7f7f7f8a : {{39'd0},
    _read_csr_data_T_26};
  wire [102:0] _read_csr_data_T_30 = 12'hf11 == io_req_bits_addr ? 103'h60a : _read_csr_data_T_28;
  wire [102:0] _read_csr_data_T_32 = 12'hf14 == io_req_bits_addr ? {{39'd0}, reg_mhartid} : _read_csr_data_T_30;
  wire [102:0] _read_csr_data_T_34 = 12'h300 == io_req_bits_addr ? {{39'd0}, reg_mstatus} : _read_csr_data_T_32;
  wire [102:0] _read_csr_data_T_36 = 12'h301 == io_req_bits_addr ? {{39'd0}, reg_misa} : _read_csr_data_T_34;
  wire [102:0] _read_csr_data_T_38 = 12'h302 == io_req_bits_addr ? {{39'd0}, reg_medeleg} : _read_csr_data_T_36;
  wire [102:0] _read_csr_data_T_40 = 12'h303 == io_req_bits_addr ? {{39'd0}, reg_mideleg} : _read_csr_data_T_38;
  wire [102:0] _read_csr_data_T_42 = 12'h304 == io_req_bits_addr ? {{39'd0}, reg_mie} : _read_csr_data_T_40;
  wire [102:0] _read_csr_data_T_44 = 12'h305 == io_req_bits_addr ? {{39'd0}, _read_csr_data_T} : _read_csr_data_T_42;
  wire [102:0] _read_csr_data_T_46 = 12'h340 == io_req_bits_addr ? {{39'd0}, reg_mscratch} : _read_csr_data_T_44;
  wire [102:0] _read_csr_data_T_48 = 12'h341 == io_req_bits_addr ? {{39'd0}, reg_mepc} : _read_csr_data_T_46;
  wire [102:0] _read_csr_data_T_50 = 12'h342 == io_req_bits_addr ? {{39'd0}, _read_csr_data_T_1} : _read_csr_data_T_48;
  wire [102:0] _read_csr_data_T_52 = 12'h343 == io_req_bits_addr ? {{39'd0}, reg_mtval} : _read_csr_data_T_50;
  wire [102:0] _read_csr_data_T_54 = 12'h344 == io_req_bits_addr ? {{27'd0}, _read_csr_data_T_2} : _read_csr_data_T_52;
  wire [102:0] _read_csr_data_T_56 = 12'h3a0 == io_req_bits_addr ? {{39'd0}, reg_pmpcfg0} : _read_csr_data_T_54;
  wire [102:0] _read_csr_data_T_58 = 12'h3a1 == io_req_bits_addr ? {{39'd0}, reg_pmpcfg1} : _read_csr_data_T_56;
  wire [102:0] _read_csr_data_T_60 = 12'h3a2 == io_req_bits_addr ? {{39'd0}, reg_pmpcfg2} : _read_csr_data_T_58;
  wire [102:0] _read_csr_data_T_62 = 12'h3a3 == io_req_bits_addr ? {{39'd0}, reg_pmpcfg3} : _read_csr_data_T_60;
  wire [102:0] _read_csr_data_T_64 = 12'h3b0 == io_req_bits_addr ? {{39'd0}, reg_pmpaddr0} : _read_csr_data_T_62;
  wire [102:0] _read_csr_data_T_66 = 12'hb00 == io_req_bits_addr ? {{39'd0}, mcycle} : _read_csr_data_T_64;
  wire [63:0] read_csr_data = _read_csr_data_T_66[63:0];
  wire [63:0] _write_data_T_3 = read_csr_data | io_req_bits_wdata;
  wire [63:0] _write_data_T_5 = ~io_req_bits_wdata;
  wire [63:0] _write_data_T_6 = read_csr_data & _write_data_T_5;
  wire [63:0] _write_data_T_8 = 6'h2e == io_req_bits_cmd ? io_req_bits_wdata : 64'h0;
  wire [63:0] _write_data_T_10 = 6'h2f == io_req_bits_cmd ? _write_data_T_3 : _write_data_T_8;
  wire [63:0] write_data = 6'h30 == io_req_bits_cmd ? _write_data_T_6 : _write_data_T_10;
  wire  system_ins = io_req_bits_cmd == 6'h31;
  wire  cpu_ren = io_req_bits_cmd != 6'h2d & ~system_ins;
  wire  wen = io_req_valid & cpu_ren & io_req_bits_cmd != 6'h32;
  wire [7:0] opcode = 8'h1 << io_req_bits_addr[2:0];
  wire  _isEcall_T = io_req_valid & system_ins;
  wire  isEcall = io_req_valid & system_ins & opcode[0];
  wire  is_break = _isEcall_T & opcode[1];
  wire  insn_ret = _isEcall_T & opcode[2];
  wire  isMret = io_req_valid & insn_ret & ~io_req_bits_addr[10];
  wire  _raiseExceptionVec_11_T = mode == 2'h3;
  wire  raiseExceptionVec_11 = mode == 2'h3 & isEcall;
  wire  raiseExceptionVec_8 = mode == 2'h0 & isEcall;
  wire [15:0] _raiseException_T = {4'h0,raiseExceptionVec_11,1'h0,1'h0,raiseExceptionVec_8,4'h0,is_break,1'h0,2'h0};
  wire  raiseException = |_raiseException_T;
  wire [3:0] _exceptionNO_T_6 = raiseExceptionVec_8 ? 4'h8 : 4'h0;
  wire [3:0] _exceptionNO_T_8 = raiseExceptionVec_11 ? 4'hb : _exceptionNO_T_6;
  wire [3:0] exceptionNO = is_break ? 4'h3 : _exceptionNO_T_8;
  wire  intrVecEnable_0 = mstatusStruct_IE_m & _raiseExceptionVec_11_T | mode < 2'h3;
  wire [5:0] intrVec_lo = {mip2_t_s,mip2_t_u,mip2_s_m,mip2_s_h,mip2_s_s,mip2_s_u};
  wire [11:0] _intrVec_T_1 = {mip2_e_m,mip2_e_h,mip2_e_s,mip2_e_u,mip2_t_m,mip2_t_h,intrVec_lo};
  wire [11:0] _intrVec_T_2 = reg_mie[11:0] & _intrVec_T_1;
  wire [5:0] intrVec_lo_1 = {intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,
    intrVecEnable_0};
  wire [11:0] _intrVec_T_3 = {intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,intrVecEnable_0,
    intrVecEnable_0,intrVec_lo_1};
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3;
  wire  raiseIntr = |intrVec;
  wire [2:0] _intrNO_T_1 = intrVec[4] ? 3'h4 : 3'h0;
  wire [3:0] _intrNO_T_3 = intrVec[8] ? 4'h8 : {{1'd0}, _intrNO_T_1};
  wire [3:0] _intrNO_T_5 = intrVec[0] ? 4'h0 : _intrNO_T_3;
  wire [3:0] _intrNO_T_7 = intrVec[5] ? 4'h5 : _intrNO_T_5;
  wire [3:0] _intrNO_T_9 = intrVec[9] ? 4'h9 : _intrNO_T_7;
  wire [3:0] _intrNO_T_11 = intrVec[1] ? 4'h1 : _intrNO_T_9;
  wire [3:0] _intrNO_T_13 = intrVec[7] ? 4'h7 : _intrNO_T_11;
  wire [3:0] _intrNO_T_15 = intrVec[11] ? 4'hb : _intrNO_T_13;
  wire [3:0] intrNO = intrVec[3] ? 4'h3 : _intrNO_T_15;
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0};
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO;
  wire [63:0] _GEN_1124 = {{60'd0}, _causeNO_T_1};
  wire [63:0] causeNO = _causeNO_T | _GEN_1124;
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_req_bits_valid;
  wire [10:0] reg_mstatus_lo = {mstatusStruct_reserved_2,mstatusStruct_SPP,mstatusStruct_IE_m,mstatusStruct_PIE_h,
    mstatusStruct_PIE_s,mstatusStruct_PIE_u,1'h0,mstatusStruct_IE_h,mstatusStruct_IE_s,mstatusStruct_IE_u};
  wire [7:0] reg_mstatus_hi_lo = {mstatusStruct_SUM,mstatusStruct_MPRV,mstatusStruct_XS,mstatusStruct_FS,mode};
  wire [63:0] _reg_mstatus_T = {mstatusStruct_SD,mstatusStruct_reserved,mstatusStruct_TSR,mstatusStruct_TW,
    mstatusStruct_TVM,mstatusStruct_MXR,reg_mstatus_hi_lo,reg_mstatus_lo};
  wire  _GEN_0 = raiseExceptionIntr ? causeNO[63] : reg_mcause_interrupt;
  wire [62:0] _GEN_1 = raiseExceptionIntr ? causeNO[62:0] : reg_mcause_exc_code;
  wire [63:0] _GEN_2 = raiseExceptionIntr ? {{32'd0}, io_req_bits_pc} : reg_mepc;
  wire [63:0] _GEN_4 = raiseExceptionIntr ? _reg_mstatus_T : reg_mstatus;
  wire [10:0] reg_mstatus_lo_1 = {mstatusStruct_reserved_2,mstatusStruct_SPP,1'h1,mstatusStruct_PIE_h,
    mstatusStruct_PIE_s,mstatusStruct_PIE_u,mstatusStruct_PIE_m,mstatusStruct_IE_h,mstatusStruct_IE_s,mstatusStruct_IE_u
    };
  wire [7:0] reg_mstatus_hi_lo_1 = {mstatusStruct_SUM,1'h0,mstatusStruct_XS,mstatusStruct_FS,2'h0};
  wire [63:0] _reg_mstatus_T_1 = {mstatusStruct_SD,mstatusStruct_reserved,mstatusStruct_TSR,mstatusStruct_TW,
    mstatusStruct_TVM,mstatusStruct_MXR,reg_mstatus_hi_lo_1,reg_mstatus_lo_1};
  wire [63:0] _GEN_6 = isMret ? _reg_mstatus_T_1 : _GEN_4;
  wire [63:0] _trapTarget_T_2 = {reg_mtvec_BASE,2'h0};
  wire [63:0] _trapTarget_T_7 = _trapTarget_T_2 + _read_csr_data_T_1;
  wire [65:0] _GEN_1125 = {_trapTarget_T_7, 2'h0};
  wire [66:0] _trapTarget_T_8 = {{1'd0}, _GEN_1125};
  wire [66:0] trapTarget = reg_mtvec_MODE == 2'h0 ? {{3'd0}, _trapTarget_T_2} : _trapTarget_T_8;
  wire [31:0] retTarget = reg_mepc[31:0];
  wire [66:0] _io_redirect_target_T = raiseExceptionIntr ? trapTarget : {{35'd0}, retTarget};
  wire [1:0] wMstatus_FS = write_data[14:13];
  wire  wMstatus_SD = write_data[63];
  wire  _reg_mstatus_T_2 = wMstatus_FS == 2'h3;
  wire [63:0] _reg_mstatus_T_4 = {_reg_mstatus_T_2,write_data[62:0]};
  wire  _T_20 = io_req_bits_addr == 12'h341;
  wire [75:0] _reg_mip_WIRE_2 = {{12'd0}, write_data};
  wire [63:0] _GEN_8 = io_req_bits_addr == 12'h3b0 ? write_data : reg_pmpaddr0;
  wire [63:0] _GEN_9 = io_req_bits_addr == 12'h3a3 ? write_data : reg_pmpcfg3;
  wire [63:0] _GEN_10 = io_req_bits_addr == 12'h3a3 ? reg_pmpaddr0 : _GEN_8;
  wire [63:0] _GEN_11 = io_req_bits_addr == 12'h3a2 ? write_data : reg_pmpcfg2;
  wire [63:0] _GEN_12 = io_req_bits_addr == 12'h3a2 ? reg_pmpcfg3 : _GEN_9;
  wire [63:0] _GEN_13 = io_req_bits_addr == 12'h3a2 ? reg_pmpaddr0 : _GEN_10;
  wire [63:0] _GEN_14 = io_req_bits_addr == 12'h3a1 ? write_data : reg_pmpcfg1;
  wire [63:0] _GEN_15 = io_req_bits_addr == 12'h3a1 ? reg_pmpcfg2 : _GEN_11;
  wire [63:0] _GEN_16 = io_req_bits_addr == 12'h3a1 ? reg_pmpcfg3 : _GEN_12;
  wire [63:0] _GEN_17 = io_req_bits_addr == 12'h3a1 ? reg_pmpaddr0 : _GEN_13;
  wire [63:0] _GEN_18 = io_req_bits_addr == 12'h3a0 ? write_data : reg_pmpcfg0;
  wire [63:0] _GEN_19 = io_req_bits_addr == 12'h3a0 ? reg_pmpcfg1 : _GEN_14;
  wire [63:0] _GEN_20 = io_req_bits_addr == 12'h3a0 ? reg_pmpcfg2 : _GEN_15;
  wire [63:0] _GEN_21 = io_req_bits_addr == 12'h3a0 ? reg_pmpcfg3 : _GEN_16;
  wire [63:0] _GEN_22 = io_req_bits_addr == 12'h3a0 ? reg_pmpaddr0 : _GEN_17;
  wire [63:0] _GEN_23 = _T_20 ? write_data : _GEN_2;
  wire [63:0] _GEN_24 = _T_20 ? reg_pmpcfg0 : _GEN_18;
  wire [63:0] _GEN_25 = _T_20 ? reg_pmpcfg1 : _GEN_19;
  wire [63:0] _GEN_26 = _T_20 ? reg_pmpcfg2 : _GEN_20;
  wire [63:0] _GEN_27 = _T_20 ? reg_pmpcfg3 : _GEN_21;
  wire [63:0] _GEN_28 = _T_20 ? reg_pmpaddr0 : _GEN_22;
  wire [51:0] _GEN_29 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[75:24] : reg_mip_reserved;
  wire  _GEN_30 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[23] : reg_mip_intr_e_m;
  wire  _GEN_31 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[22] : reg_mip_intr_e_h;
  wire  _GEN_32 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[21] : reg_mip_intr_e_s;
  wire  _GEN_33 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[20] : reg_mip_intr_e_u;
  wire  _GEN_34 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[19] : reg_mip_intr_t_m;
  wire  _GEN_35 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[18] : reg_mip_intr_t_h;
  wire  _GEN_36 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[17] : reg_mip_intr_t_s;
  wire  _GEN_37 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[16] : reg_mip_intr_t_u;
  wire  _GEN_38 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[15] : reg_mip_intr_s_m;
  wire  _GEN_39 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[14] : reg_mip_intr_s_h;
  wire  _GEN_40 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[13] : reg_mip_intr_s_s;
  wire  _GEN_41 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[12] : reg_mip_intr_s_u;
  wire  _GEN_42 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[11] : reg_mip_MEIP;
  wire  _GEN_43 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[10] : reg_mip_reserved_2;
  wire  _GEN_44 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[9] : reg_mip_SEIP;
  wire  _GEN_45 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[8] : reg_mip_UEIP;
  wire  _GEN_46 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[7] : reg_mip_MTIP;
  wire  _GEN_47 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[6] : reg_mip_reserved_3;
  wire  _GEN_48 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[5] : reg_mip_STIP;
  wire  _GEN_49 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[4] : reg_mip_UTIP;
  wire  _GEN_50 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[3] : reg_mip_MSIP;
  wire  _GEN_51 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[2] : reg_mip_reserved_4;
  wire  _GEN_52 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[1] : reg_mip_SSIP;
  wire  _GEN_53 = io_req_bits_addr == 12'h344 ? _reg_mip_WIRE_2[0] : reg_mip_USIP;
  wire [63:0] _GEN_54 = io_req_bits_addr == 12'h344 ? _GEN_2 : _GEN_23;
  wire [63:0] _GEN_55 = io_req_bits_addr == 12'h344 ? reg_pmpcfg0 : _GEN_24;
  wire [63:0] _GEN_56 = io_req_bits_addr == 12'h344 ? reg_pmpcfg1 : _GEN_25;
  wire [63:0] _GEN_57 = io_req_bits_addr == 12'h344 ? reg_pmpcfg2 : _GEN_26;
  wire [63:0] _GEN_58 = io_req_bits_addr == 12'h344 ? reg_pmpcfg3 : _GEN_27;
  wire [63:0] _GEN_59 = io_req_bits_addr == 12'h344 ? reg_pmpaddr0 : _GEN_28;
  wire [63:0] _GEN_60 = io_req_bits_addr == 12'h343 ? write_data : reg_mtval;
  wire [51:0] _GEN_61 = io_req_bits_addr == 12'h343 ? reg_mip_reserved : _GEN_29;
  wire  _GEN_62 = io_req_bits_addr == 12'h343 ? reg_mip_intr_e_m : _GEN_30;
  wire  _GEN_63 = io_req_bits_addr == 12'h343 ? reg_mip_intr_e_h : _GEN_31;
  wire  _GEN_64 = io_req_bits_addr == 12'h343 ? reg_mip_intr_e_s : _GEN_32;
  wire  _GEN_65 = io_req_bits_addr == 12'h343 ? reg_mip_intr_e_u : _GEN_33;
  wire  _GEN_66 = io_req_bits_addr == 12'h343 ? reg_mip_intr_t_m : _GEN_34;
  wire  _GEN_67 = io_req_bits_addr == 12'h343 ? reg_mip_intr_t_h : _GEN_35;
  wire  _GEN_68 = io_req_bits_addr == 12'h343 ? reg_mip_intr_t_s : _GEN_36;
  wire  _GEN_69 = io_req_bits_addr == 12'h343 ? reg_mip_intr_t_u : _GEN_37;
  wire  _GEN_70 = io_req_bits_addr == 12'h343 ? reg_mip_intr_s_m : _GEN_38;
  wire  _GEN_71 = io_req_bits_addr == 12'h343 ? reg_mip_intr_s_h : _GEN_39;
  wire  _GEN_72 = io_req_bits_addr == 12'h343 ? reg_mip_intr_s_s : _GEN_40;
  wire  _GEN_73 = io_req_bits_addr == 12'h343 ? reg_mip_intr_s_u : _GEN_41;
  wire  _GEN_74 = io_req_bits_addr == 12'h343 ? reg_mip_MEIP : _GEN_42;
  wire  _GEN_75 = io_req_bits_addr == 12'h343 ? reg_mip_reserved_2 : _GEN_43;
  wire  _GEN_76 = io_req_bits_addr == 12'h343 ? reg_mip_SEIP : _GEN_44;
  wire  _GEN_77 = io_req_bits_addr == 12'h343 ? reg_mip_UEIP : _GEN_45;
  wire  _GEN_78 = io_req_bits_addr == 12'h343 ? reg_mip_MTIP : _GEN_46;
  wire  _GEN_79 = io_req_bits_addr == 12'h343 ? reg_mip_reserved_3 : _GEN_47;
  wire  _GEN_80 = io_req_bits_addr == 12'h343 ? reg_mip_STIP : _GEN_48;
  wire  _GEN_81 = io_req_bits_addr == 12'h343 ? reg_mip_UTIP : _GEN_49;
  wire  _GEN_82 = io_req_bits_addr == 12'h343 ? reg_mip_MSIP : _GEN_50;
  wire  _GEN_83 = io_req_bits_addr == 12'h343 ? reg_mip_reserved_4 : _GEN_51;
  wire  _GEN_84 = io_req_bits_addr == 12'h343 ? reg_mip_SSIP : _GEN_52;
  wire  _GEN_85 = io_req_bits_addr == 12'h343 ? reg_mip_USIP : _GEN_53;
  wire [63:0] _GEN_86 = io_req_bits_addr == 12'h343 ? _GEN_2 : _GEN_54;
  wire [63:0] _GEN_87 = io_req_bits_addr == 12'h343 ? reg_pmpcfg0 : _GEN_55;
  wire [63:0] _GEN_88 = io_req_bits_addr == 12'h343 ? reg_pmpcfg1 : _GEN_56;
  wire [63:0] _GEN_89 = io_req_bits_addr == 12'h343 ? reg_pmpcfg2 : _GEN_57;
  wire [63:0] _GEN_90 = io_req_bits_addr == 12'h343 ? reg_pmpcfg3 : _GEN_58;
  wire [63:0] _GEN_91 = io_req_bits_addr == 12'h343 ? reg_pmpaddr0 : _GEN_59;
  wire  _GEN_92 = io_req_bits_addr == 12'h342 ? wMstatus_SD : _GEN_0;
  wire [62:0] _GEN_93 = io_req_bits_addr == 12'h342 ? write_data[62:0] : _GEN_1;
  wire [63:0] _GEN_94 = io_req_bits_addr == 12'h342 ? reg_mtval : _GEN_60;
  wire [51:0] _GEN_95 = io_req_bits_addr == 12'h342 ? reg_mip_reserved : _GEN_61;
  wire  _GEN_96 = io_req_bits_addr == 12'h342 ? reg_mip_intr_e_m : _GEN_62;
  wire  _GEN_97 = io_req_bits_addr == 12'h342 ? reg_mip_intr_e_h : _GEN_63;
  wire  _GEN_98 = io_req_bits_addr == 12'h342 ? reg_mip_intr_e_s : _GEN_64;
  wire  _GEN_99 = io_req_bits_addr == 12'h342 ? reg_mip_intr_e_u : _GEN_65;
  wire  _GEN_100 = io_req_bits_addr == 12'h342 ? reg_mip_intr_t_m : _GEN_66;
  wire  _GEN_101 = io_req_bits_addr == 12'h342 ? reg_mip_intr_t_h : _GEN_67;
  wire  _GEN_102 = io_req_bits_addr == 12'h342 ? reg_mip_intr_t_s : _GEN_68;
  wire  _GEN_103 = io_req_bits_addr == 12'h342 ? reg_mip_intr_t_u : _GEN_69;
  wire  _GEN_104 = io_req_bits_addr == 12'h342 ? reg_mip_intr_s_m : _GEN_70;
  wire  _GEN_105 = io_req_bits_addr == 12'h342 ? reg_mip_intr_s_h : _GEN_71;
  wire  _GEN_106 = io_req_bits_addr == 12'h342 ? reg_mip_intr_s_s : _GEN_72;
  wire  _GEN_107 = io_req_bits_addr == 12'h342 ? reg_mip_intr_s_u : _GEN_73;
  wire  _GEN_108 = io_req_bits_addr == 12'h342 ? reg_mip_MEIP : _GEN_74;
  wire  _GEN_109 = io_req_bits_addr == 12'h342 ? reg_mip_reserved_2 : _GEN_75;
  wire  _GEN_110 = io_req_bits_addr == 12'h342 ? reg_mip_SEIP : _GEN_76;
  wire  _GEN_111 = io_req_bits_addr == 12'h342 ? reg_mip_UEIP : _GEN_77;
  wire  _GEN_112 = io_req_bits_addr == 12'h342 ? reg_mip_MTIP : _GEN_78;
  wire  _GEN_113 = io_req_bits_addr == 12'h342 ? reg_mip_reserved_3 : _GEN_79;
  wire  _GEN_114 = io_req_bits_addr == 12'h342 ? reg_mip_STIP : _GEN_80;
  wire  _GEN_115 = io_req_bits_addr == 12'h342 ? reg_mip_UTIP : _GEN_81;
  wire  _GEN_116 = io_req_bits_addr == 12'h342 ? reg_mip_MSIP : _GEN_82;
  wire  _GEN_117 = io_req_bits_addr == 12'h342 ? reg_mip_reserved_4 : _GEN_83;
  wire  _GEN_118 = io_req_bits_addr == 12'h342 ? reg_mip_SSIP : _GEN_84;
  wire  _GEN_119 = io_req_bits_addr == 12'h342 ? reg_mip_USIP : _GEN_85;
  wire [63:0] _GEN_120 = io_req_bits_addr == 12'h342 ? _GEN_2 : _GEN_86;
  wire [63:0] _GEN_121 = io_req_bits_addr == 12'h342 ? reg_pmpcfg0 : _GEN_87;
  wire [63:0] _GEN_122 = io_req_bits_addr == 12'h342 ? reg_pmpcfg1 : _GEN_88;
  wire [63:0] _GEN_123 = io_req_bits_addr == 12'h342 ? reg_pmpcfg2 : _GEN_89;
  wire [63:0] _GEN_124 = io_req_bits_addr == 12'h342 ? reg_pmpcfg3 : _GEN_90;
  wire [63:0] _GEN_125 = io_req_bits_addr == 12'h342 ? reg_pmpaddr0 : _GEN_91;
  wire [63:0] _GEN_126 = io_req_bits_addr == 12'h341 ? write_data : _GEN_120;
  wire  _GEN_127 = io_req_bits_addr == 12'h341 ? _GEN_0 : _GEN_92;
  wire [62:0] _GEN_128 = io_req_bits_addr == 12'h341 ? _GEN_1 : _GEN_93;
  wire [63:0] _GEN_129 = io_req_bits_addr == 12'h341 ? reg_mtval : _GEN_94;
  wire [51:0] _GEN_130 = io_req_bits_addr == 12'h341 ? reg_mip_reserved : _GEN_95;
  wire  _GEN_131 = io_req_bits_addr == 12'h341 ? reg_mip_intr_e_m : _GEN_96;
  wire  _GEN_132 = io_req_bits_addr == 12'h341 ? reg_mip_intr_e_h : _GEN_97;
  wire  _GEN_133 = io_req_bits_addr == 12'h341 ? reg_mip_intr_e_s : _GEN_98;
  wire  _GEN_134 = io_req_bits_addr == 12'h341 ? reg_mip_intr_e_u : _GEN_99;
  wire  _GEN_135 = io_req_bits_addr == 12'h341 ? reg_mip_intr_t_m : _GEN_100;
  wire  _GEN_136 = io_req_bits_addr == 12'h341 ? reg_mip_intr_t_h : _GEN_101;
  wire  _GEN_137 = io_req_bits_addr == 12'h341 ? reg_mip_intr_t_s : _GEN_102;
  wire  _GEN_138 = io_req_bits_addr == 12'h341 ? reg_mip_intr_t_u : _GEN_103;
  wire  _GEN_139 = io_req_bits_addr == 12'h341 ? reg_mip_intr_s_m : _GEN_104;
  wire  _GEN_140 = io_req_bits_addr == 12'h341 ? reg_mip_intr_s_h : _GEN_105;
  wire  _GEN_141 = io_req_bits_addr == 12'h341 ? reg_mip_intr_s_s : _GEN_106;
  wire  _GEN_142 = io_req_bits_addr == 12'h341 ? reg_mip_intr_s_u : _GEN_107;
  wire  _GEN_143 = io_req_bits_addr == 12'h341 ? reg_mip_MEIP : _GEN_108;
  wire  _GEN_144 = io_req_bits_addr == 12'h341 ? reg_mip_reserved_2 : _GEN_109;
  wire  _GEN_145 = io_req_bits_addr == 12'h341 ? reg_mip_SEIP : _GEN_110;
  wire  _GEN_146 = io_req_bits_addr == 12'h341 ? reg_mip_UEIP : _GEN_111;
  wire  _GEN_147 = io_req_bits_addr == 12'h341 ? reg_mip_MTIP : _GEN_112;
  wire  _GEN_148 = io_req_bits_addr == 12'h341 ? reg_mip_reserved_3 : _GEN_113;
  wire  _GEN_149 = io_req_bits_addr == 12'h341 ? reg_mip_STIP : _GEN_114;
  wire  _GEN_150 = io_req_bits_addr == 12'h341 ? reg_mip_UTIP : _GEN_115;
  wire  _GEN_151 = io_req_bits_addr == 12'h341 ? reg_mip_MSIP : _GEN_116;
  wire  _GEN_152 = io_req_bits_addr == 12'h341 ? reg_mip_reserved_4 : _GEN_117;
  wire  _GEN_153 = io_req_bits_addr == 12'h341 ? reg_mip_SSIP : _GEN_118;
  wire  _GEN_154 = io_req_bits_addr == 12'h341 ? reg_mip_USIP : _GEN_119;
  wire [63:0] _GEN_155 = io_req_bits_addr == 12'h341 ? reg_pmpcfg0 : _GEN_121;
  wire [63:0] _GEN_156 = io_req_bits_addr == 12'h341 ? reg_pmpcfg1 : _GEN_122;
  wire [63:0] _GEN_157 = io_req_bits_addr == 12'h341 ? reg_pmpcfg2 : _GEN_123;
  wire [63:0] _GEN_158 = io_req_bits_addr == 12'h341 ? reg_pmpcfg3 : _GEN_124;
  wire [63:0] _GEN_159 = io_req_bits_addr == 12'h341 ? reg_pmpaddr0 : _GEN_125;
  wire [63:0] _GEN_160 = io_req_bits_addr == 12'h340 ? write_data : reg_mscratch;
  wire [63:0] _GEN_161 = io_req_bits_addr == 12'h340 ? _GEN_2 : _GEN_126;
  wire  _GEN_162 = io_req_bits_addr == 12'h340 ? _GEN_0 : _GEN_127;
  wire [62:0] _GEN_163 = io_req_bits_addr == 12'h340 ? _GEN_1 : _GEN_128;
  wire [63:0] _GEN_164 = io_req_bits_addr == 12'h340 ? reg_mtval : _GEN_129;
  wire [51:0] _GEN_165 = io_req_bits_addr == 12'h340 ? reg_mip_reserved : _GEN_130;
  wire  _GEN_166 = io_req_bits_addr == 12'h340 ? reg_mip_intr_e_m : _GEN_131;
  wire  _GEN_167 = io_req_bits_addr == 12'h340 ? reg_mip_intr_e_h : _GEN_132;
  wire  _GEN_168 = io_req_bits_addr == 12'h340 ? reg_mip_intr_e_s : _GEN_133;
  wire  _GEN_169 = io_req_bits_addr == 12'h340 ? reg_mip_intr_e_u : _GEN_134;
  wire  _GEN_170 = io_req_bits_addr == 12'h340 ? reg_mip_intr_t_m : _GEN_135;
  wire  _GEN_171 = io_req_bits_addr == 12'h340 ? reg_mip_intr_t_h : _GEN_136;
  wire  _GEN_172 = io_req_bits_addr == 12'h340 ? reg_mip_intr_t_s : _GEN_137;
  wire  _GEN_173 = io_req_bits_addr == 12'h340 ? reg_mip_intr_t_u : _GEN_138;
  wire  _GEN_174 = io_req_bits_addr == 12'h340 ? reg_mip_intr_s_m : _GEN_139;
  wire  _GEN_175 = io_req_bits_addr == 12'h340 ? reg_mip_intr_s_h : _GEN_140;
  wire  _GEN_176 = io_req_bits_addr == 12'h340 ? reg_mip_intr_s_s : _GEN_141;
  wire  _GEN_177 = io_req_bits_addr == 12'h340 ? reg_mip_intr_s_u : _GEN_142;
  wire  _GEN_178 = io_req_bits_addr == 12'h340 ? reg_mip_MEIP : _GEN_143;
  wire  _GEN_179 = io_req_bits_addr == 12'h340 ? reg_mip_reserved_2 : _GEN_144;
  wire  _GEN_180 = io_req_bits_addr == 12'h340 ? reg_mip_SEIP : _GEN_145;
  wire  _GEN_181 = io_req_bits_addr == 12'h340 ? reg_mip_UEIP : _GEN_146;
  wire  _GEN_182 = io_req_bits_addr == 12'h340 ? reg_mip_MTIP : _GEN_147;
  wire  _GEN_183 = io_req_bits_addr == 12'h340 ? reg_mip_reserved_3 : _GEN_148;
  wire  _GEN_184 = io_req_bits_addr == 12'h340 ? reg_mip_STIP : _GEN_149;
  wire  _GEN_185 = io_req_bits_addr == 12'h340 ? reg_mip_UTIP : _GEN_150;
  wire  _GEN_186 = io_req_bits_addr == 12'h340 ? reg_mip_MSIP : _GEN_151;
  wire  _GEN_187 = io_req_bits_addr == 12'h340 ? reg_mip_reserved_4 : _GEN_152;
  wire  _GEN_188 = io_req_bits_addr == 12'h340 ? reg_mip_SSIP : _GEN_153;
  wire  _GEN_189 = io_req_bits_addr == 12'h340 ? reg_mip_USIP : _GEN_154;
  wire [63:0] _GEN_190 = io_req_bits_addr == 12'h340 ? reg_pmpcfg0 : _GEN_155;
  wire [63:0] _GEN_191 = io_req_bits_addr == 12'h340 ? reg_pmpcfg1 : _GEN_156;
  wire [63:0] _GEN_192 = io_req_bits_addr == 12'h340 ? reg_pmpcfg2 : _GEN_157;
  wire [63:0] _GEN_193 = io_req_bits_addr == 12'h340 ? reg_pmpcfg3 : _GEN_158;
  wire [63:0] _GEN_194 = io_req_bits_addr == 12'h340 ? reg_pmpaddr0 : _GEN_159;
  wire [61:0] _GEN_195 = io_req_bits_addr == 12'h305 ? write_data[63:2] : reg_mtvec_BASE;
  wire [1:0] _GEN_196 = io_req_bits_addr == 12'h305 ? write_data[1:0] : reg_mtvec_MODE;
  wire [63:0] _GEN_197 = io_req_bits_addr == 12'h305 ? reg_mscratch : _GEN_160;
  wire [63:0] _GEN_198 = io_req_bits_addr == 12'h305 ? _GEN_2 : _GEN_161;
  wire  _GEN_199 = io_req_bits_addr == 12'h305 ? _GEN_0 : _GEN_162;
  wire [62:0] _GEN_200 = io_req_bits_addr == 12'h305 ? _GEN_1 : _GEN_163;
  wire [63:0] _GEN_201 = io_req_bits_addr == 12'h305 ? reg_mtval : _GEN_164;
  wire [51:0] _GEN_202 = io_req_bits_addr == 12'h305 ? reg_mip_reserved : _GEN_165;
  wire  _GEN_203 = io_req_bits_addr == 12'h305 ? reg_mip_intr_e_m : _GEN_166;
  wire  _GEN_204 = io_req_bits_addr == 12'h305 ? reg_mip_intr_e_h : _GEN_167;
  wire  _GEN_205 = io_req_bits_addr == 12'h305 ? reg_mip_intr_e_s : _GEN_168;
  wire  _GEN_206 = io_req_bits_addr == 12'h305 ? reg_mip_intr_e_u : _GEN_169;
  wire  _GEN_207 = io_req_bits_addr == 12'h305 ? reg_mip_intr_t_m : _GEN_170;
  wire  _GEN_208 = io_req_bits_addr == 12'h305 ? reg_mip_intr_t_h : _GEN_171;
  wire  _GEN_209 = io_req_bits_addr == 12'h305 ? reg_mip_intr_t_s : _GEN_172;
  wire  _GEN_210 = io_req_bits_addr == 12'h305 ? reg_mip_intr_t_u : _GEN_173;
  wire  _GEN_211 = io_req_bits_addr == 12'h305 ? reg_mip_intr_s_m : _GEN_174;
  wire  _GEN_212 = io_req_bits_addr == 12'h305 ? reg_mip_intr_s_h : _GEN_175;
  wire  _GEN_213 = io_req_bits_addr == 12'h305 ? reg_mip_intr_s_s : _GEN_176;
  wire  _GEN_214 = io_req_bits_addr == 12'h305 ? reg_mip_intr_s_u : _GEN_177;
  wire  _GEN_215 = io_req_bits_addr == 12'h305 ? reg_mip_MEIP : _GEN_178;
  wire  _GEN_216 = io_req_bits_addr == 12'h305 ? reg_mip_reserved_2 : _GEN_179;
  wire  _GEN_217 = io_req_bits_addr == 12'h305 ? reg_mip_SEIP : _GEN_180;
  wire  _GEN_218 = io_req_bits_addr == 12'h305 ? reg_mip_UEIP : _GEN_181;
  wire  _GEN_219 = io_req_bits_addr == 12'h305 ? reg_mip_MTIP : _GEN_182;
  wire  _GEN_220 = io_req_bits_addr == 12'h305 ? reg_mip_reserved_3 : _GEN_183;
  wire  _GEN_221 = io_req_bits_addr == 12'h305 ? reg_mip_STIP : _GEN_184;
  wire  _GEN_222 = io_req_bits_addr == 12'h305 ? reg_mip_UTIP : _GEN_185;
  wire  _GEN_223 = io_req_bits_addr == 12'h305 ? reg_mip_MSIP : _GEN_186;
  wire  _GEN_224 = io_req_bits_addr == 12'h305 ? reg_mip_reserved_4 : _GEN_187;
  wire  _GEN_225 = io_req_bits_addr == 12'h305 ? reg_mip_SSIP : _GEN_188;
  wire  _GEN_226 = io_req_bits_addr == 12'h305 ? reg_mip_USIP : _GEN_189;
  wire [63:0] _GEN_227 = io_req_bits_addr == 12'h305 ? reg_pmpcfg0 : _GEN_190;
  wire [63:0] _GEN_228 = io_req_bits_addr == 12'h305 ? reg_pmpcfg1 : _GEN_191;
  wire [63:0] _GEN_229 = io_req_bits_addr == 12'h305 ? reg_pmpcfg2 : _GEN_192;
  wire [63:0] _GEN_230 = io_req_bits_addr == 12'h305 ? reg_pmpcfg3 : _GEN_193;
  wire [63:0] _GEN_231 = io_req_bits_addr == 12'h305 ? reg_pmpaddr0 : _GEN_194;
  wire [63:0] _GEN_232 = io_req_bits_addr == 12'h304 ? write_data : reg_mie;
  wire [61:0] _GEN_233 = io_req_bits_addr == 12'h304 ? reg_mtvec_BASE : _GEN_195;
  wire [1:0] _GEN_234 = io_req_bits_addr == 12'h304 ? reg_mtvec_MODE : _GEN_196;
  wire [63:0] _GEN_235 = io_req_bits_addr == 12'h304 ? reg_mscratch : _GEN_197;
  wire [63:0] _GEN_236 = io_req_bits_addr == 12'h304 ? _GEN_2 : _GEN_198;
  wire  _GEN_237 = io_req_bits_addr == 12'h304 ? _GEN_0 : _GEN_199;
  wire [62:0] _GEN_238 = io_req_bits_addr == 12'h304 ? _GEN_1 : _GEN_200;
  wire [63:0] _GEN_239 = io_req_bits_addr == 12'h304 ? reg_mtval : _GEN_201;
  wire [51:0] _GEN_240 = io_req_bits_addr == 12'h304 ? reg_mip_reserved : _GEN_202;
  wire  _GEN_241 = io_req_bits_addr == 12'h304 ? reg_mip_intr_e_m : _GEN_203;
  wire  _GEN_242 = io_req_bits_addr == 12'h304 ? reg_mip_intr_e_h : _GEN_204;
  wire  _GEN_243 = io_req_bits_addr == 12'h304 ? reg_mip_intr_e_s : _GEN_205;
  wire  _GEN_244 = io_req_bits_addr == 12'h304 ? reg_mip_intr_e_u : _GEN_206;
  wire  _GEN_245 = io_req_bits_addr == 12'h304 ? reg_mip_intr_t_m : _GEN_207;
  wire  _GEN_246 = io_req_bits_addr == 12'h304 ? reg_mip_intr_t_h : _GEN_208;
  wire  _GEN_247 = io_req_bits_addr == 12'h304 ? reg_mip_intr_t_s : _GEN_209;
  wire  _GEN_248 = io_req_bits_addr == 12'h304 ? reg_mip_intr_t_u : _GEN_210;
  wire  _GEN_249 = io_req_bits_addr == 12'h304 ? reg_mip_intr_s_m : _GEN_211;
  wire  _GEN_250 = io_req_bits_addr == 12'h304 ? reg_mip_intr_s_h : _GEN_212;
  wire  _GEN_251 = io_req_bits_addr == 12'h304 ? reg_mip_intr_s_s : _GEN_213;
  wire  _GEN_252 = io_req_bits_addr == 12'h304 ? reg_mip_intr_s_u : _GEN_214;
  wire  _GEN_253 = io_req_bits_addr == 12'h304 ? reg_mip_MEIP : _GEN_215;
  wire  _GEN_254 = io_req_bits_addr == 12'h304 ? reg_mip_reserved_2 : _GEN_216;
  wire  _GEN_255 = io_req_bits_addr == 12'h304 ? reg_mip_SEIP : _GEN_217;
  wire  _GEN_256 = io_req_bits_addr == 12'h304 ? reg_mip_UEIP : _GEN_218;
  wire  _GEN_257 = io_req_bits_addr == 12'h304 ? reg_mip_MTIP : _GEN_219;
  wire  _GEN_258 = io_req_bits_addr == 12'h304 ? reg_mip_reserved_3 : _GEN_220;
  wire  _GEN_259 = io_req_bits_addr == 12'h304 ? reg_mip_STIP : _GEN_221;
  wire  _GEN_260 = io_req_bits_addr == 12'h304 ? reg_mip_UTIP : _GEN_222;
  wire  _GEN_261 = io_req_bits_addr == 12'h304 ? reg_mip_MSIP : _GEN_223;
  wire  _GEN_262 = io_req_bits_addr == 12'h304 ? reg_mip_reserved_4 : _GEN_224;
  wire  _GEN_263 = io_req_bits_addr == 12'h304 ? reg_mip_SSIP : _GEN_225;
  wire  _GEN_264 = io_req_bits_addr == 12'h304 ? reg_mip_USIP : _GEN_226;
  wire [63:0] _GEN_265 = io_req_bits_addr == 12'h304 ? reg_pmpcfg0 : _GEN_227;
  wire [63:0] _GEN_266 = io_req_bits_addr == 12'h304 ? reg_pmpcfg1 : _GEN_228;
  wire [63:0] _GEN_267 = io_req_bits_addr == 12'h304 ? reg_pmpcfg2 : _GEN_229;
  wire [63:0] _GEN_268 = io_req_bits_addr == 12'h304 ? reg_pmpcfg3 : _GEN_230;
  wire [63:0] _GEN_269 = io_req_bits_addr == 12'h304 ? reg_pmpaddr0 : _GEN_231;
  wire [63:0] _GEN_270 = io_req_bits_addr == 12'h303 ? write_data : reg_mideleg;
  wire [63:0] _GEN_271 = io_req_bits_addr == 12'h303 ? reg_mie : _GEN_232;
  wire [61:0] _GEN_272 = io_req_bits_addr == 12'h303 ? reg_mtvec_BASE : _GEN_233;
  wire [1:0] _GEN_273 = io_req_bits_addr == 12'h303 ? reg_mtvec_MODE : _GEN_234;
  wire [63:0] _GEN_274 = io_req_bits_addr == 12'h303 ? reg_mscratch : _GEN_235;
  wire [63:0] _GEN_275 = io_req_bits_addr == 12'h303 ? _GEN_2 : _GEN_236;
  wire  _GEN_276 = io_req_bits_addr == 12'h303 ? _GEN_0 : _GEN_237;
  wire [62:0] _GEN_277 = io_req_bits_addr == 12'h303 ? _GEN_1 : _GEN_238;
  wire [63:0] _GEN_278 = io_req_bits_addr == 12'h303 ? reg_mtval : _GEN_239;
  wire [51:0] _GEN_279 = io_req_bits_addr == 12'h303 ? reg_mip_reserved : _GEN_240;
  wire  _GEN_280 = io_req_bits_addr == 12'h303 ? reg_mip_intr_e_m : _GEN_241;
  wire  _GEN_281 = io_req_bits_addr == 12'h303 ? reg_mip_intr_e_h : _GEN_242;
  wire  _GEN_282 = io_req_bits_addr == 12'h303 ? reg_mip_intr_e_s : _GEN_243;
  wire  _GEN_283 = io_req_bits_addr == 12'h303 ? reg_mip_intr_e_u : _GEN_244;
  wire  _GEN_284 = io_req_bits_addr == 12'h303 ? reg_mip_intr_t_m : _GEN_245;
  wire  _GEN_285 = io_req_bits_addr == 12'h303 ? reg_mip_intr_t_h : _GEN_246;
  wire  _GEN_286 = io_req_bits_addr == 12'h303 ? reg_mip_intr_t_s : _GEN_247;
  wire  _GEN_287 = io_req_bits_addr == 12'h303 ? reg_mip_intr_t_u : _GEN_248;
  wire  _GEN_288 = io_req_bits_addr == 12'h303 ? reg_mip_intr_s_m : _GEN_249;
  wire  _GEN_289 = io_req_bits_addr == 12'h303 ? reg_mip_intr_s_h : _GEN_250;
  wire  _GEN_290 = io_req_bits_addr == 12'h303 ? reg_mip_intr_s_s : _GEN_251;
  wire  _GEN_291 = io_req_bits_addr == 12'h303 ? reg_mip_intr_s_u : _GEN_252;
  wire  _GEN_292 = io_req_bits_addr == 12'h303 ? reg_mip_MEIP : _GEN_253;
  wire  _GEN_293 = io_req_bits_addr == 12'h303 ? reg_mip_reserved_2 : _GEN_254;
  wire  _GEN_294 = io_req_bits_addr == 12'h303 ? reg_mip_SEIP : _GEN_255;
  wire  _GEN_295 = io_req_bits_addr == 12'h303 ? reg_mip_UEIP : _GEN_256;
  wire  _GEN_296 = io_req_bits_addr == 12'h303 ? reg_mip_MTIP : _GEN_257;
  wire  _GEN_297 = io_req_bits_addr == 12'h303 ? reg_mip_reserved_3 : _GEN_258;
  wire  _GEN_298 = io_req_bits_addr == 12'h303 ? reg_mip_STIP : _GEN_259;
  wire  _GEN_299 = io_req_bits_addr == 12'h303 ? reg_mip_UTIP : _GEN_260;
  wire  _GEN_300 = io_req_bits_addr == 12'h303 ? reg_mip_MSIP : _GEN_261;
  wire  _GEN_301 = io_req_bits_addr == 12'h303 ? reg_mip_reserved_4 : _GEN_262;
  wire  _GEN_302 = io_req_bits_addr == 12'h303 ? reg_mip_SSIP : _GEN_263;
  wire  _GEN_303 = io_req_bits_addr == 12'h303 ? reg_mip_USIP : _GEN_264;
  wire [63:0] _GEN_304 = io_req_bits_addr == 12'h303 ? reg_pmpcfg0 : _GEN_265;
  wire [63:0] _GEN_305 = io_req_bits_addr == 12'h303 ? reg_pmpcfg1 : _GEN_266;
  wire [63:0] _GEN_306 = io_req_bits_addr == 12'h303 ? reg_pmpcfg2 : _GEN_267;
  wire [63:0] _GEN_307 = io_req_bits_addr == 12'h303 ? reg_pmpcfg3 : _GEN_268;
  wire [63:0] _GEN_308 = io_req_bits_addr == 12'h303 ? reg_pmpaddr0 : _GEN_269;
  wire [63:0] _GEN_309 = io_req_bits_addr == 12'h302 ? write_data : reg_medeleg;
  wire [63:0] _GEN_310 = io_req_bits_addr == 12'h302 ? reg_mideleg : _GEN_270;
  wire [63:0] _GEN_311 = io_req_bits_addr == 12'h302 ? reg_mie : _GEN_271;
  wire [61:0] _GEN_312 = io_req_bits_addr == 12'h302 ? reg_mtvec_BASE : _GEN_272;
  wire [1:0] _GEN_313 = io_req_bits_addr == 12'h302 ? reg_mtvec_MODE : _GEN_273;
  wire [63:0] _GEN_314 = io_req_bits_addr == 12'h302 ? reg_mscratch : _GEN_274;
  wire [63:0] _GEN_315 = io_req_bits_addr == 12'h302 ? _GEN_2 : _GEN_275;
  wire  _GEN_316 = io_req_bits_addr == 12'h302 ? _GEN_0 : _GEN_276;
  wire [62:0] _GEN_317 = io_req_bits_addr == 12'h302 ? _GEN_1 : _GEN_277;
  wire [63:0] _GEN_318 = io_req_bits_addr == 12'h302 ? reg_mtval : _GEN_278;
  wire [51:0] _GEN_319 = io_req_bits_addr == 12'h302 ? reg_mip_reserved : _GEN_279;
  wire  _GEN_320 = io_req_bits_addr == 12'h302 ? reg_mip_intr_e_m : _GEN_280;
  wire  _GEN_321 = io_req_bits_addr == 12'h302 ? reg_mip_intr_e_h : _GEN_281;
  wire  _GEN_322 = io_req_bits_addr == 12'h302 ? reg_mip_intr_e_s : _GEN_282;
  wire  _GEN_323 = io_req_bits_addr == 12'h302 ? reg_mip_intr_e_u : _GEN_283;
  wire  _GEN_324 = io_req_bits_addr == 12'h302 ? reg_mip_intr_t_m : _GEN_284;
  wire  _GEN_325 = io_req_bits_addr == 12'h302 ? reg_mip_intr_t_h : _GEN_285;
  wire  _GEN_326 = io_req_bits_addr == 12'h302 ? reg_mip_intr_t_s : _GEN_286;
  wire  _GEN_327 = io_req_bits_addr == 12'h302 ? reg_mip_intr_t_u : _GEN_287;
  wire  _GEN_328 = io_req_bits_addr == 12'h302 ? reg_mip_intr_s_m : _GEN_288;
  wire  _GEN_329 = io_req_bits_addr == 12'h302 ? reg_mip_intr_s_h : _GEN_289;
  wire  _GEN_330 = io_req_bits_addr == 12'h302 ? reg_mip_intr_s_s : _GEN_290;
  wire  _GEN_331 = io_req_bits_addr == 12'h302 ? reg_mip_intr_s_u : _GEN_291;
  wire  _GEN_332 = io_req_bits_addr == 12'h302 ? reg_mip_MEIP : _GEN_292;
  wire  _GEN_333 = io_req_bits_addr == 12'h302 ? reg_mip_reserved_2 : _GEN_293;
  wire  _GEN_334 = io_req_bits_addr == 12'h302 ? reg_mip_SEIP : _GEN_294;
  wire  _GEN_335 = io_req_bits_addr == 12'h302 ? reg_mip_UEIP : _GEN_295;
  wire  _GEN_336 = io_req_bits_addr == 12'h302 ? reg_mip_MTIP : _GEN_296;
  wire  _GEN_337 = io_req_bits_addr == 12'h302 ? reg_mip_reserved_3 : _GEN_297;
  wire  _GEN_338 = io_req_bits_addr == 12'h302 ? reg_mip_STIP : _GEN_298;
  wire  _GEN_339 = io_req_bits_addr == 12'h302 ? reg_mip_UTIP : _GEN_299;
  wire  _GEN_340 = io_req_bits_addr == 12'h302 ? reg_mip_MSIP : _GEN_300;
  wire  _GEN_341 = io_req_bits_addr == 12'h302 ? reg_mip_reserved_4 : _GEN_301;
  wire  _GEN_342 = io_req_bits_addr == 12'h302 ? reg_mip_SSIP : _GEN_302;
  wire  _GEN_343 = io_req_bits_addr == 12'h302 ? reg_mip_USIP : _GEN_303;
  wire [63:0] _GEN_344 = io_req_bits_addr == 12'h302 ? reg_pmpcfg0 : _GEN_304;
  wire [63:0] _GEN_345 = io_req_bits_addr == 12'h302 ? reg_pmpcfg1 : _GEN_305;
  wire [63:0] _GEN_346 = io_req_bits_addr == 12'h302 ? reg_pmpcfg2 : _GEN_306;
  wire [63:0] _GEN_347 = io_req_bits_addr == 12'h302 ? reg_pmpcfg3 : _GEN_307;
  wire [63:0] _GEN_348 = io_req_bits_addr == 12'h302 ? reg_pmpaddr0 : _GEN_308;
  wire [63:0] _GEN_349 = io_req_bits_addr == 12'h301 ? write_data : reg_misa;
  wire [63:0] _GEN_350 = io_req_bits_addr == 12'h301 ? reg_medeleg : _GEN_309;
  wire [63:0] _GEN_351 = io_req_bits_addr == 12'h301 ? reg_mideleg : _GEN_310;
  wire [63:0] _GEN_352 = io_req_bits_addr == 12'h301 ? reg_mie : _GEN_311;
  wire [61:0] _GEN_353 = io_req_bits_addr == 12'h301 ? reg_mtvec_BASE : _GEN_312;
  wire [1:0] _GEN_354 = io_req_bits_addr == 12'h301 ? reg_mtvec_MODE : _GEN_313;
  wire [63:0] _GEN_355 = io_req_bits_addr == 12'h301 ? reg_mscratch : _GEN_314;
  wire [63:0] _GEN_356 = io_req_bits_addr == 12'h301 ? _GEN_2 : _GEN_315;
  wire  _GEN_357 = io_req_bits_addr == 12'h301 ? _GEN_0 : _GEN_316;
  wire [62:0] _GEN_358 = io_req_bits_addr == 12'h301 ? _GEN_1 : _GEN_317;
  wire [63:0] _GEN_359 = io_req_bits_addr == 12'h301 ? reg_mtval : _GEN_318;
  wire [51:0] _GEN_360 = io_req_bits_addr == 12'h301 ? reg_mip_reserved : _GEN_319;
  wire  _GEN_361 = io_req_bits_addr == 12'h301 ? reg_mip_intr_e_m : _GEN_320;
  wire  _GEN_362 = io_req_bits_addr == 12'h301 ? reg_mip_intr_e_h : _GEN_321;
  wire  _GEN_363 = io_req_bits_addr == 12'h301 ? reg_mip_intr_e_s : _GEN_322;
  wire  _GEN_364 = io_req_bits_addr == 12'h301 ? reg_mip_intr_e_u : _GEN_323;
  wire  _GEN_365 = io_req_bits_addr == 12'h301 ? reg_mip_intr_t_m : _GEN_324;
  wire  _GEN_366 = io_req_bits_addr == 12'h301 ? reg_mip_intr_t_h : _GEN_325;
  wire  _GEN_367 = io_req_bits_addr == 12'h301 ? reg_mip_intr_t_s : _GEN_326;
  wire  _GEN_368 = io_req_bits_addr == 12'h301 ? reg_mip_intr_t_u : _GEN_327;
  wire  _GEN_369 = io_req_bits_addr == 12'h301 ? reg_mip_intr_s_m : _GEN_328;
  wire  _GEN_370 = io_req_bits_addr == 12'h301 ? reg_mip_intr_s_h : _GEN_329;
  wire  _GEN_371 = io_req_bits_addr == 12'h301 ? reg_mip_intr_s_s : _GEN_330;
  wire  _GEN_372 = io_req_bits_addr == 12'h301 ? reg_mip_intr_s_u : _GEN_331;
  wire  _GEN_373 = io_req_bits_addr == 12'h301 ? reg_mip_MEIP : _GEN_332;
  wire  _GEN_374 = io_req_bits_addr == 12'h301 ? reg_mip_reserved_2 : _GEN_333;
  wire  _GEN_375 = io_req_bits_addr == 12'h301 ? reg_mip_SEIP : _GEN_334;
  wire  _GEN_376 = io_req_bits_addr == 12'h301 ? reg_mip_UEIP : _GEN_335;
  wire  _GEN_377 = io_req_bits_addr == 12'h301 ? reg_mip_MTIP : _GEN_336;
  wire  _GEN_378 = io_req_bits_addr == 12'h301 ? reg_mip_reserved_3 : _GEN_337;
  wire  _GEN_379 = io_req_bits_addr == 12'h301 ? reg_mip_STIP : _GEN_338;
  wire  _GEN_380 = io_req_bits_addr == 12'h301 ? reg_mip_UTIP : _GEN_339;
  wire  _GEN_381 = io_req_bits_addr == 12'h301 ? reg_mip_MSIP : _GEN_340;
  wire  _GEN_382 = io_req_bits_addr == 12'h301 ? reg_mip_reserved_4 : _GEN_341;
  wire  _GEN_383 = io_req_bits_addr == 12'h301 ? reg_mip_SSIP : _GEN_342;
  wire  _GEN_384 = io_req_bits_addr == 12'h301 ? reg_mip_USIP : _GEN_343;
  wire [63:0] _GEN_385 = io_req_bits_addr == 12'h301 ? reg_pmpcfg0 : _GEN_344;
  wire [63:0] _GEN_386 = io_req_bits_addr == 12'h301 ? reg_pmpcfg1 : _GEN_345;
  wire [63:0] _GEN_387 = io_req_bits_addr == 12'h301 ? reg_pmpcfg2 : _GEN_346;
  wire [63:0] _GEN_388 = io_req_bits_addr == 12'h301 ? reg_pmpcfg3 : _GEN_347;
  wire [63:0] _GEN_389 = io_req_bits_addr == 12'h301 ? reg_pmpaddr0 : _GEN_348;
  wire [63:0] _GEN_390 = io_req_bits_addr == 12'h300 ? _reg_mstatus_T_4 : _GEN_6;
  wire [63:0] _GEN_391 = io_req_bits_addr == 12'h300 ? reg_misa : _GEN_349;
  wire [63:0] _GEN_392 = io_req_bits_addr == 12'h300 ? reg_medeleg : _GEN_350;
  wire [63:0] _GEN_393 = io_req_bits_addr == 12'h300 ? reg_mideleg : _GEN_351;
  wire [63:0] _GEN_394 = io_req_bits_addr == 12'h300 ? reg_mie : _GEN_352;
  wire [61:0] _GEN_395 = io_req_bits_addr == 12'h300 ? reg_mtvec_BASE : _GEN_353;
  wire [1:0] _GEN_396 = io_req_bits_addr == 12'h300 ? reg_mtvec_MODE : _GEN_354;
  wire [63:0] _GEN_397 = io_req_bits_addr == 12'h300 ? reg_mscratch : _GEN_355;
  wire [63:0] _GEN_398 = io_req_bits_addr == 12'h300 ? _GEN_2 : _GEN_356;
  wire  _GEN_399 = io_req_bits_addr == 12'h300 ? _GEN_0 : _GEN_357;
  wire [62:0] _GEN_400 = io_req_bits_addr == 12'h300 ? _GEN_1 : _GEN_358;
  wire [63:0] _GEN_401 = io_req_bits_addr == 12'h300 ? reg_mtval : _GEN_359;
  wire [51:0] _GEN_402 = io_req_bits_addr == 12'h300 ? reg_mip_reserved : _GEN_360;
  wire  _GEN_403 = io_req_bits_addr == 12'h300 ? reg_mip_intr_e_m : _GEN_361;
  wire  _GEN_404 = io_req_bits_addr == 12'h300 ? reg_mip_intr_e_h : _GEN_362;
  wire  _GEN_405 = io_req_bits_addr == 12'h300 ? reg_mip_intr_e_s : _GEN_363;
  wire  _GEN_406 = io_req_bits_addr == 12'h300 ? reg_mip_intr_e_u : _GEN_364;
  wire  _GEN_407 = io_req_bits_addr == 12'h300 ? reg_mip_intr_t_m : _GEN_365;
  wire  _GEN_408 = io_req_bits_addr == 12'h300 ? reg_mip_intr_t_h : _GEN_366;
  wire  _GEN_409 = io_req_bits_addr == 12'h300 ? reg_mip_intr_t_s : _GEN_367;
  wire  _GEN_410 = io_req_bits_addr == 12'h300 ? reg_mip_intr_t_u : _GEN_368;
  wire  _GEN_411 = io_req_bits_addr == 12'h300 ? reg_mip_intr_s_m : _GEN_369;
  wire  _GEN_412 = io_req_bits_addr == 12'h300 ? reg_mip_intr_s_h : _GEN_370;
  wire  _GEN_413 = io_req_bits_addr == 12'h300 ? reg_mip_intr_s_s : _GEN_371;
  wire  _GEN_414 = io_req_bits_addr == 12'h300 ? reg_mip_intr_s_u : _GEN_372;
  wire  _GEN_415 = io_req_bits_addr == 12'h300 ? reg_mip_MEIP : _GEN_373;
  wire  _GEN_416 = io_req_bits_addr == 12'h300 ? reg_mip_reserved_2 : _GEN_374;
  wire  _GEN_417 = io_req_bits_addr == 12'h300 ? reg_mip_SEIP : _GEN_375;
  wire  _GEN_418 = io_req_bits_addr == 12'h300 ? reg_mip_UEIP : _GEN_376;
  wire  _GEN_419 = io_req_bits_addr == 12'h300 ? reg_mip_MTIP : _GEN_377;
  wire  _GEN_420 = io_req_bits_addr == 12'h300 ? reg_mip_reserved_3 : _GEN_378;
  wire  _GEN_421 = io_req_bits_addr == 12'h300 ? reg_mip_STIP : _GEN_379;
  wire  _GEN_422 = io_req_bits_addr == 12'h300 ? reg_mip_UTIP : _GEN_380;
  wire  _GEN_423 = io_req_bits_addr == 12'h300 ? reg_mip_MSIP : _GEN_381;
  wire  _GEN_424 = io_req_bits_addr == 12'h300 ? reg_mip_reserved_4 : _GEN_382;
  wire  _GEN_425 = io_req_bits_addr == 12'h300 ? reg_mip_SSIP : _GEN_383;
  wire  _GEN_426 = io_req_bits_addr == 12'h300 ? reg_mip_USIP : _GEN_384;
  wire [63:0] _GEN_427 = io_req_bits_addr == 12'h300 ? reg_pmpcfg0 : _GEN_385;
  wire [63:0] _GEN_428 = io_req_bits_addr == 12'h300 ? reg_pmpcfg1 : _GEN_386;
  wire [63:0] _GEN_429 = io_req_bits_addr == 12'h300 ? reg_pmpcfg2 : _GEN_387;
  wire [63:0] _GEN_430 = io_req_bits_addr == 12'h300 ? reg_pmpcfg3 : _GEN_388;
  wire [63:0] _GEN_431 = io_req_bits_addr == 12'h300 ? reg_pmpaddr0 : _GEN_389;
  wire [63:0] _GEN_432 = io_req_bits_addr == 12'h144 ? write_data : reg_sip;
  wire [63:0] _GEN_433 = io_req_bits_addr == 12'h144 ? _GEN_6 : _GEN_390;
  wire [63:0] _GEN_434 = io_req_bits_addr == 12'h144 ? reg_misa : _GEN_391;
  wire [63:0] _GEN_435 = io_req_bits_addr == 12'h144 ? reg_medeleg : _GEN_392;
  wire [63:0] _GEN_436 = io_req_bits_addr == 12'h144 ? reg_mideleg : _GEN_393;
  wire [63:0] _GEN_437 = io_req_bits_addr == 12'h144 ? reg_mie : _GEN_394;
  wire [61:0] _GEN_438 = io_req_bits_addr == 12'h144 ? reg_mtvec_BASE : _GEN_395;
  wire [1:0] _GEN_439 = io_req_bits_addr == 12'h144 ? reg_mtvec_MODE : _GEN_396;
  wire [63:0] _GEN_440 = io_req_bits_addr == 12'h144 ? reg_mscratch : _GEN_397;
  wire [63:0] _GEN_441 = io_req_bits_addr == 12'h144 ? _GEN_2 : _GEN_398;
  wire  _GEN_442 = io_req_bits_addr == 12'h144 ? _GEN_0 : _GEN_399;
  wire [62:0] _GEN_443 = io_req_bits_addr == 12'h144 ? _GEN_1 : _GEN_400;
  wire [63:0] _GEN_444 = io_req_bits_addr == 12'h144 ? reg_mtval : _GEN_401;
  wire [51:0] _GEN_445 = io_req_bits_addr == 12'h144 ? reg_mip_reserved : _GEN_402;
  wire  _GEN_446 = io_req_bits_addr == 12'h144 ? reg_mip_intr_e_m : _GEN_403;
  wire  _GEN_447 = io_req_bits_addr == 12'h144 ? reg_mip_intr_e_h : _GEN_404;
  wire  _GEN_448 = io_req_bits_addr == 12'h144 ? reg_mip_intr_e_s : _GEN_405;
  wire  _GEN_449 = io_req_bits_addr == 12'h144 ? reg_mip_intr_e_u : _GEN_406;
  wire  _GEN_450 = io_req_bits_addr == 12'h144 ? reg_mip_intr_t_m : _GEN_407;
  wire  _GEN_451 = io_req_bits_addr == 12'h144 ? reg_mip_intr_t_h : _GEN_408;
  wire  _GEN_452 = io_req_bits_addr == 12'h144 ? reg_mip_intr_t_s : _GEN_409;
  wire  _GEN_453 = io_req_bits_addr == 12'h144 ? reg_mip_intr_t_u : _GEN_410;
  wire  _GEN_454 = io_req_bits_addr == 12'h144 ? reg_mip_intr_s_m : _GEN_411;
  wire  _GEN_455 = io_req_bits_addr == 12'h144 ? reg_mip_intr_s_h : _GEN_412;
  wire  _GEN_456 = io_req_bits_addr == 12'h144 ? reg_mip_intr_s_s : _GEN_413;
  wire  _GEN_457 = io_req_bits_addr == 12'h144 ? reg_mip_intr_s_u : _GEN_414;
  wire  _GEN_458 = io_req_bits_addr == 12'h144 ? reg_mip_MEIP : _GEN_415;
  wire  _GEN_459 = io_req_bits_addr == 12'h144 ? reg_mip_reserved_2 : _GEN_416;
  wire  _GEN_460 = io_req_bits_addr == 12'h144 ? reg_mip_SEIP : _GEN_417;
  wire  _GEN_461 = io_req_bits_addr == 12'h144 ? reg_mip_UEIP : _GEN_418;
  wire  _GEN_462 = io_req_bits_addr == 12'h144 ? reg_mip_MTIP : _GEN_419;
  wire  _GEN_463 = io_req_bits_addr == 12'h144 ? reg_mip_reserved_3 : _GEN_420;
  wire  _GEN_464 = io_req_bits_addr == 12'h144 ? reg_mip_STIP : _GEN_421;
  wire  _GEN_465 = io_req_bits_addr == 12'h144 ? reg_mip_UTIP : _GEN_422;
  wire  _GEN_466 = io_req_bits_addr == 12'h144 ? reg_mip_MSIP : _GEN_423;
  wire  _GEN_467 = io_req_bits_addr == 12'h144 ? reg_mip_reserved_4 : _GEN_424;
  wire  _GEN_468 = io_req_bits_addr == 12'h144 ? reg_mip_SSIP : _GEN_425;
  wire  _GEN_469 = io_req_bits_addr == 12'h144 ? reg_mip_USIP : _GEN_426;
  wire [63:0] _GEN_470 = io_req_bits_addr == 12'h144 ? reg_pmpcfg0 : _GEN_427;
  wire [63:0] _GEN_471 = io_req_bits_addr == 12'h144 ? reg_pmpcfg1 : _GEN_428;
  wire [63:0] _GEN_472 = io_req_bits_addr == 12'h144 ? reg_pmpcfg2 : _GEN_429;
  wire [63:0] _GEN_473 = io_req_bits_addr == 12'h144 ? reg_pmpcfg3 : _GEN_430;
  wire [63:0] _GEN_474 = io_req_bits_addr == 12'h144 ? reg_pmpaddr0 : _GEN_431;
  wire [63:0] _GEN_475 = io_req_bits_addr == 12'h143 ? write_data : reg_stval;
  wire [63:0] _GEN_476 = io_req_bits_addr == 12'h143 ? reg_sip : _GEN_432;
  wire [63:0] _GEN_477 = io_req_bits_addr == 12'h143 ? _GEN_6 : _GEN_433;
  wire [63:0] _GEN_478 = io_req_bits_addr == 12'h143 ? reg_misa : _GEN_434;
  wire [63:0] _GEN_479 = io_req_bits_addr == 12'h143 ? reg_medeleg : _GEN_435;
  wire [63:0] _GEN_480 = io_req_bits_addr == 12'h143 ? reg_mideleg : _GEN_436;
  wire [63:0] _GEN_481 = io_req_bits_addr == 12'h143 ? reg_mie : _GEN_437;
  wire [61:0] _GEN_482 = io_req_bits_addr == 12'h143 ? reg_mtvec_BASE : _GEN_438;
  wire [1:0] _GEN_483 = io_req_bits_addr == 12'h143 ? reg_mtvec_MODE : _GEN_439;
  wire [63:0] _GEN_484 = io_req_bits_addr == 12'h143 ? reg_mscratch : _GEN_440;
  wire [63:0] _GEN_485 = io_req_bits_addr == 12'h143 ? _GEN_2 : _GEN_441;
  wire  _GEN_486 = io_req_bits_addr == 12'h143 ? _GEN_0 : _GEN_442;
  wire [62:0] _GEN_487 = io_req_bits_addr == 12'h143 ? _GEN_1 : _GEN_443;
  wire [63:0] _GEN_488 = io_req_bits_addr == 12'h143 ? reg_mtval : _GEN_444;
  wire [51:0] _GEN_489 = io_req_bits_addr == 12'h143 ? reg_mip_reserved : _GEN_445;
  wire  _GEN_490 = io_req_bits_addr == 12'h143 ? reg_mip_intr_e_m : _GEN_446;
  wire  _GEN_491 = io_req_bits_addr == 12'h143 ? reg_mip_intr_e_h : _GEN_447;
  wire  _GEN_492 = io_req_bits_addr == 12'h143 ? reg_mip_intr_e_s : _GEN_448;
  wire  _GEN_493 = io_req_bits_addr == 12'h143 ? reg_mip_intr_e_u : _GEN_449;
  wire  _GEN_494 = io_req_bits_addr == 12'h143 ? reg_mip_intr_t_m : _GEN_450;
  wire  _GEN_495 = io_req_bits_addr == 12'h143 ? reg_mip_intr_t_h : _GEN_451;
  wire  _GEN_496 = io_req_bits_addr == 12'h143 ? reg_mip_intr_t_s : _GEN_452;
  wire  _GEN_497 = io_req_bits_addr == 12'h143 ? reg_mip_intr_t_u : _GEN_453;
  wire  _GEN_498 = io_req_bits_addr == 12'h143 ? reg_mip_intr_s_m : _GEN_454;
  wire  _GEN_499 = io_req_bits_addr == 12'h143 ? reg_mip_intr_s_h : _GEN_455;
  wire  _GEN_500 = io_req_bits_addr == 12'h143 ? reg_mip_intr_s_s : _GEN_456;
  wire  _GEN_501 = io_req_bits_addr == 12'h143 ? reg_mip_intr_s_u : _GEN_457;
  wire  _GEN_502 = io_req_bits_addr == 12'h143 ? reg_mip_MEIP : _GEN_458;
  wire  _GEN_503 = io_req_bits_addr == 12'h143 ? reg_mip_reserved_2 : _GEN_459;
  wire  _GEN_504 = io_req_bits_addr == 12'h143 ? reg_mip_SEIP : _GEN_460;
  wire  _GEN_505 = io_req_bits_addr == 12'h143 ? reg_mip_UEIP : _GEN_461;
  wire  _GEN_506 = io_req_bits_addr == 12'h143 ? reg_mip_MTIP : _GEN_462;
  wire  _GEN_507 = io_req_bits_addr == 12'h143 ? reg_mip_reserved_3 : _GEN_463;
  wire  _GEN_508 = io_req_bits_addr == 12'h143 ? reg_mip_STIP : _GEN_464;
  wire  _GEN_509 = io_req_bits_addr == 12'h143 ? reg_mip_UTIP : _GEN_465;
  wire  _GEN_510 = io_req_bits_addr == 12'h143 ? reg_mip_MSIP : _GEN_466;
  wire  _GEN_511 = io_req_bits_addr == 12'h143 ? reg_mip_reserved_4 : _GEN_467;
  wire  _GEN_512 = io_req_bits_addr == 12'h143 ? reg_mip_SSIP : _GEN_468;
  wire  _GEN_513 = io_req_bits_addr == 12'h143 ? reg_mip_USIP : _GEN_469;
  wire [63:0] _GEN_514 = io_req_bits_addr == 12'h143 ? reg_pmpcfg0 : _GEN_470;
  wire [63:0] _GEN_515 = io_req_bits_addr == 12'h143 ? reg_pmpcfg1 : _GEN_471;
  wire [63:0] _GEN_516 = io_req_bits_addr == 12'h143 ? reg_pmpcfg2 : _GEN_472;
  wire [63:0] _GEN_517 = io_req_bits_addr == 12'h143 ? reg_pmpcfg3 : _GEN_473;
  wire [63:0] _GEN_518 = io_req_bits_addr == 12'h143 ? reg_pmpaddr0 : _GEN_474;
  wire [63:0] _GEN_519 = io_req_bits_addr == 12'h142 ? write_data : reg_scause;
  wire [63:0] _GEN_520 = io_req_bits_addr == 12'h142 ? reg_stval : _GEN_475;
  wire [63:0] _GEN_521 = io_req_bits_addr == 12'h142 ? reg_sip : _GEN_476;
  wire [63:0] _GEN_522 = io_req_bits_addr == 12'h142 ? _GEN_6 : _GEN_477;
  wire [63:0] _GEN_523 = io_req_bits_addr == 12'h142 ? reg_misa : _GEN_478;
  wire [63:0] _GEN_524 = io_req_bits_addr == 12'h142 ? reg_medeleg : _GEN_479;
  wire [63:0] _GEN_525 = io_req_bits_addr == 12'h142 ? reg_mideleg : _GEN_480;
  wire [63:0] _GEN_526 = io_req_bits_addr == 12'h142 ? reg_mie : _GEN_481;
  wire [61:0] _GEN_527 = io_req_bits_addr == 12'h142 ? reg_mtvec_BASE : _GEN_482;
  wire [1:0] _GEN_528 = io_req_bits_addr == 12'h142 ? reg_mtvec_MODE : _GEN_483;
  wire [63:0] _GEN_529 = io_req_bits_addr == 12'h142 ? reg_mscratch : _GEN_484;
  wire [63:0] _GEN_530 = io_req_bits_addr == 12'h142 ? _GEN_2 : _GEN_485;
  wire  _GEN_531 = io_req_bits_addr == 12'h142 ? _GEN_0 : _GEN_486;
  wire [62:0] _GEN_532 = io_req_bits_addr == 12'h142 ? _GEN_1 : _GEN_487;
  wire [63:0] _GEN_533 = io_req_bits_addr == 12'h142 ? reg_mtval : _GEN_488;
  wire [51:0] _GEN_534 = io_req_bits_addr == 12'h142 ? reg_mip_reserved : _GEN_489;
  wire  _GEN_535 = io_req_bits_addr == 12'h142 ? reg_mip_intr_e_m : _GEN_490;
  wire  _GEN_536 = io_req_bits_addr == 12'h142 ? reg_mip_intr_e_h : _GEN_491;
  wire  _GEN_537 = io_req_bits_addr == 12'h142 ? reg_mip_intr_e_s : _GEN_492;
  wire  _GEN_538 = io_req_bits_addr == 12'h142 ? reg_mip_intr_e_u : _GEN_493;
  wire  _GEN_539 = io_req_bits_addr == 12'h142 ? reg_mip_intr_t_m : _GEN_494;
  wire  _GEN_540 = io_req_bits_addr == 12'h142 ? reg_mip_intr_t_h : _GEN_495;
  wire  _GEN_541 = io_req_bits_addr == 12'h142 ? reg_mip_intr_t_s : _GEN_496;
  wire  _GEN_542 = io_req_bits_addr == 12'h142 ? reg_mip_intr_t_u : _GEN_497;
  wire  _GEN_543 = io_req_bits_addr == 12'h142 ? reg_mip_intr_s_m : _GEN_498;
  wire  _GEN_544 = io_req_bits_addr == 12'h142 ? reg_mip_intr_s_h : _GEN_499;
  wire  _GEN_545 = io_req_bits_addr == 12'h142 ? reg_mip_intr_s_s : _GEN_500;
  wire  _GEN_546 = io_req_bits_addr == 12'h142 ? reg_mip_intr_s_u : _GEN_501;
  wire  _GEN_547 = io_req_bits_addr == 12'h142 ? reg_mip_MEIP : _GEN_502;
  wire  _GEN_548 = io_req_bits_addr == 12'h142 ? reg_mip_reserved_2 : _GEN_503;
  wire  _GEN_549 = io_req_bits_addr == 12'h142 ? reg_mip_SEIP : _GEN_504;
  wire  _GEN_550 = io_req_bits_addr == 12'h142 ? reg_mip_UEIP : _GEN_505;
  wire  _GEN_551 = io_req_bits_addr == 12'h142 ? reg_mip_MTIP : _GEN_506;
  wire  _GEN_552 = io_req_bits_addr == 12'h142 ? reg_mip_reserved_3 : _GEN_507;
  wire  _GEN_553 = io_req_bits_addr == 12'h142 ? reg_mip_STIP : _GEN_508;
  wire  _GEN_554 = io_req_bits_addr == 12'h142 ? reg_mip_UTIP : _GEN_509;
  wire  _GEN_555 = io_req_bits_addr == 12'h142 ? reg_mip_MSIP : _GEN_510;
  wire  _GEN_556 = io_req_bits_addr == 12'h142 ? reg_mip_reserved_4 : _GEN_511;
  wire  _GEN_557 = io_req_bits_addr == 12'h142 ? reg_mip_SSIP : _GEN_512;
  wire  _GEN_558 = io_req_bits_addr == 12'h142 ? reg_mip_USIP : _GEN_513;
  wire [63:0] _GEN_559 = io_req_bits_addr == 12'h142 ? reg_pmpcfg0 : _GEN_514;
  wire [63:0] _GEN_560 = io_req_bits_addr == 12'h142 ? reg_pmpcfg1 : _GEN_515;
  wire [63:0] _GEN_561 = io_req_bits_addr == 12'h142 ? reg_pmpcfg2 : _GEN_516;
  wire [63:0] _GEN_562 = io_req_bits_addr == 12'h142 ? reg_pmpcfg3 : _GEN_517;
  wire [63:0] _GEN_563 = io_req_bits_addr == 12'h142 ? reg_pmpaddr0 : _GEN_518;
  wire [63:0] _GEN_564 = io_req_bits_addr == 12'h140 ? write_data : reg_sscratch;
  wire [63:0] _GEN_565 = io_req_bits_addr == 12'h140 ? reg_scause : _GEN_519;
  wire [63:0] _GEN_566 = io_req_bits_addr == 12'h140 ? reg_stval : _GEN_520;
  wire [63:0] _GEN_567 = io_req_bits_addr == 12'h140 ? reg_sip : _GEN_521;
  wire [63:0] _GEN_568 = io_req_bits_addr == 12'h140 ? _GEN_6 : _GEN_522;
  wire [63:0] _GEN_569 = io_req_bits_addr == 12'h140 ? reg_misa : _GEN_523;
  wire [63:0] _GEN_570 = io_req_bits_addr == 12'h140 ? reg_medeleg : _GEN_524;
  wire [63:0] _GEN_571 = io_req_bits_addr == 12'h140 ? reg_mideleg : _GEN_525;
  wire [63:0] _GEN_572 = io_req_bits_addr == 12'h140 ? reg_mie : _GEN_526;
  wire [61:0] _GEN_573 = io_req_bits_addr == 12'h140 ? reg_mtvec_BASE : _GEN_527;
  wire [1:0] _GEN_574 = io_req_bits_addr == 12'h140 ? reg_mtvec_MODE : _GEN_528;
  wire [63:0] _GEN_575 = io_req_bits_addr == 12'h140 ? reg_mscratch : _GEN_529;
  wire [63:0] _GEN_576 = io_req_bits_addr == 12'h140 ? _GEN_2 : _GEN_530;
  wire  _GEN_577 = io_req_bits_addr == 12'h140 ? _GEN_0 : _GEN_531;
  wire [62:0] _GEN_578 = io_req_bits_addr == 12'h140 ? _GEN_1 : _GEN_532;
  wire [63:0] _GEN_579 = io_req_bits_addr == 12'h140 ? reg_mtval : _GEN_533;
  wire [51:0] _GEN_580 = io_req_bits_addr == 12'h140 ? reg_mip_reserved : _GEN_534;
  wire  _GEN_581 = io_req_bits_addr == 12'h140 ? reg_mip_intr_e_m : _GEN_535;
  wire  _GEN_582 = io_req_bits_addr == 12'h140 ? reg_mip_intr_e_h : _GEN_536;
  wire  _GEN_583 = io_req_bits_addr == 12'h140 ? reg_mip_intr_e_s : _GEN_537;
  wire  _GEN_584 = io_req_bits_addr == 12'h140 ? reg_mip_intr_e_u : _GEN_538;
  wire  _GEN_585 = io_req_bits_addr == 12'h140 ? reg_mip_intr_t_m : _GEN_539;
  wire  _GEN_586 = io_req_bits_addr == 12'h140 ? reg_mip_intr_t_h : _GEN_540;
  wire  _GEN_587 = io_req_bits_addr == 12'h140 ? reg_mip_intr_t_s : _GEN_541;
  wire  _GEN_588 = io_req_bits_addr == 12'h140 ? reg_mip_intr_t_u : _GEN_542;
  wire  _GEN_589 = io_req_bits_addr == 12'h140 ? reg_mip_intr_s_m : _GEN_543;
  wire  _GEN_590 = io_req_bits_addr == 12'h140 ? reg_mip_intr_s_h : _GEN_544;
  wire  _GEN_591 = io_req_bits_addr == 12'h140 ? reg_mip_intr_s_s : _GEN_545;
  wire  _GEN_592 = io_req_bits_addr == 12'h140 ? reg_mip_intr_s_u : _GEN_546;
  wire  _GEN_593 = io_req_bits_addr == 12'h140 ? reg_mip_MEIP : _GEN_547;
  wire  _GEN_594 = io_req_bits_addr == 12'h140 ? reg_mip_reserved_2 : _GEN_548;
  wire  _GEN_595 = io_req_bits_addr == 12'h140 ? reg_mip_SEIP : _GEN_549;
  wire  _GEN_596 = io_req_bits_addr == 12'h140 ? reg_mip_UEIP : _GEN_550;
  wire  _GEN_597 = io_req_bits_addr == 12'h140 ? reg_mip_MTIP : _GEN_551;
  wire  _GEN_598 = io_req_bits_addr == 12'h140 ? reg_mip_reserved_3 : _GEN_552;
  wire  _GEN_599 = io_req_bits_addr == 12'h140 ? reg_mip_STIP : _GEN_553;
  wire  _GEN_600 = io_req_bits_addr == 12'h140 ? reg_mip_UTIP : _GEN_554;
  wire  _GEN_601 = io_req_bits_addr == 12'h140 ? reg_mip_MSIP : _GEN_555;
  wire  _GEN_602 = io_req_bits_addr == 12'h140 ? reg_mip_reserved_4 : _GEN_556;
  wire  _GEN_603 = io_req_bits_addr == 12'h140 ? reg_mip_SSIP : _GEN_557;
  wire  _GEN_604 = io_req_bits_addr == 12'h140 ? reg_mip_USIP : _GEN_558;
  wire [63:0] _GEN_605 = io_req_bits_addr == 12'h140 ? reg_pmpcfg0 : _GEN_559;
  wire [63:0] _GEN_606 = io_req_bits_addr == 12'h140 ? reg_pmpcfg1 : _GEN_560;
  wire [63:0] _GEN_607 = io_req_bits_addr == 12'h140 ? reg_pmpcfg2 : _GEN_561;
  wire [63:0] _GEN_608 = io_req_bits_addr == 12'h140 ? reg_pmpcfg3 : _GEN_562;
  wire [63:0] _GEN_609 = io_req_bits_addr == 12'h140 ? reg_pmpaddr0 : _GEN_563;
  wire [63:0] _GEN_610 = io_req_bits_addr == 12'h106 ? write_data : reg_scounteren;
  wire [63:0] _GEN_611 = io_req_bits_addr == 12'h106 ? reg_sscratch : _GEN_564;
  wire [63:0] _GEN_612 = io_req_bits_addr == 12'h106 ? reg_scause : _GEN_565;
  wire [63:0] _GEN_613 = io_req_bits_addr == 12'h106 ? reg_stval : _GEN_566;
  wire [63:0] _GEN_614 = io_req_bits_addr == 12'h106 ? reg_sip : _GEN_567;
  wire [63:0] _GEN_615 = io_req_bits_addr == 12'h106 ? _GEN_6 : _GEN_568;
  wire [63:0] _GEN_616 = io_req_bits_addr == 12'h106 ? reg_misa : _GEN_569;
  wire [63:0] _GEN_617 = io_req_bits_addr == 12'h106 ? reg_medeleg : _GEN_570;
  wire [63:0] _GEN_618 = io_req_bits_addr == 12'h106 ? reg_mideleg : _GEN_571;
  wire [63:0] _GEN_619 = io_req_bits_addr == 12'h106 ? reg_mie : _GEN_572;
  wire [61:0] _GEN_620 = io_req_bits_addr == 12'h106 ? reg_mtvec_BASE : _GEN_573;
  wire [1:0] _GEN_621 = io_req_bits_addr == 12'h106 ? reg_mtvec_MODE : _GEN_574;
  wire [63:0] _GEN_622 = io_req_bits_addr == 12'h106 ? reg_mscratch : _GEN_575;
  wire [63:0] _GEN_623 = io_req_bits_addr == 12'h106 ? _GEN_2 : _GEN_576;
  wire  _GEN_624 = io_req_bits_addr == 12'h106 ? _GEN_0 : _GEN_577;
  wire [62:0] _GEN_625 = io_req_bits_addr == 12'h106 ? _GEN_1 : _GEN_578;
  wire [63:0] _GEN_626 = io_req_bits_addr == 12'h106 ? reg_mtval : _GEN_579;
  wire [51:0] _GEN_627 = io_req_bits_addr == 12'h106 ? reg_mip_reserved : _GEN_580;
  wire  _GEN_628 = io_req_bits_addr == 12'h106 ? reg_mip_intr_e_m : _GEN_581;
  wire  _GEN_629 = io_req_bits_addr == 12'h106 ? reg_mip_intr_e_h : _GEN_582;
  wire  _GEN_630 = io_req_bits_addr == 12'h106 ? reg_mip_intr_e_s : _GEN_583;
  wire  _GEN_631 = io_req_bits_addr == 12'h106 ? reg_mip_intr_e_u : _GEN_584;
  wire  _GEN_632 = io_req_bits_addr == 12'h106 ? reg_mip_intr_t_m : _GEN_585;
  wire  _GEN_633 = io_req_bits_addr == 12'h106 ? reg_mip_intr_t_h : _GEN_586;
  wire  _GEN_634 = io_req_bits_addr == 12'h106 ? reg_mip_intr_t_s : _GEN_587;
  wire  _GEN_635 = io_req_bits_addr == 12'h106 ? reg_mip_intr_t_u : _GEN_588;
  wire  _GEN_636 = io_req_bits_addr == 12'h106 ? reg_mip_intr_s_m : _GEN_589;
  wire  _GEN_637 = io_req_bits_addr == 12'h106 ? reg_mip_intr_s_h : _GEN_590;
  wire  _GEN_638 = io_req_bits_addr == 12'h106 ? reg_mip_intr_s_s : _GEN_591;
  wire  _GEN_639 = io_req_bits_addr == 12'h106 ? reg_mip_intr_s_u : _GEN_592;
  wire  _GEN_640 = io_req_bits_addr == 12'h106 ? reg_mip_MEIP : _GEN_593;
  wire  _GEN_641 = io_req_bits_addr == 12'h106 ? reg_mip_reserved_2 : _GEN_594;
  wire  _GEN_642 = io_req_bits_addr == 12'h106 ? reg_mip_SEIP : _GEN_595;
  wire  _GEN_643 = io_req_bits_addr == 12'h106 ? reg_mip_UEIP : _GEN_596;
  wire  _GEN_644 = io_req_bits_addr == 12'h106 ? reg_mip_MTIP : _GEN_597;
  wire  _GEN_645 = io_req_bits_addr == 12'h106 ? reg_mip_reserved_3 : _GEN_598;
  wire  _GEN_646 = io_req_bits_addr == 12'h106 ? reg_mip_STIP : _GEN_599;
  wire  _GEN_647 = io_req_bits_addr == 12'h106 ? reg_mip_UTIP : _GEN_600;
  wire  _GEN_648 = io_req_bits_addr == 12'h106 ? reg_mip_MSIP : _GEN_601;
  wire  _GEN_649 = io_req_bits_addr == 12'h106 ? reg_mip_reserved_4 : _GEN_602;
  wire  _GEN_650 = io_req_bits_addr == 12'h106 ? reg_mip_SSIP : _GEN_603;
  wire  _GEN_651 = io_req_bits_addr == 12'h106 ? reg_mip_USIP : _GEN_604;
  wire [63:0] _GEN_652 = io_req_bits_addr == 12'h106 ? reg_pmpcfg0 : _GEN_605;
  wire [63:0] _GEN_653 = io_req_bits_addr == 12'h106 ? reg_pmpcfg1 : _GEN_606;
  wire [63:0] _GEN_654 = io_req_bits_addr == 12'h106 ? reg_pmpcfg2 : _GEN_607;
  wire [63:0] _GEN_655 = io_req_bits_addr == 12'h106 ? reg_pmpcfg3 : _GEN_608;
  wire [63:0] _GEN_656 = io_req_bits_addr == 12'h106 ? reg_pmpaddr0 : _GEN_609;
  wire [63:0] _GEN_657 = io_req_bits_addr == 12'h105 ? write_data : reg_stvec;
  wire [63:0] _GEN_658 = io_req_bits_addr == 12'h105 ? reg_scounteren : _GEN_610;
  wire [63:0] _GEN_659 = io_req_bits_addr == 12'h105 ? reg_sscratch : _GEN_611;
  wire [63:0] _GEN_660 = io_req_bits_addr == 12'h105 ? reg_scause : _GEN_612;
  wire [63:0] _GEN_661 = io_req_bits_addr == 12'h105 ? reg_stval : _GEN_613;
  wire [63:0] _GEN_662 = io_req_bits_addr == 12'h105 ? reg_sip : _GEN_614;
  wire [63:0] _GEN_663 = io_req_bits_addr == 12'h105 ? _GEN_6 : _GEN_615;
  wire [63:0] _GEN_664 = io_req_bits_addr == 12'h105 ? reg_misa : _GEN_616;
  wire [63:0] _GEN_665 = io_req_bits_addr == 12'h105 ? reg_medeleg : _GEN_617;
  wire [63:0] _GEN_666 = io_req_bits_addr == 12'h105 ? reg_mideleg : _GEN_618;
  wire [63:0] _GEN_667 = io_req_bits_addr == 12'h105 ? reg_mie : _GEN_619;
  wire [61:0] _GEN_668 = io_req_bits_addr == 12'h105 ? reg_mtvec_BASE : _GEN_620;
  wire [1:0] _GEN_669 = io_req_bits_addr == 12'h105 ? reg_mtvec_MODE : _GEN_621;
  wire [63:0] _GEN_670 = io_req_bits_addr == 12'h105 ? reg_mscratch : _GEN_622;
  wire [63:0] _GEN_671 = io_req_bits_addr == 12'h105 ? _GEN_2 : _GEN_623;
  wire  _GEN_672 = io_req_bits_addr == 12'h105 ? _GEN_0 : _GEN_624;
  wire [62:0] _GEN_673 = io_req_bits_addr == 12'h105 ? _GEN_1 : _GEN_625;
  wire [63:0] _GEN_674 = io_req_bits_addr == 12'h105 ? reg_mtval : _GEN_626;
  wire [51:0] _GEN_675 = io_req_bits_addr == 12'h105 ? reg_mip_reserved : _GEN_627;
  wire  _GEN_676 = io_req_bits_addr == 12'h105 ? reg_mip_intr_e_m : _GEN_628;
  wire  _GEN_677 = io_req_bits_addr == 12'h105 ? reg_mip_intr_e_h : _GEN_629;
  wire  _GEN_678 = io_req_bits_addr == 12'h105 ? reg_mip_intr_e_s : _GEN_630;
  wire  _GEN_679 = io_req_bits_addr == 12'h105 ? reg_mip_intr_e_u : _GEN_631;
  wire  _GEN_680 = io_req_bits_addr == 12'h105 ? reg_mip_intr_t_m : _GEN_632;
  wire  _GEN_681 = io_req_bits_addr == 12'h105 ? reg_mip_intr_t_h : _GEN_633;
  wire  _GEN_682 = io_req_bits_addr == 12'h105 ? reg_mip_intr_t_s : _GEN_634;
  wire  _GEN_683 = io_req_bits_addr == 12'h105 ? reg_mip_intr_t_u : _GEN_635;
  wire  _GEN_684 = io_req_bits_addr == 12'h105 ? reg_mip_intr_s_m : _GEN_636;
  wire  _GEN_685 = io_req_bits_addr == 12'h105 ? reg_mip_intr_s_h : _GEN_637;
  wire  _GEN_686 = io_req_bits_addr == 12'h105 ? reg_mip_intr_s_s : _GEN_638;
  wire  _GEN_687 = io_req_bits_addr == 12'h105 ? reg_mip_intr_s_u : _GEN_639;
  wire  _GEN_688 = io_req_bits_addr == 12'h105 ? reg_mip_MEIP : _GEN_640;
  wire  _GEN_689 = io_req_bits_addr == 12'h105 ? reg_mip_reserved_2 : _GEN_641;
  wire  _GEN_690 = io_req_bits_addr == 12'h105 ? reg_mip_SEIP : _GEN_642;
  wire  _GEN_691 = io_req_bits_addr == 12'h105 ? reg_mip_UEIP : _GEN_643;
  wire  _GEN_692 = io_req_bits_addr == 12'h105 ? reg_mip_MTIP : _GEN_644;
  wire  _GEN_693 = io_req_bits_addr == 12'h105 ? reg_mip_reserved_3 : _GEN_645;
  wire  _GEN_694 = io_req_bits_addr == 12'h105 ? reg_mip_STIP : _GEN_646;
  wire  _GEN_695 = io_req_bits_addr == 12'h105 ? reg_mip_UTIP : _GEN_647;
  wire  _GEN_696 = io_req_bits_addr == 12'h105 ? reg_mip_MSIP : _GEN_648;
  wire  _GEN_697 = io_req_bits_addr == 12'h105 ? reg_mip_reserved_4 : _GEN_649;
  wire  _GEN_698 = io_req_bits_addr == 12'h105 ? reg_mip_SSIP : _GEN_650;
  wire  _GEN_699 = io_req_bits_addr == 12'h105 ? reg_mip_USIP : _GEN_651;
  wire [63:0] _GEN_700 = io_req_bits_addr == 12'h105 ? reg_pmpcfg0 : _GEN_652;
  wire [63:0] _GEN_701 = io_req_bits_addr == 12'h105 ? reg_pmpcfg1 : _GEN_653;
  wire [63:0] _GEN_702 = io_req_bits_addr == 12'h105 ? reg_pmpcfg2 : _GEN_654;
  wire [63:0] _GEN_703 = io_req_bits_addr == 12'h105 ? reg_pmpcfg3 : _GEN_655;
  wire [63:0] _GEN_704 = io_req_bits_addr == 12'h105 ? reg_pmpaddr0 : _GEN_656;
  wire [63:0] _GEN_705 = io_req_bits_addr == 12'h104 ? write_data : reg_sie;
  wire [63:0] _GEN_706 = io_req_bits_addr == 12'h104 ? reg_stvec : _GEN_657;
  wire [63:0] _GEN_707 = io_req_bits_addr == 12'h104 ? reg_scounteren : _GEN_658;
  wire [63:0] _GEN_708 = io_req_bits_addr == 12'h104 ? reg_sscratch : _GEN_659;
  wire [63:0] _GEN_709 = io_req_bits_addr == 12'h104 ? reg_scause : _GEN_660;
  wire [63:0] _GEN_710 = io_req_bits_addr == 12'h104 ? reg_stval : _GEN_661;
  wire [63:0] _GEN_711 = io_req_bits_addr == 12'h104 ? reg_sip : _GEN_662;
  wire [63:0] _GEN_712 = io_req_bits_addr == 12'h104 ? _GEN_6 : _GEN_663;
  wire [63:0] _GEN_713 = io_req_bits_addr == 12'h104 ? reg_misa : _GEN_664;
  wire [63:0] _GEN_714 = io_req_bits_addr == 12'h104 ? reg_medeleg : _GEN_665;
  wire [63:0] _GEN_715 = io_req_bits_addr == 12'h104 ? reg_mideleg : _GEN_666;
  wire [63:0] _GEN_716 = io_req_bits_addr == 12'h104 ? reg_mie : _GEN_667;
  wire [61:0] _GEN_717 = io_req_bits_addr == 12'h104 ? reg_mtvec_BASE : _GEN_668;
  wire [1:0] _GEN_718 = io_req_bits_addr == 12'h104 ? reg_mtvec_MODE : _GEN_669;
  wire [63:0] _GEN_719 = io_req_bits_addr == 12'h104 ? reg_mscratch : _GEN_670;
  wire [63:0] _GEN_720 = io_req_bits_addr == 12'h104 ? _GEN_2 : _GEN_671;
  wire  _GEN_721 = io_req_bits_addr == 12'h104 ? _GEN_0 : _GEN_672;
  wire [62:0] _GEN_722 = io_req_bits_addr == 12'h104 ? _GEN_1 : _GEN_673;
  wire [63:0] _GEN_723 = io_req_bits_addr == 12'h104 ? reg_mtval : _GEN_674;
  wire [51:0] _GEN_724 = io_req_bits_addr == 12'h104 ? reg_mip_reserved : _GEN_675;
  wire  _GEN_725 = io_req_bits_addr == 12'h104 ? reg_mip_intr_e_m : _GEN_676;
  wire  _GEN_726 = io_req_bits_addr == 12'h104 ? reg_mip_intr_e_h : _GEN_677;
  wire  _GEN_727 = io_req_bits_addr == 12'h104 ? reg_mip_intr_e_s : _GEN_678;
  wire  _GEN_728 = io_req_bits_addr == 12'h104 ? reg_mip_intr_e_u : _GEN_679;
  wire  _GEN_729 = io_req_bits_addr == 12'h104 ? reg_mip_intr_t_m : _GEN_680;
  wire  _GEN_730 = io_req_bits_addr == 12'h104 ? reg_mip_intr_t_h : _GEN_681;
  wire  _GEN_731 = io_req_bits_addr == 12'h104 ? reg_mip_intr_t_s : _GEN_682;
  wire  _GEN_732 = io_req_bits_addr == 12'h104 ? reg_mip_intr_t_u : _GEN_683;
  wire  _GEN_733 = io_req_bits_addr == 12'h104 ? reg_mip_intr_s_m : _GEN_684;
  wire  _GEN_734 = io_req_bits_addr == 12'h104 ? reg_mip_intr_s_h : _GEN_685;
  wire  _GEN_735 = io_req_bits_addr == 12'h104 ? reg_mip_intr_s_s : _GEN_686;
  wire  _GEN_736 = io_req_bits_addr == 12'h104 ? reg_mip_intr_s_u : _GEN_687;
  wire  _GEN_737 = io_req_bits_addr == 12'h104 ? reg_mip_MEIP : _GEN_688;
  wire  _GEN_738 = io_req_bits_addr == 12'h104 ? reg_mip_reserved_2 : _GEN_689;
  wire  _GEN_739 = io_req_bits_addr == 12'h104 ? reg_mip_SEIP : _GEN_690;
  wire  _GEN_740 = io_req_bits_addr == 12'h104 ? reg_mip_UEIP : _GEN_691;
  wire  _GEN_741 = io_req_bits_addr == 12'h104 ? reg_mip_MTIP : _GEN_692;
  wire  _GEN_742 = io_req_bits_addr == 12'h104 ? reg_mip_reserved_3 : _GEN_693;
  wire  _GEN_743 = io_req_bits_addr == 12'h104 ? reg_mip_STIP : _GEN_694;
  wire  _GEN_744 = io_req_bits_addr == 12'h104 ? reg_mip_UTIP : _GEN_695;
  wire  _GEN_745 = io_req_bits_addr == 12'h104 ? reg_mip_MSIP : _GEN_696;
  wire  _GEN_746 = io_req_bits_addr == 12'h104 ? reg_mip_reserved_4 : _GEN_697;
  wire  _GEN_747 = io_req_bits_addr == 12'h104 ? reg_mip_SSIP : _GEN_698;
  wire  _GEN_748 = io_req_bits_addr == 12'h104 ? reg_mip_USIP : _GEN_699;
  wire [63:0] _GEN_749 = io_req_bits_addr == 12'h104 ? reg_pmpcfg0 : _GEN_700;
  wire [63:0] _GEN_750 = io_req_bits_addr == 12'h104 ? reg_pmpcfg1 : _GEN_701;
  wire [63:0] _GEN_751 = io_req_bits_addr == 12'h104 ? reg_pmpcfg2 : _GEN_702;
  wire [63:0] _GEN_752 = io_req_bits_addr == 12'h104 ? reg_pmpcfg3 : _GEN_703;
  wire [63:0] _GEN_753 = io_req_bits_addr == 12'h104 ? reg_pmpaddr0 : _GEN_704;
  wire [63:0] _GEN_754 = io_req_bits_addr == 12'h103 ? write_data : reg_sideleg;
  wire [63:0] _GEN_755 = io_req_bits_addr == 12'h103 ? reg_sie : _GEN_705;
  wire [63:0] _GEN_756 = io_req_bits_addr == 12'h103 ? reg_stvec : _GEN_706;
  wire [63:0] _GEN_757 = io_req_bits_addr == 12'h103 ? reg_scounteren : _GEN_707;
  wire [63:0] _GEN_758 = io_req_bits_addr == 12'h103 ? reg_sscratch : _GEN_708;
  wire [63:0] _GEN_759 = io_req_bits_addr == 12'h103 ? reg_scause : _GEN_709;
  wire [63:0] _GEN_760 = io_req_bits_addr == 12'h103 ? reg_stval : _GEN_710;
  wire [63:0] _GEN_761 = io_req_bits_addr == 12'h103 ? reg_sip : _GEN_711;
  wire [63:0] _GEN_762 = io_req_bits_addr == 12'h103 ? _GEN_6 : _GEN_712;
  wire [63:0] _GEN_763 = io_req_bits_addr == 12'h103 ? reg_misa : _GEN_713;
  wire [63:0] _GEN_764 = io_req_bits_addr == 12'h103 ? reg_medeleg : _GEN_714;
  wire [63:0] _GEN_765 = io_req_bits_addr == 12'h103 ? reg_mideleg : _GEN_715;
  wire [63:0] _GEN_766 = io_req_bits_addr == 12'h103 ? reg_mie : _GEN_716;
  wire [61:0] _GEN_767 = io_req_bits_addr == 12'h103 ? reg_mtvec_BASE : _GEN_717;
  wire [1:0] _GEN_768 = io_req_bits_addr == 12'h103 ? reg_mtvec_MODE : _GEN_718;
  wire [63:0] _GEN_769 = io_req_bits_addr == 12'h103 ? reg_mscratch : _GEN_719;
  wire [63:0] _GEN_770 = io_req_bits_addr == 12'h103 ? _GEN_2 : _GEN_720;
  wire  _GEN_771 = io_req_bits_addr == 12'h103 ? _GEN_0 : _GEN_721;
  wire [62:0] _GEN_772 = io_req_bits_addr == 12'h103 ? _GEN_1 : _GEN_722;
  wire [63:0] _GEN_773 = io_req_bits_addr == 12'h103 ? reg_mtval : _GEN_723;
  wire [51:0] _GEN_774 = io_req_bits_addr == 12'h103 ? reg_mip_reserved : _GEN_724;
  wire  _GEN_775 = io_req_bits_addr == 12'h103 ? reg_mip_intr_e_m : _GEN_725;
  wire  _GEN_776 = io_req_bits_addr == 12'h103 ? reg_mip_intr_e_h : _GEN_726;
  wire  _GEN_777 = io_req_bits_addr == 12'h103 ? reg_mip_intr_e_s : _GEN_727;
  wire  _GEN_778 = io_req_bits_addr == 12'h103 ? reg_mip_intr_e_u : _GEN_728;
  wire  _GEN_779 = io_req_bits_addr == 12'h103 ? reg_mip_intr_t_m : _GEN_729;
  wire  _GEN_780 = io_req_bits_addr == 12'h103 ? reg_mip_intr_t_h : _GEN_730;
  wire  _GEN_781 = io_req_bits_addr == 12'h103 ? reg_mip_intr_t_s : _GEN_731;
  wire  _GEN_782 = io_req_bits_addr == 12'h103 ? reg_mip_intr_t_u : _GEN_732;
  wire  _GEN_783 = io_req_bits_addr == 12'h103 ? reg_mip_intr_s_m : _GEN_733;
  wire  _GEN_784 = io_req_bits_addr == 12'h103 ? reg_mip_intr_s_h : _GEN_734;
  wire  _GEN_785 = io_req_bits_addr == 12'h103 ? reg_mip_intr_s_s : _GEN_735;
  wire  _GEN_786 = io_req_bits_addr == 12'h103 ? reg_mip_intr_s_u : _GEN_736;
  wire  _GEN_787 = io_req_bits_addr == 12'h103 ? reg_mip_MEIP : _GEN_737;
  wire  _GEN_788 = io_req_bits_addr == 12'h103 ? reg_mip_reserved_2 : _GEN_738;
  wire  _GEN_789 = io_req_bits_addr == 12'h103 ? reg_mip_SEIP : _GEN_739;
  wire  _GEN_790 = io_req_bits_addr == 12'h103 ? reg_mip_UEIP : _GEN_740;
  wire  _GEN_791 = io_req_bits_addr == 12'h103 ? reg_mip_MTIP : _GEN_741;
  wire  _GEN_792 = io_req_bits_addr == 12'h103 ? reg_mip_reserved_3 : _GEN_742;
  wire  _GEN_793 = io_req_bits_addr == 12'h103 ? reg_mip_STIP : _GEN_743;
  wire  _GEN_794 = io_req_bits_addr == 12'h103 ? reg_mip_UTIP : _GEN_744;
  wire  _GEN_795 = io_req_bits_addr == 12'h103 ? reg_mip_MSIP : _GEN_745;
  wire  _GEN_796 = io_req_bits_addr == 12'h103 ? reg_mip_reserved_4 : _GEN_746;
  wire  _GEN_797 = io_req_bits_addr == 12'h103 ? reg_mip_SSIP : _GEN_747;
  wire  _GEN_798 = io_req_bits_addr == 12'h103 ? reg_mip_USIP : _GEN_748;
  wire [63:0] _GEN_799 = io_req_bits_addr == 12'h103 ? reg_pmpcfg0 : _GEN_749;
  wire [63:0] _GEN_800 = io_req_bits_addr == 12'h103 ? reg_pmpcfg1 : _GEN_750;
  wire [63:0] _GEN_801 = io_req_bits_addr == 12'h103 ? reg_pmpcfg2 : _GEN_751;
  wire [63:0] _GEN_802 = io_req_bits_addr == 12'h103 ? reg_pmpcfg3 : _GEN_752;
  wire [63:0] _GEN_803 = io_req_bits_addr == 12'h103 ? reg_pmpaddr0 : _GEN_753;
  wire [63:0] _GEN_804 = io_req_bits_addr == 12'h102 ? write_data : reg_sedeleg;
  wire [63:0] _GEN_805 = io_req_bits_addr == 12'h102 ? reg_sideleg : _GEN_754;
  wire [63:0] _GEN_806 = io_req_bits_addr == 12'h102 ? reg_sie : _GEN_755;
  wire [63:0] _GEN_807 = io_req_bits_addr == 12'h102 ? reg_stvec : _GEN_756;
  wire [63:0] _GEN_808 = io_req_bits_addr == 12'h102 ? reg_scounteren : _GEN_757;
  wire [63:0] _GEN_809 = io_req_bits_addr == 12'h102 ? reg_sscratch : _GEN_758;
  wire [63:0] _GEN_810 = io_req_bits_addr == 12'h102 ? reg_scause : _GEN_759;
  wire [63:0] _GEN_811 = io_req_bits_addr == 12'h102 ? reg_stval : _GEN_760;
  wire [63:0] _GEN_812 = io_req_bits_addr == 12'h102 ? reg_sip : _GEN_761;
  wire [63:0] _GEN_813 = io_req_bits_addr == 12'h102 ? _GEN_6 : _GEN_762;
  wire [63:0] _GEN_814 = io_req_bits_addr == 12'h102 ? reg_misa : _GEN_763;
  wire [63:0] _GEN_815 = io_req_bits_addr == 12'h102 ? reg_medeleg : _GEN_764;
  wire [63:0] _GEN_816 = io_req_bits_addr == 12'h102 ? reg_mideleg : _GEN_765;
  wire [63:0] _GEN_817 = io_req_bits_addr == 12'h102 ? reg_mie : _GEN_766;
  wire [61:0] _GEN_818 = io_req_bits_addr == 12'h102 ? reg_mtvec_BASE : _GEN_767;
  wire [1:0] _GEN_819 = io_req_bits_addr == 12'h102 ? reg_mtvec_MODE : _GEN_768;
  wire [63:0] _GEN_820 = io_req_bits_addr == 12'h102 ? reg_mscratch : _GEN_769;
  wire [63:0] _GEN_821 = io_req_bits_addr == 12'h102 ? _GEN_2 : _GEN_770;
  wire  _GEN_822 = io_req_bits_addr == 12'h102 ? _GEN_0 : _GEN_771;
  wire [62:0] _GEN_823 = io_req_bits_addr == 12'h102 ? _GEN_1 : _GEN_772;
  wire [63:0] _GEN_824 = io_req_bits_addr == 12'h102 ? reg_mtval : _GEN_773;
  wire [51:0] _GEN_825 = io_req_bits_addr == 12'h102 ? reg_mip_reserved : _GEN_774;
  wire  _GEN_826 = io_req_bits_addr == 12'h102 ? reg_mip_intr_e_m : _GEN_775;
  wire  _GEN_827 = io_req_bits_addr == 12'h102 ? reg_mip_intr_e_h : _GEN_776;
  wire  _GEN_828 = io_req_bits_addr == 12'h102 ? reg_mip_intr_e_s : _GEN_777;
  wire  _GEN_829 = io_req_bits_addr == 12'h102 ? reg_mip_intr_e_u : _GEN_778;
  wire  _GEN_830 = io_req_bits_addr == 12'h102 ? reg_mip_intr_t_m : _GEN_779;
  wire  _GEN_831 = io_req_bits_addr == 12'h102 ? reg_mip_intr_t_h : _GEN_780;
  wire  _GEN_832 = io_req_bits_addr == 12'h102 ? reg_mip_intr_t_s : _GEN_781;
  wire  _GEN_833 = io_req_bits_addr == 12'h102 ? reg_mip_intr_t_u : _GEN_782;
  wire  _GEN_834 = io_req_bits_addr == 12'h102 ? reg_mip_intr_s_m : _GEN_783;
  wire  _GEN_835 = io_req_bits_addr == 12'h102 ? reg_mip_intr_s_h : _GEN_784;
  wire  _GEN_836 = io_req_bits_addr == 12'h102 ? reg_mip_intr_s_s : _GEN_785;
  wire  _GEN_837 = io_req_bits_addr == 12'h102 ? reg_mip_intr_s_u : _GEN_786;
  wire  _GEN_838 = io_req_bits_addr == 12'h102 ? reg_mip_MEIP : _GEN_787;
  wire  _GEN_839 = io_req_bits_addr == 12'h102 ? reg_mip_reserved_2 : _GEN_788;
  wire  _GEN_840 = io_req_bits_addr == 12'h102 ? reg_mip_SEIP : _GEN_789;
  wire  _GEN_841 = io_req_bits_addr == 12'h102 ? reg_mip_UEIP : _GEN_790;
  wire  _GEN_842 = io_req_bits_addr == 12'h102 ? reg_mip_MTIP : _GEN_791;
  wire  _GEN_843 = io_req_bits_addr == 12'h102 ? reg_mip_reserved_3 : _GEN_792;
  wire  _GEN_844 = io_req_bits_addr == 12'h102 ? reg_mip_STIP : _GEN_793;
  wire  _GEN_845 = io_req_bits_addr == 12'h102 ? reg_mip_UTIP : _GEN_794;
  wire  _GEN_846 = io_req_bits_addr == 12'h102 ? reg_mip_MSIP : _GEN_795;
  wire  _GEN_847 = io_req_bits_addr == 12'h102 ? reg_mip_reserved_4 : _GEN_796;
  wire  _GEN_848 = io_req_bits_addr == 12'h102 ? reg_mip_SSIP : _GEN_797;
  wire  _GEN_849 = io_req_bits_addr == 12'h102 ? reg_mip_USIP : _GEN_798;
  wire [63:0] _GEN_850 = io_req_bits_addr == 12'h102 ? reg_pmpcfg0 : _GEN_799;
  wire [63:0] _GEN_851 = io_req_bits_addr == 12'h102 ? reg_pmpcfg1 : _GEN_800;
  wire [63:0] _GEN_852 = io_req_bits_addr == 12'h102 ? reg_pmpcfg2 : _GEN_801;
  wire [63:0] _GEN_853 = io_req_bits_addr == 12'h102 ? reg_pmpcfg3 : _GEN_802;
  wire [63:0] _GEN_854 = io_req_bits_addr == 12'h102 ? reg_pmpaddr0 : _GEN_803;
  wire [63:0] _GEN_855 = io_req_bits_addr == 12'h100 ? write_data : reg_sstatus;
  wire [63:0] _GEN_856 = io_req_bits_addr == 12'h100 ? reg_sedeleg : _GEN_804;
  wire [63:0] _GEN_857 = io_req_bits_addr == 12'h100 ? reg_sideleg : _GEN_805;
  wire [63:0] _GEN_858 = io_req_bits_addr == 12'h100 ? reg_sie : _GEN_806;
  wire [63:0] _GEN_859 = io_req_bits_addr == 12'h100 ? reg_stvec : _GEN_807;
  wire [63:0] _GEN_860 = io_req_bits_addr == 12'h100 ? reg_scounteren : _GEN_808;
  wire [63:0] _GEN_861 = io_req_bits_addr == 12'h100 ? reg_sscratch : _GEN_809;
  wire [63:0] _GEN_862 = io_req_bits_addr == 12'h100 ? reg_scause : _GEN_810;
  wire [63:0] _GEN_863 = io_req_bits_addr == 12'h100 ? reg_stval : _GEN_811;
  wire [63:0] _GEN_864 = io_req_bits_addr == 12'h100 ? reg_sip : _GEN_812;
  wire [63:0] _GEN_865 = io_req_bits_addr == 12'h100 ? _GEN_6 : _GEN_813;
  wire [63:0] _GEN_866 = io_req_bits_addr == 12'h100 ? reg_misa : _GEN_814;
  wire [63:0] _GEN_867 = io_req_bits_addr == 12'h100 ? reg_medeleg : _GEN_815;
  wire [63:0] _GEN_868 = io_req_bits_addr == 12'h100 ? reg_mideleg : _GEN_816;
  wire [63:0] _GEN_869 = io_req_bits_addr == 12'h100 ? reg_mie : _GEN_817;
  wire [61:0] _GEN_870 = io_req_bits_addr == 12'h100 ? reg_mtvec_BASE : _GEN_818;
  wire [1:0] _GEN_871 = io_req_bits_addr == 12'h100 ? reg_mtvec_MODE : _GEN_819;
  wire [63:0] _GEN_872 = io_req_bits_addr == 12'h100 ? reg_mscratch : _GEN_820;
  wire [63:0] _GEN_873 = io_req_bits_addr == 12'h100 ? _GEN_2 : _GEN_821;
  wire  _GEN_874 = io_req_bits_addr == 12'h100 ? _GEN_0 : _GEN_822;
  wire [62:0] _GEN_875 = io_req_bits_addr == 12'h100 ? _GEN_1 : _GEN_823;
  wire [63:0] _GEN_876 = io_req_bits_addr == 12'h100 ? reg_mtval : _GEN_824;
  wire [51:0] _GEN_877 = io_req_bits_addr == 12'h100 ? reg_mip_reserved : _GEN_825;
  wire  _GEN_878 = io_req_bits_addr == 12'h100 ? reg_mip_intr_e_m : _GEN_826;
  wire  _GEN_879 = io_req_bits_addr == 12'h100 ? reg_mip_intr_e_h : _GEN_827;
  wire  _GEN_880 = io_req_bits_addr == 12'h100 ? reg_mip_intr_e_s : _GEN_828;
  wire  _GEN_881 = io_req_bits_addr == 12'h100 ? reg_mip_intr_e_u : _GEN_829;
  wire  _GEN_882 = io_req_bits_addr == 12'h100 ? reg_mip_intr_t_m : _GEN_830;
  wire  _GEN_883 = io_req_bits_addr == 12'h100 ? reg_mip_intr_t_h : _GEN_831;
  wire  _GEN_884 = io_req_bits_addr == 12'h100 ? reg_mip_intr_t_s : _GEN_832;
  wire  _GEN_885 = io_req_bits_addr == 12'h100 ? reg_mip_intr_t_u : _GEN_833;
  wire  _GEN_886 = io_req_bits_addr == 12'h100 ? reg_mip_intr_s_m : _GEN_834;
  wire  _GEN_887 = io_req_bits_addr == 12'h100 ? reg_mip_intr_s_h : _GEN_835;
  wire  _GEN_888 = io_req_bits_addr == 12'h100 ? reg_mip_intr_s_s : _GEN_836;
  wire  _GEN_889 = io_req_bits_addr == 12'h100 ? reg_mip_intr_s_u : _GEN_837;
  wire  _GEN_890 = io_req_bits_addr == 12'h100 ? reg_mip_MEIP : _GEN_838;
  wire  _GEN_891 = io_req_bits_addr == 12'h100 ? reg_mip_reserved_2 : _GEN_839;
  wire  _GEN_892 = io_req_bits_addr == 12'h100 ? reg_mip_SEIP : _GEN_840;
  wire  _GEN_893 = io_req_bits_addr == 12'h100 ? reg_mip_UEIP : _GEN_841;
  wire  _GEN_894 = io_req_bits_addr == 12'h100 ? reg_mip_MTIP : _GEN_842;
  wire  _GEN_895 = io_req_bits_addr == 12'h100 ? reg_mip_reserved_3 : _GEN_843;
  wire  _GEN_896 = io_req_bits_addr == 12'h100 ? reg_mip_STIP : _GEN_844;
  wire  _GEN_897 = io_req_bits_addr == 12'h100 ? reg_mip_UTIP : _GEN_845;
  wire  _GEN_898 = io_req_bits_addr == 12'h100 ? reg_mip_MSIP : _GEN_846;
  wire  _GEN_899 = io_req_bits_addr == 12'h100 ? reg_mip_reserved_4 : _GEN_847;
  wire  _GEN_900 = io_req_bits_addr == 12'h100 ? reg_mip_SSIP : _GEN_848;
  wire  _GEN_901 = io_req_bits_addr == 12'h100 ? reg_mip_USIP : _GEN_849;
  wire [63:0] _GEN_902 = io_req_bits_addr == 12'h100 ? reg_pmpcfg0 : _GEN_850;
  wire [63:0] _GEN_903 = io_req_bits_addr == 12'h100 ? reg_pmpcfg1 : _GEN_851;
  wire [63:0] _GEN_904 = io_req_bits_addr == 12'h100 ? reg_pmpcfg2 : _GEN_852;
  wire [63:0] _GEN_905 = io_req_bits_addr == 12'h100 ? reg_pmpcfg3 : _GEN_853;
  wire [63:0] _GEN_906 = io_req_bits_addr == 12'h100 ? reg_pmpaddr0 : _GEN_854;
  wire [63:0] _GEN_907 = io_req_bits_addr == 12'hf14 ? write_data : reg_mhartid;
  wire [63:0] _GEN_908 = io_req_bits_addr == 12'hf14 ? reg_sstatus : _GEN_855;
  wire [63:0] _GEN_909 = io_req_bits_addr == 12'hf14 ? reg_sedeleg : _GEN_856;
  wire [63:0] _GEN_910 = io_req_bits_addr == 12'hf14 ? reg_sideleg : _GEN_857;
  wire [63:0] _GEN_911 = io_req_bits_addr == 12'hf14 ? reg_sie : _GEN_858;
  wire [63:0] _GEN_912 = io_req_bits_addr == 12'hf14 ? reg_stvec : _GEN_859;
  wire [63:0] _GEN_913 = io_req_bits_addr == 12'hf14 ? reg_scounteren : _GEN_860;
  wire [63:0] _GEN_914 = io_req_bits_addr == 12'hf14 ? reg_sscratch : _GEN_861;
  wire [63:0] _GEN_915 = io_req_bits_addr == 12'hf14 ? reg_scause : _GEN_862;
  wire [63:0] _GEN_916 = io_req_bits_addr == 12'hf14 ? reg_stval : _GEN_863;
  wire [63:0] _GEN_917 = io_req_bits_addr == 12'hf14 ? reg_sip : _GEN_864;
  wire [63:0] _GEN_918 = io_req_bits_addr == 12'hf14 ? _GEN_6 : _GEN_865;
  wire [63:0] _GEN_919 = io_req_bits_addr == 12'hf14 ? reg_misa : _GEN_866;
  wire [63:0] _GEN_920 = io_req_bits_addr == 12'hf14 ? reg_medeleg : _GEN_867;
  wire [63:0] _GEN_921 = io_req_bits_addr == 12'hf14 ? reg_mideleg : _GEN_868;
  wire [63:0] _GEN_922 = io_req_bits_addr == 12'hf14 ? reg_mie : _GEN_869;
  wire [61:0] _GEN_923 = io_req_bits_addr == 12'hf14 ? reg_mtvec_BASE : _GEN_870;
  wire [1:0] _GEN_924 = io_req_bits_addr == 12'hf14 ? reg_mtvec_MODE : _GEN_871;
  wire [63:0] _GEN_925 = io_req_bits_addr == 12'hf14 ? reg_mscratch : _GEN_872;
  wire [63:0] _GEN_926 = io_req_bits_addr == 12'hf14 ? _GEN_2 : _GEN_873;
  wire  _GEN_927 = io_req_bits_addr == 12'hf14 ? _GEN_0 : _GEN_874;
  wire [62:0] _GEN_928 = io_req_bits_addr == 12'hf14 ? _GEN_1 : _GEN_875;
  wire [63:0] _GEN_929 = io_req_bits_addr == 12'hf14 ? reg_mtval : _GEN_876;
  wire [51:0] _GEN_930 = io_req_bits_addr == 12'hf14 ? reg_mip_reserved : _GEN_877;
  wire  _GEN_931 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_e_m : _GEN_878;
  wire  _GEN_932 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_e_h : _GEN_879;
  wire  _GEN_933 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_e_s : _GEN_880;
  wire  _GEN_934 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_e_u : _GEN_881;
  wire  _GEN_935 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_t_m : _GEN_882;
  wire  _GEN_936 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_t_h : _GEN_883;
  wire  _GEN_937 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_t_s : _GEN_884;
  wire  _GEN_938 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_t_u : _GEN_885;
  wire  _GEN_939 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_s_m : _GEN_886;
  wire  _GEN_940 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_s_h : _GEN_887;
  wire  _GEN_941 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_s_s : _GEN_888;
  wire  _GEN_942 = io_req_bits_addr == 12'hf14 ? reg_mip_intr_s_u : _GEN_889;
  wire  _GEN_943 = io_req_bits_addr == 12'hf14 ? reg_mip_MEIP : _GEN_890;
  wire  _GEN_944 = io_req_bits_addr == 12'hf14 ? reg_mip_reserved_2 : _GEN_891;
  wire  _GEN_945 = io_req_bits_addr == 12'hf14 ? reg_mip_SEIP : _GEN_892;
  wire  _GEN_946 = io_req_bits_addr == 12'hf14 ? reg_mip_UEIP : _GEN_893;
  wire  _GEN_947 = io_req_bits_addr == 12'hf14 ? reg_mip_MTIP : _GEN_894;
  wire  _GEN_948 = io_req_bits_addr == 12'hf14 ? reg_mip_reserved_3 : _GEN_895;
  wire  _GEN_949 = io_req_bits_addr == 12'hf14 ? reg_mip_STIP : _GEN_896;
  wire  _GEN_950 = io_req_bits_addr == 12'hf14 ? reg_mip_UTIP : _GEN_897;
  wire  _GEN_951 = io_req_bits_addr == 12'hf14 ? reg_mip_MSIP : _GEN_898;
  wire  _GEN_952 = io_req_bits_addr == 12'hf14 ? reg_mip_reserved_4 : _GEN_899;
  wire  _GEN_953 = io_req_bits_addr == 12'hf14 ? reg_mip_SSIP : _GEN_900;
  wire  _GEN_954 = io_req_bits_addr == 12'hf14 ? reg_mip_USIP : _GEN_901;
  wire [63:0] _GEN_955 = io_req_bits_addr == 12'hf14 ? reg_pmpcfg0 : _GEN_902;
  wire [63:0] _GEN_956 = io_req_bits_addr == 12'hf14 ? reg_pmpcfg1 : _GEN_903;
  wire [63:0] _GEN_957 = io_req_bits_addr == 12'hf14 ? reg_pmpcfg2 : _GEN_904;
  wire [63:0] _GEN_958 = io_req_bits_addr == 12'hf14 ? reg_pmpcfg3 : _GEN_905;
  wire [63:0] _GEN_959 = io_req_bits_addr == 12'hf14 ? reg_pmpaddr0 : _GEN_906;
  assign io_resp_bits_rdata = io_req_bits_rd == 5'h0 ? 64'h0 : read_csr_data;
  assign io_redirect_valid = raiseExceptionIntr | isMret;
  assign io_redirect_target = _io_redirect_target_T[31:0];
  assign io_en = |_raiseException_T;
  assign io_raiseIntr = |intrVec;
  always @(posedge clock) begin
    if (reset) begin
      mode <= 2'h3;
    end else if (isMret) begin
      mode <= mstatusStruct_MPP;
    end else if (raiseExceptionIntr) begin
      mode <= 2'h3;
    end
    if (reset) begin
      reg_satp <= 64'h0;
    end else if (wen) begin
      if (io_req_bits_addr == 12'h180) begin
        if (6'h30 == io_req_bits_cmd) begin
          reg_satp <= _write_data_T_6;
        end else begin
          reg_satp <= _write_data_T_10;
        end
      end
    end
    if (reset) begin
      reg_sepc <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (io_req_bits_addr == 12'h141) begin
          reg_sepc <= write_data;
        end
      end
    end
    if (reset) begin
      reg_sstatus <= 64'h200000000;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sstatus <= _GEN_908;
        end
      end
    end
    if (reset) begin
      reg_sedeleg <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sedeleg <= _GEN_909;
        end
      end
    end
    if (reset) begin
      reg_sideleg <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sideleg <= _GEN_910;
        end
      end
    end
    if (reset) begin
      reg_sie <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sie <= _GEN_911;
        end
      end
    end
    if (reset) begin
      reg_stvec <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_stvec <= _GEN_912;
        end
      end
    end
    if (reset) begin
      reg_scounteren <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_scounteren <= _GEN_913;
        end
      end
    end
    if (reset) begin
      reg_sscratch <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sscratch <= _GEN_914;
        end
      end
    end
    if (reset) begin
      reg_scause <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_scause <= _GEN_915;
        end
      end
    end
    if (reset) begin
      reg_stval <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_stval <= _GEN_916;
        end
      end
    end
    if (reset) begin
      reg_sip <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_sip <= _GEN_917;
        end
      end
    end
    if (reset) begin
      reg_mhartid <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mhartid <= _GEN_907;
        end
      end
    end
    if (reset) begin
      reg_mstatus <= 64'ha00001800;
    end else if (wen) begin
      if (io_req_bits_addr == 12'h180) begin
        reg_mstatus <= _GEN_6;
      end else if (io_req_bits_addr == 12'h141) begin
        reg_mstatus <= _GEN_6;
      end else begin
        reg_mstatus <= _GEN_918;
      end
    end else begin
      reg_mstatus <= _GEN_6;
    end
    if (reset) begin
      reg_misa <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_misa <= _GEN_919;
        end
      end
    end
    if (reset) begin
      reg_medeleg <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_medeleg <= _GEN_920;
        end
      end
    end
    if (reset) begin
      reg_mideleg <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mideleg <= _GEN_921;
        end
      end
    end
    if (reset) begin
      reg_mie <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mie <= _GEN_922;
        end
      end
    end
    if (reset) begin
      reg_mtvec_BASE <= 62'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mtvec_BASE <= _GEN_923;
        end
      end
    end
    if (reset) begin
      reg_mtvec_MODE <= 2'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mtvec_MODE <= _GEN_924;
        end
      end
    end
    if (reset) begin
      reg_mscratch <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mscratch <= _GEN_925;
        end
      end
    end
    if (reset) begin
      reg_mepc <= 64'h0;
    end else if (wen) begin
      if (io_req_bits_addr == 12'h180) begin
        reg_mepc <= _GEN_2;
      end else if (io_req_bits_addr == 12'h141) begin
        reg_mepc <= _GEN_2;
      end else begin
        reg_mepc <= _GEN_926;
      end
    end else begin
      reg_mepc <= _GEN_2;
    end
    if (reset) begin
      reg_mcause_interrupt <= 1'h0;
    end else if (wen) begin
      if (io_req_bits_addr == 12'h180) begin
        reg_mcause_interrupt <= _GEN_0;
      end else if (io_req_bits_addr == 12'h141) begin
        reg_mcause_interrupt <= _GEN_0;
      end else begin
        reg_mcause_interrupt <= _GEN_927;
      end
    end else begin
      reg_mcause_interrupt <= _GEN_0;
    end
    if (reset) begin
      reg_mcause_exc_code <= 63'h0;
    end else if (wen) begin
      if (io_req_bits_addr == 12'h180) begin
        reg_mcause_exc_code <= _GEN_1;
      end else if (io_req_bits_addr == 12'h141) begin
        reg_mcause_exc_code <= _GEN_1;
      end else begin
        reg_mcause_exc_code <= _GEN_928;
      end
    end else begin
      reg_mcause_exc_code <= _GEN_1;
    end
    if (reset) begin
      reg_mtval <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mtval <= _GEN_929;
        end
      end
    end
    if (reset) begin
      reg_mip_reserved <= 52'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_reserved <= _GEN_930;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_e_m <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_e_m <= _GEN_931;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_e_h <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_e_h <= _GEN_932;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_e_s <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_e_s <= _GEN_933;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_e_u <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_e_u <= _GEN_934;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_t_m <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_t_m <= _GEN_935;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_t_h <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_t_h <= _GEN_936;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_t_s <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_t_s <= _GEN_937;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_t_u <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_t_u <= _GEN_938;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_s_m <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_s_m <= _GEN_939;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_s_h <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_s_h <= _GEN_940;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_s_s <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_s_s <= _GEN_941;
        end
      end
    end
    if (reset) begin
      reg_mip_intr_s_u <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_intr_s_u <= _GEN_942;
        end
      end
    end
    if (reset) begin
      reg_mip_MEIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_MEIP <= _GEN_943;
        end
      end
    end
    if (reset) begin
      reg_mip_reserved_2 <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_reserved_2 <= _GEN_944;
        end
      end
    end
    if (reset) begin
      reg_mip_SEIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_SEIP <= _GEN_945;
        end
      end
    end
    if (reset) begin
      reg_mip_UEIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_UEIP <= _GEN_946;
        end
      end
    end
    if (reset) begin
      reg_mip_MTIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_MTIP <= _GEN_947;
        end
      end
    end
    if (reset) begin
      reg_mip_reserved_3 <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_reserved_3 <= _GEN_948;
        end
      end
    end
    if (reset) begin
      reg_mip_STIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_STIP <= _GEN_949;
        end
      end
    end
    if (reset) begin
      reg_mip_UTIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_UTIP <= _GEN_950;
        end
      end
    end
    if (reset) begin
      reg_mip_MSIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_MSIP <= _GEN_951;
        end
      end
    end
    if (reset) begin
      reg_mip_reserved_4 <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_reserved_4 <= _GEN_952;
        end
      end
    end
    if (reset) begin
      reg_mip_SSIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_SSIP <= _GEN_953;
        end
      end
    end
    if (reset) begin
      reg_mip_USIP <= 1'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_mip_USIP <= _GEN_954;
        end
      end
    end
    if (reset) begin
      reg_pmpcfg0 <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_pmpcfg0 <= _GEN_955;
        end
      end
    end
    if (reset) begin
      reg_pmpcfg1 <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_pmpcfg1 <= _GEN_956;
        end
      end
    end
    if (reset) begin
      reg_pmpcfg2 <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_pmpcfg2 <= _GEN_957;
        end
      end
    end
    if (reset) begin
      reg_pmpcfg3 <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_pmpcfg3 <= _GEN_958;
        end
      end
    end
    if (reset) begin
      reg_pmpaddr0 <= 64'h0;
    end else if (wen) begin
      if (!(io_req_bits_addr == 12'h180)) begin
        if (!(io_req_bits_addr == 12'h141)) begin
          reg_pmpaddr0 <= _GEN_959;
        end
      end
    end
    if (reset) begin
      mcycle <= 64'h0;
    end else begin
      mcycle <= _mcycle_T_1;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mode = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  reg_satp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  reg_sepc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_sstatus = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  reg_sedeleg = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_sideleg = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  reg_sie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_stvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  reg_scounteren = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  reg_sscratch = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  reg_scause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  reg_stval = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  reg_sip = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  reg_mhartid = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  reg_mstatus = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  reg_misa = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  reg_medeleg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  reg_mideleg = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_mie = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_mtvec_BASE = _RAND_19[61:0];
  _RAND_20 = {1{`RANDOM}};
  reg_mtvec_MODE = _RAND_20[1:0];
  _RAND_21 = {2{`RANDOM}};
  reg_mscratch = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  reg_mepc = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  reg_mcause_interrupt = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  reg_mcause_exc_code = _RAND_24[62:0];
  _RAND_25 = {2{`RANDOM}};
  reg_mtval = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  reg_mip_reserved = _RAND_26[51:0];
  _RAND_27 = {1{`RANDOM}};
  reg_mip_intr_e_m = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  reg_mip_intr_e_h = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  reg_mip_intr_e_s = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  reg_mip_intr_e_u = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  reg_mip_intr_t_m = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  reg_mip_intr_t_h = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  reg_mip_intr_t_s = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  reg_mip_intr_t_u = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  reg_mip_intr_s_m = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  reg_mip_intr_s_h = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  reg_mip_intr_s_s = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  reg_mip_intr_s_u = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  reg_mip_MEIP = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  reg_mip_reserved_2 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  reg_mip_SEIP = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  reg_mip_UEIP = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  reg_mip_MTIP = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  reg_mip_reserved_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  reg_mip_STIP = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  reg_mip_UTIP = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  reg_mip_MSIP = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  reg_mip_reserved_4 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  reg_mip_SSIP = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  reg_mip_USIP = _RAND_50[0:0];
  _RAND_51 = {2{`RANDOM}};
  reg_pmpcfg0 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  reg_pmpcfg1 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  reg_pmpcfg2 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  reg_pmpcfg3 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  reg_pmpaddr0 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  mcycle = _RAND_56[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Mou(
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [5:0]  io_in_bits_func,
  output        io_out_bits_redirect_valid,
  output [31:0] io_out_bits_redirect_target,
  output        flushICache_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 6'h2b;
  assign io_out_bits_redirect_valid = io_in_valid;
  assign io_out_bits_redirect_target = io_in_bits_pc + 32'h4;
  assign flushICache_0 = flushICache;
endmodule
module ysyx_040656_ExecuteStage(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [31:0] io_in_bits_inst,
  input         io_in_bits_valid,
  input         io_in_bits_bubble,
  input  [2:0]  io_in_bits_opcode_type,
  input  [5:0]  io_in_bits_opcode_func,
  input  [3:0]  io_in_bits_br_type,
  input         io_in_bits_rf_en,
  input  [4:0]  io_in_bits_wb_addr,
  input  [1:0]  io_in_bits_wb_stage,
  input  [63:0] io_in_bits_op1_data,
  input  [63:0] io_in_bits_op2_data,
  input  [63:0] io_in_bits_rs1_data,
  input  [63:0] io_in_bits_rs2_data,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [1:0]  io_dmem_req_bits_size,
  output [2:0]  io_dmem_req_bits_cmd,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [63:0] io_mmio_req_bits_wdata,
  output [1:0]  io_mmio_req_bits_size,
  output [2:0]  io_mmio_req_bits_cmd,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_valid,
  output        io_out_bits_wen,
  output [4:0]  io_out_bits_wb_addr,
  output [63:0] io_out_bits_wb_data,
  output        io_out_bits_redirect_valid,
  output [31:0] io_out_bits_redirect_target,
  output        io_bypass_rf_wen,
  output [4:0]  io_bypass_addr,
  output [63:0] io_bypass_data,
  output        flushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif
  wire [63:0] alu_io_in_bits_op1_data;
  wire [63:0] alu_io_in_bits_op2_data;
  wire [5:0] alu_io_in_bits_func;
  wire [63:0] alu_io_out_bits;
  wire  jmp_io_in_valid;
  wire [63:0] jmp_io_in_bits_op1_data;
  wire [63:0] jmp_io_in_bits_op2_data;
  wire [63:0] jmp_io_in_bits_rs1_data;
  wire [63:0] jmp_io_in_bits_rs2_data;
  wire [3:0] jmp_io_in_bits_br_type;
  wire [31:0] jmp_io_in_bits_pc;
  wire  jmp_io_out_bits_redirect_valid;
  wire [31:0] jmp_io_out_bits_redirect_target;
  wire  mdu_clock;
  wire  mdu_reset;
  wire  mdu_io_in_valid;
  wire [63:0] mdu_io_in_bits_op1_data;
  wire [63:0] mdu_io_in_bits_op2_data;
  wire [5:0] mdu_io_in_bits_func;
  wire  mdu_io_out_valid;
  wire [63:0] mdu_io_out_bits;
  wire  lsu_clock;
  wire  lsu_reset;
  wire  lsu_io_in_valid;
  wire [31:0] lsu_io_in_bits_addr;
  wire [5:0] lsu_io_in_bits_func;
  wire [63:0] lsu_io_in_bits_rs2_data;
  wire  lsu_io_out_valid;
  wire [63:0] lsu_io_out_bits_data;
  wire  lsu_io_dmem_req_ready;
  wire  lsu_io_dmem_req_valid;
  wire [31:0] lsu_io_dmem_req_bits_addr;
  wire [63:0] lsu_io_dmem_req_bits_wdata;
  wire [1:0] lsu_io_dmem_req_bits_size;
  wire [2:0] lsu_io_dmem_req_bits_cmd;
  wire  lsu_io_dmem_resp_ready;
  wire  lsu_io_dmem_resp_valid;
  wire [63:0] lsu_io_dmem_resp_bits_rdata;
  wire  lsu_io_mmio_req_ready;
  wire  lsu_io_mmio_req_valid;
  wire [31:0] lsu_io_mmio_req_bits_addr;
  wire [63:0] lsu_io_mmio_req_bits_wdata;
  wire [1:0] lsu_io_mmio_req_bits_size;
  wire [2:0] lsu_io_mmio_req_bits_cmd;
  wire  lsu_io_mmio_resp_ready;
  wire  lsu_io_mmio_resp_valid;
  wire [63:0] lsu_io_mmio_resp_bits_rdata;
  wire  csr_clock;
  wire  csr_reset;
  wire  csr_io_req_valid;
  wire [31:0] csr_io_req_bits_pc;
  wire [5:0] csr_io_req_bits_cmd;
  wire [11:0] csr_io_req_bits_addr;
  wire [63:0] csr_io_req_bits_wdata;
  wire [4:0] csr_io_req_bits_rd;
  wire  csr_io_req_bits_valid;
  wire [63:0] csr_io_resp_bits_rdata;
  wire  csr_io_redirect_valid;
  wire [31:0] csr_io_redirect_target;
  wire  csr_io_en;
  wire  csr_io_raiseIntr;
  wire  mou_io_in_valid;
  wire [31:0] mou_io_in_bits_pc;
  wire [5:0] mou_io_in_bits_func;
  wire  mou_io_out_bits_redirect_valid;
  wire [31:0] mou_io_out_bits_redirect_target;
  wire  mou_flushICache_0;
  reg  executeNop_valid;
  reg  executeNop_bubble;
  reg [2:0] executeNop_opcode_type;
  reg [5:0] executeNop_opcode_func;
  reg [31:0] executeBuffer_pc;
  reg [31:0] executeBuffer_inst;
  reg  executeBuffer_valid;
  reg  executeBuffer_bubble;
  reg [2:0] executeBuffer_opcode_type;
  reg [5:0] executeBuffer_opcode_func;
  reg [3:0] executeBuffer_br_type;
  reg  executeBuffer_rf_en;
  reg [4:0] executeBuffer_wb_addr;
  reg [1:0] executeBuffer_wb_stage;
  reg [63:0] executeBuffer_op1_data;
  reg [63:0] executeBuffer_op2_data;
  reg [63:0] executeBuffer_rs1_data;
  reg [63:0] executeBuffer_rs2_data;
  wire  _T_1 = ~io_flush;
  wire  isLSU = executeBuffer_opcode_type == 3'h2 & _T_1;
  wire  isCSR = executeBuffer_opcode_type == 3'h3 & _T_1;
  wire  isMDU = executeBuffer_opcode_type == 3'h5 & _T_1;
  wire  _lsuOut_T_1 = isLSU & ~csr_io_raiseIntr;
  wire [63:0] _lsuOut_T_3 = executeBuffer_op1_data + executeBuffer_op2_data;
  wire [63:0] _executeOutput_T_7 = 3'h1 == executeBuffer_opcode_type ? alu_io_out_bits : 64'h0;
  wire [63:0] _executeOutput_T_9 = 3'h2 == executeBuffer_opcode_type ? lsu_io_out_bits_data : _executeOutput_T_7;
  wire [63:0] _executeOutput_T_11 = 3'h5 == executeBuffer_opcode_type ? mdu_io_out_bits : _executeOutput_T_9;
  wire [63:0] _executeOutput_T_13 = 3'h6 == executeBuffer_opcode_type ? {{32'd0}, jmp_io_out_bits_redirect_target} :
    _executeOutput_T_11;
  wire [63:0] executeOutput = 3'h3 == executeBuffer_opcode_type ? csr_io_resp_bits_rdata : _executeOutput_T_13;
  wire  _outValid_T_2 = isMDU ? mdu_io_out_valid : 1'h1;
  wire [31:0] _wb_data_T_4 = executeBuffer_pc + 32'h4;
  wire [63:0] _wb_data_T_7 = 2'h1 == executeBuffer_wb_stage ? executeOutput : 64'h0;
  wire [63:0] _wb_data_T_9 = 2'h2 == executeBuffer_wb_stage ? {{32'd0}, _wb_data_T_4} : _wb_data_T_7;
  wire [31:0] _io_out_bits_redirect_target_T = csr_io_redirect_valid ? csr_io_redirect_target :
    jmp_io_out_bits_redirect_target;
  ysyx_040656_Alu alu (
    .io_in_bits_op1_data(alu_io_in_bits_op1_data),
    .io_in_bits_op2_data(alu_io_in_bits_op2_data),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_bits(alu_io_out_bits)
  );
  ysyx_040656_Jmp jmp (
    .io_in_valid(jmp_io_in_valid),
    .io_in_bits_op1_data(jmp_io_in_bits_op1_data),
    .io_in_bits_op2_data(jmp_io_in_bits_op2_data),
    .io_in_bits_rs1_data(jmp_io_in_bits_rs1_data),
    .io_in_bits_rs2_data(jmp_io_in_bits_rs2_data),
    .io_in_bits_br_type(jmp_io_in_bits_br_type),
    .io_in_bits_pc(jmp_io_in_bits_pc),
    .io_out_bits_redirect_valid(jmp_io_out_bits_redirect_valid),
    .io_out_bits_redirect_target(jmp_io_out_bits_redirect_target)
  );
  ysyx_040656_Mdu mdu (
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_op1_data(mdu_io_in_bits_op1_data),
    .io_in_bits_op2_data(mdu_io_in_bits_op2_data),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  ysyx_040656_Lsu lsu (
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_in_valid(lsu_io_in_valid),
    .io_in_bits_addr(lsu_io_in_bits_addr),
    .io_in_bits_func(lsu_io_in_bits_func),
    .io_in_bits_rs2_data(lsu_io_in_bits_rs2_data),
    .io_out_valid(lsu_io_out_valid),
    .io_out_bits_data(lsu_io_out_bits_data),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_addr(lsu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(lsu_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_size(lsu_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(lsu_io_dmem_req_bits_cmd),
    .io_dmem_resp_ready(lsu_io_dmem_resp_ready),
    .io_dmem_resp_valid(lsu_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(lsu_io_dmem_resp_bits_rdata),
    .io_mmio_req_ready(lsu_io_mmio_req_ready),
    .io_mmio_req_valid(lsu_io_mmio_req_valid),
    .io_mmio_req_bits_addr(lsu_io_mmio_req_bits_addr),
    .io_mmio_req_bits_wdata(lsu_io_mmio_req_bits_wdata),
    .io_mmio_req_bits_size(lsu_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(lsu_io_mmio_req_bits_cmd),
    .io_mmio_resp_ready(lsu_io_mmio_resp_ready),
    .io_mmio_resp_valid(lsu_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(lsu_io_mmio_resp_bits_rdata)
  );
  ysyx_040656_Csr csr (
    .clock(csr_clock),
    .reset(csr_reset),
    .io_req_valid(csr_io_req_valid),
    .io_req_bits_pc(csr_io_req_bits_pc),
    .io_req_bits_cmd(csr_io_req_bits_cmd),
    .io_req_bits_addr(csr_io_req_bits_addr),
    .io_req_bits_wdata(csr_io_req_bits_wdata),
    .io_req_bits_rd(csr_io_req_bits_rd),
    .io_req_bits_valid(csr_io_req_bits_valid),
    .io_resp_bits_rdata(csr_io_resp_bits_rdata),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_redirect_target(csr_io_redirect_target),
    .io_en(csr_io_en),
    .io_raiseIntr(csr_io_raiseIntr)
  );
  ysyx_040656_Mou mou (
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_pc(mou_io_in_bits_pc),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_out_bits_redirect_valid(mou_io_out_bits_redirect_valid),
    .io_out_bits_redirect_target(mou_io_out_bits_redirect_target),
    .flushICache_0(mou_flushICache_0)
  );
  assign io_in_ready = io_out_valid | executeBuffer_bubble;
  assign io_dmem_req_valid = lsu_io_dmem_req_valid;
  assign io_dmem_req_bits_addr = lsu_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_wdata = lsu_io_dmem_req_bits_wdata;
  assign io_dmem_req_bits_size = lsu_io_dmem_req_bits_size;
  assign io_dmem_req_bits_cmd = lsu_io_dmem_req_bits_cmd;
  assign io_mmio_req_valid = lsu_io_mmio_req_valid;
  assign io_mmio_req_bits_addr = lsu_io_mmio_req_bits_addr;
  assign io_mmio_req_bits_wdata = lsu_io_mmio_req_bits_wdata;
  assign io_mmio_req_bits_size = lsu_io_mmio_req_bits_size;
  assign io_mmio_req_bits_cmd = lsu_io_mmio_req_bits_cmd;
  assign io_out_valid = _lsuOut_T_1 ? lsu_io_out_valid : _outValid_T_2;
  assign io_out_bits_valid = executeBuffer_valid & ~executeBuffer_bubble;
  assign io_out_bits_wen = executeBuffer_rf_en & ~csr_io_en & executeBuffer_wb_addr >= 5'h1;
  assign io_out_bits_wb_addr = executeBuffer_wb_addr;
  assign io_out_bits_wb_data = 2'h0 == executeBuffer_wb_stage ? 64'h0 : _wb_data_T_9;
  assign io_out_bits_redirect_valid = jmp_io_out_bits_redirect_valid | csr_io_redirect_valid |
    mou_io_out_bits_redirect_valid;
  assign io_out_bits_redirect_target = mou_io_out_bits_redirect_valid ? mou_io_out_bits_redirect_target :
    _io_out_bits_redirect_target_T;
  assign io_bypass_rf_wen = executeBuffer_rf_en & ~csr_io_en & executeBuffer_wb_addr >= 5'h1;
  assign io_bypass_addr = executeBuffer_wb_addr;
  assign io_bypass_data = 2'h0 == executeBuffer_wb_stage ? 64'h0 : _wb_data_T_9;
  assign flushICache = mou_flushICache_0;
  assign alu_io_in_bits_op1_data = executeBuffer_op1_data;
  assign alu_io_in_bits_op2_data = executeBuffer_op2_data;
  assign alu_io_in_bits_func = executeBuffer_opcode_func;
  assign jmp_io_in_valid = executeBuffer_opcode_type == 3'h6 & _T_1;
  assign jmp_io_in_bits_op1_data = executeBuffer_op1_data;
  assign jmp_io_in_bits_op2_data = executeBuffer_op2_data;
  assign jmp_io_in_bits_rs1_data = executeBuffer_rs2_data;
  assign jmp_io_in_bits_rs2_data = executeBuffer_rs1_data;
  assign jmp_io_in_bits_br_type = executeBuffer_br_type;
  assign jmp_io_in_bits_pc = executeBuffer_pc;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = executeBuffer_opcode_type == 3'h5 & _T_1;
  assign mdu_io_in_bits_op1_data = executeBuffer_op1_data;
  assign mdu_io_in_bits_op2_data = executeBuffer_op2_data;
  assign mdu_io_in_bits_func = executeBuffer_opcode_func;
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_in_valid = isLSU & ~csr_io_raiseIntr;
  assign lsu_io_in_bits_addr = _lsuOut_T_3[31:0];
  assign lsu_io_in_bits_func = executeBuffer_opcode_func;
  assign lsu_io_in_bits_rs2_data = executeBuffer_rs2_data;
  assign lsu_io_dmem_req_ready = io_dmem_req_ready;
  assign lsu_io_dmem_resp_valid = io_dmem_resp_valid;
  assign lsu_io_dmem_resp_bits_rdata = io_dmem_resp_bits_rdata;
  assign lsu_io_mmio_req_ready = io_mmio_req_ready;
  assign lsu_io_mmio_resp_valid = io_mmio_resp_valid;
  assign lsu_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_req_valid = executeBuffer_opcode_type == 3'h3 & _T_1;
  assign csr_io_req_bits_pc = executeBuffer_pc;
  assign csr_io_req_bits_cmd = isCSR ? executeBuffer_opcode_func : 6'h2d;
  assign csr_io_req_bits_addr = executeBuffer_opcode_func == 6'h2d & isCSR ? 12'h0 : executeBuffer_inst[31:20];
  assign csr_io_req_bits_wdata = executeBuffer_op1_data;
  assign csr_io_req_bits_rd = executeBuffer_wb_addr;
  assign csr_io_req_bits_valid = executeBuffer_opcode_type == 3'h3 & _T_1;
  assign mou_io_in_valid = executeBuffer_opcode_type == 3'h4 & _T_1;
  assign mou_io_in_bits_pc = executeBuffer_pc;
  assign mou_io_in_bits_func = executeBuffer_opcode_func;
  always @(posedge clock) begin
    if (reset) begin
      executeNop_valid <= 1'h0;
    end else begin
      executeNop_valid <= 1'h1;
    end
    if (reset) begin
      executeNop_bubble <= 1'h0;
    end else begin
      executeNop_bubble <= 1'h1;
    end
    if (reset) begin
      executeNop_opcode_type <= 3'h0;
    end else begin
      executeNop_opcode_type <= 3'h1;
    end
    if (reset) begin
      executeNop_opcode_func <= 6'h0;
    end else begin
      executeNop_opcode_func <= 6'h2;
    end
    if (reset) begin
      executeBuffer_pc <= 32'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_pc <= 32'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_pc <= io_in_bits_pc;
    end else if (io_out_valid) begin
      executeBuffer_pc <= 32'h0;
    end
    if (reset) begin
      executeBuffer_inst <= 32'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_inst <= 32'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_inst <= io_in_bits_inst;
    end else if (io_out_valid) begin
      executeBuffer_inst <= 32'h0;
    end
    if (reset) begin
      executeBuffer_valid <= executeNop_valid;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_valid <= executeNop_valid;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_valid <= io_in_bits_valid;
    end else if (io_out_valid) begin
      executeBuffer_valid <= executeNop_valid;
    end
    if (reset) begin
      executeBuffer_bubble <= executeNop_bubble;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_bubble <= executeNop_bubble;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_bubble <= io_in_bits_bubble;
    end else if (io_out_valid) begin
      executeBuffer_bubble <= executeNop_bubble;
    end
    if (reset) begin
      executeBuffer_opcode_type <= executeNop_opcode_type;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_opcode_type <= executeNop_opcode_type;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_opcode_type <= io_in_bits_opcode_type;
    end else if (io_out_valid) begin
      executeBuffer_opcode_type <= executeNop_opcode_type;
    end
    if (reset) begin
      executeBuffer_opcode_func <= executeNop_opcode_func;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_opcode_func <= executeNop_opcode_func;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_opcode_func <= io_in_bits_opcode_func;
    end else if (io_out_valid) begin
      executeBuffer_opcode_func <= executeNop_opcode_func;
    end
    if (reset) begin
      executeBuffer_br_type <= 4'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_br_type <= 4'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_br_type <= io_in_bits_br_type;
    end else if (io_out_valid) begin
      executeBuffer_br_type <= 4'h0;
    end
    if (reset) begin
      executeBuffer_rf_en <= 1'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_rf_en <= 1'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_rf_en <= io_in_bits_rf_en;
    end else if (io_out_valid) begin
      executeBuffer_rf_en <= 1'h0;
    end
    if (reset) begin
      executeBuffer_wb_addr <= 5'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_wb_addr <= 5'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_wb_addr <= io_in_bits_wb_addr;
    end else if (io_out_valid) begin
      executeBuffer_wb_addr <= 5'h0;
    end
    if (reset) begin
      executeBuffer_wb_stage <= 2'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_wb_stage <= 2'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_wb_stage <= io_in_bits_wb_stage;
    end else if (io_out_valid) begin
      executeBuffer_wb_stage <= 2'h0;
    end
    if (reset) begin
      executeBuffer_op1_data <= 64'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_op1_data <= 64'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_op1_data <= io_in_bits_op1_data;
    end else if (io_out_valid) begin
      executeBuffer_op1_data <= 64'h0;
    end
    if (reset) begin
      executeBuffer_op2_data <= 64'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_op2_data <= 64'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_op2_data <= io_in_bits_op2_data;
    end else if (io_out_valid) begin
      executeBuffer_op2_data <= 64'h0;
    end
    if (reset) begin
      executeBuffer_rs1_data <= 64'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_rs1_data <= 64'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_rs1_data <= io_in_bits_rs1_data;
    end else if (io_out_valid) begin
      executeBuffer_rs1_data <= 64'h0;
    end
    if (reset) begin
      executeBuffer_rs2_data <= 64'h0;
    end else if (io_out_bits_redirect_valid) begin
      executeBuffer_rs2_data <= 64'h0;
    end else if (io_in_ready & ~io_flush & io_in_bits_valid) begin
      executeBuffer_rs2_data <= io_in_bits_rs2_data;
    end else if (io_out_valid) begin
      executeBuffer_rs2_data <= 64'h0;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  executeNop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  executeNop_bubble = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  executeNop_opcode_type = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  executeNop_opcode_func = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  executeBuffer_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  executeBuffer_inst = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  executeBuffer_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  executeBuffer_bubble = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  executeBuffer_opcode_type = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  executeBuffer_opcode_func = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  executeBuffer_br_type = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  executeBuffer_rf_en = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  executeBuffer_wb_addr = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  executeBuffer_wb_stage = _RAND_13[1:0];
  _RAND_14 = {2{`RANDOM}};
  executeBuffer_op1_data = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  executeBuffer_op2_data = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  executeBuffer_rs1_data = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  executeBuffer_rs2_data = _RAND_17[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_WriteBackUnit(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_valid,
  input         io_in_bits_wen,
  input  [4:0]  io_in_bits_wb_addr,
  input  [63:0] io_in_bits_wb_data,
  input         io_in_bits_redirect_valid,
  input  [31:0] io_in_bits_redirect_target,
  input         io_in_bits_flush,
  output [4:0]  io_regFile_w_addr,
  output [63:0] io_regFile_w_data,
  output        io_regFile_wen,
  output        io_bypass_rf_wen,
  output [4:0]  io_bypass_addr,
  output [63:0] io_bypass_data,
  output        io_redirect_valid,
  output [31:0] io_redirect_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif
  reg  writeBackBuffer_valid;
  reg  writeBackBuffer_wen;
  reg [4:0] writeBackBuffer_wb_addr;
  reg [63:0] writeBackBuffer_wb_data;
  reg  writeBackBuffer_redirect_valid;
  reg [31:0] writeBackBuffer_redirect_target;
  wire  _T = io_in_ready & io_in_valid;
  wire  _GEN_0 = _T & ~io_in_bits_flush & io_in_bits_valid;
  wire  _GEN_3 = _T & ~io_in_bits_flush & io_in_bits_wen;
  wire  _GEN_7 = _T & ~io_in_bits_flush & io_in_bits_redirect_valid;
  reg [63:0] instrCnt;
  wire [63:0] _instrCnt_T_1 = instrCnt + 64'h1;
  assign io_in_ready = 1'h1;
  assign io_regFile_w_addr = writeBackBuffer_wb_addr;
  assign io_regFile_w_data = writeBackBuffer_wb_data;
  assign io_regFile_wen = writeBackBuffer_valid & writeBackBuffer_wen;
  assign io_bypass_rf_wen = writeBackBuffer_wen;
  assign io_bypass_addr = writeBackBuffer_wb_addr;
  assign io_bypass_data = writeBackBuffer_wb_data;
  assign io_redirect_valid = writeBackBuffer_redirect_valid;
  assign io_redirect_target = writeBackBuffer_redirect_target;
  always @(posedge clock) begin
    if (reset) begin
      writeBackBuffer_valid <= 1'h0;
    end else begin
      writeBackBuffer_valid <= _GEN_0;
    end
    if (reset) begin
      writeBackBuffer_wen <= 1'h0;
    end else begin
      writeBackBuffer_wen <= _GEN_3;
    end
    if (reset) begin
      writeBackBuffer_wb_addr <= 5'h0;
    end else if (_T & ~io_in_bits_flush) begin
      writeBackBuffer_wb_addr <= io_in_bits_wb_addr;
    end else begin
      writeBackBuffer_wb_addr <= 5'h0;
    end
    if (reset) begin
      writeBackBuffer_wb_data <= 64'h0;
    end else if (_T & ~io_in_bits_flush) begin
      writeBackBuffer_wb_data <= io_in_bits_wb_data;
    end else begin
      writeBackBuffer_wb_data <= 64'h0;
    end
    if (reset) begin
      writeBackBuffer_redirect_valid <= 1'h0;
    end else begin
      writeBackBuffer_redirect_valid <= _GEN_7;
    end
    if (reset) begin
      writeBackBuffer_redirect_target <= 32'h0;
    end else if (_T & ~io_in_bits_flush) begin
      writeBackBuffer_redirect_target <= io_in_bits_redirect_target;
    end else begin
      writeBackBuffer_redirect_target <= 32'h0;
    end
    if (reset) begin
      instrCnt <= 64'h0;
    end else if (writeBackBuffer_valid) begin
      instrCnt <= _instrCnt_T_1;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeBackBuffer_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  writeBackBuffer_wen = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  writeBackBuffer_wb_addr = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  writeBackBuffer_wb_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  writeBackBuffer_redirect_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  writeBackBuffer_redirect_target = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  instrCnt = _RAND_6[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_r_rs1_addr,
  input  [4:0]  io_r_rs2_addr,
  output [63:0] io_r_rs1_data,
  output [63:0] io_r_rs2_data,
  input  [4:0]  io_w_w_addr,
  input  [63:0] io_w_w_data,
  input         io_w_wen
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif
  reg [63:0] regMem [0:31];
  wire  regMem_io_r_rs1_data_MPORT_en;
  wire [4:0] regMem_io_r_rs1_data_MPORT_addr;
  wire [63:0] regMem_io_r_rs1_data_MPORT_data;
  wire  regMem_io_r_rs2_data_MPORT_en;
  wire [4:0] regMem_io_r_rs2_data_MPORT_addr;
  wire [63:0] regMem_io_r_rs2_data_MPORT_data;
  wire [63:0] regMem_MPORT_data;
  wire [4:0] regMem_MPORT_addr;
  wire  regMem_MPORT_mask;
  wire  regMem_MPORT_en;
  wire [63:0] regMem_MPORT_1_data;
  wire [4:0] regMem_MPORT_1_addr;
  wire  regMem_MPORT_1_mask;
  wire  regMem_MPORT_1_en;
  wire [63:0] regMem_MPORT_2_data;
  wire [4:0] regMem_MPORT_2_addr;
  wire  regMem_MPORT_2_mask;
  wire  regMem_MPORT_2_en;
  wire [63:0] regMem_MPORT_3_data;
  wire [4:0] regMem_MPORT_3_addr;
  wire  regMem_MPORT_3_mask;
  wire  regMem_MPORT_3_en;
  wire [63:0] regMem_MPORT_4_data;
  wire [4:0] regMem_MPORT_4_addr;
  wire  regMem_MPORT_4_mask;
  wire  regMem_MPORT_4_en;
  wire [63:0] regMem_MPORT_5_data;
  wire [4:0] regMem_MPORT_5_addr;
  wire  regMem_MPORT_5_mask;
  wire  regMem_MPORT_5_en;
  wire [63:0] regMem_MPORT_6_data;
  wire [4:0] regMem_MPORT_6_addr;
  wire  regMem_MPORT_6_mask;
  wire  regMem_MPORT_6_en;
  wire [63:0] regMem_MPORT_7_data;
  wire [4:0] regMem_MPORT_7_addr;
  wire  regMem_MPORT_7_mask;
  wire  regMem_MPORT_7_en;
  wire [63:0] regMem_MPORT_8_data;
  wire [4:0] regMem_MPORT_8_addr;
  wire  regMem_MPORT_8_mask;
  wire  regMem_MPORT_8_en;
  wire [63:0] regMem_MPORT_9_data;
  wire [4:0] regMem_MPORT_9_addr;
  wire  regMem_MPORT_9_mask;
  wire  regMem_MPORT_9_en;
  wire [63:0] regMem_MPORT_10_data;
  wire [4:0] regMem_MPORT_10_addr;
  wire  regMem_MPORT_10_mask;
  wire  regMem_MPORT_10_en;
  wire [63:0] regMem_MPORT_11_data;
  wire [4:0] regMem_MPORT_11_addr;
  wire  regMem_MPORT_11_mask;
  wire  regMem_MPORT_11_en;
  wire [63:0] regMem_MPORT_12_data;
  wire [4:0] regMem_MPORT_12_addr;
  wire  regMem_MPORT_12_mask;
  wire  regMem_MPORT_12_en;
  wire [63:0] regMem_MPORT_13_data;
  wire [4:0] regMem_MPORT_13_addr;
  wire  regMem_MPORT_13_mask;
  wire  regMem_MPORT_13_en;
  wire [63:0] regMem_MPORT_14_data;
  wire [4:0] regMem_MPORT_14_addr;
  wire  regMem_MPORT_14_mask;
  wire  regMem_MPORT_14_en;
  wire [63:0] regMem_MPORT_15_data;
  wire [4:0] regMem_MPORT_15_addr;
  wire  regMem_MPORT_15_mask;
  wire  regMem_MPORT_15_en;
  wire [63:0] regMem_MPORT_16_data;
  wire [4:0] regMem_MPORT_16_addr;
  wire  regMem_MPORT_16_mask;
  wire  regMem_MPORT_16_en;
  wire [63:0] regMem_MPORT_17_data;
  wire [4:0] regMem_MPORT_17_addr;
  wire  regMem_MPORT_17_mask;
  wire  regMem_MPORT_17_en;
  wire [63:0] regMem_MPORT_18_data;
  wire [4:0] regMem_MPORT_18_addr;
  wire  regMem_MPORT_18_mask;
  wire  regMem_MPORT_18_en;
  wire [63:0] regMem_MPORT_19_data;
  wire [4:0] regMem_MPORT_19_addr;
  wire  regMem_MPORT_19_mask;
  wire  regMem_MPORT_19_en;
  wire [63:0] regMem_MPORT_20_data;
  wire [4:0] regMem_MPORT_20_addr;
  wire  regMem_MPORT_20_mask;
  wire  regMem_MPORT_20_en;
  wire [63:0] regMem_MPORT_21_data;
  wire [4:0] regMem_MPORT_21_addr;
  wire  regMem_MPORT_21_mask;
  wire  regMem_MPORT_21_en;
  wire [63:0] regMem_MPORT_22_data;
  wire [4:0] regMem_MPORT_22_addr;
  wire  regMem_MPORT_22_mask;
  wire  regMem_MPORT_22_en;
  wire [63:0] regMem_MPORT_23_data;
  wire [4:0] regMem_MPORT_23_addr;
  wire  regMem_MPORT_23_mask;
  wire  regMem_MPORT_23_en;
  wire [63:0] regMem_MPORT_24_data;
  wire [4:0] regMem_MPORT_24_addr;
  wire  regMem_MPORT_24_mask;
  wire  regMem_MPORT_24_en;
  wire [63:0] regMem_MPORT_25_data;
  wire [4:0] regMem_MPORT_25_addr;
  wire  regMem_MPORT_25_mask;
  wire  regMem_MPORT_25_en;
  wire [63:0] regMem_MPORT_26_data;
  wire [4:0] regMem_MPORT_26_addr;
  wire  regMem_MPORT_26_mask;
  wire  regMem_MPORT_26_en;
  wire [63:0] regMem_MPORT_27_data;
  wire [4:0] regMem_MPORT_27_addr;
  wire  regMem_MPORT_27_mask;
  wire  regMem_MPORT_27_en;
  wire [63:0] regMem_MPORT_28_data;
  wire [4:0] regMem_MPORT_28_addr;
  wire  regMem_MPORT_28_mask;
  wire  regMem_MPORT_28_en;
  wire [63:0] regMem_MPORT_29_data;
  wire [4:0] regMem_MPORT_29_addr;
  wire  regMem_MPORT_29_mask;
  wire  regMem_MPORT_29_en;
  wire [63:0] regMem_MPORT_30_data;
  wire [4:0] regMem_MPORT_30_addr;
  wire  regMem_MPORT_30_mask;
  wire  regMem_MPORT_30_en;
  wire [63:0] regMem_MPORT_31_data;
  wire [4:0] regMem_MPORT_31_addr;
  wire  regMem_MPORT_31_mask;
  wire  regMem_MPORT_31_en;
  wire [63:0] regMem_MPORT_32_data;
  wire [4:0] regMem_MPORT_32_addr;
  wire  regMem_MPORT_32_mask;
  wire  regMem_MPORT_32_en;
  wire  _T = io_w_w_addr >= 5'h1;
  assign regMem_io_r_rs1_data_MPORT_en = 1'h1;
  assign regMem_io_r_rs1_data_MPORT_addr = io_r_rs1_addr;
  assign regMem_io_r_rs1_data_MPORT_data = regMem[regMem_io_r_rs1_data_MPORT_addr];
  assign regMem_io_r_rs2_data_MPORT_en = 1'h1;
  assign regMem_io_r_rs2_data_MPORT_addr = io_r_rs2_addr;
  assign regMem_io_r_rs2_data_MPORT_data = regMem[regMem_io_r_rs2_data_MPORT_addr];
  assign regMem_MPORT_data = io_w_w_data;
  assign regMem_MPORT_addr = io_w_w_addr;
  assign regMem_MPORT_mask = 1'h1;
  assign regMem_MPORT_en = io_w_wen & _T;
  assign regMem_MPORT_1_data = 64'h0;
  assign regMem_MPORT_1_addr = 5'h0;
  assign regMem_MPORT_1_mask = 1'h1;
  assign regMem_MPORT_1_en = reset;
  assign regMem_MPORT_2_data = 64'h0;
  assign regMem_MPORT_2_addr = 5'h1;
  assign regMem_MPORT_2_mask = 1'h1;
  assign regMem_MPORT_2_en = reset;
  assign regMem_MPORT_3_data = 64'h0;
  assign regMem_MPORT_3_addr = 5'h2;
  assign regMem_MPORT_3_mask = 1'h1;
  assign regMem_MPORT_3_en = reset;
  assign regMem_MPORT_4_data = 64'h0;
  assign regMem_MPORT_4_addr = 5'h3;
  assign regMem_MPORT_4_mask = 1'h1;
  assign regMem_MPORT_4_en = reset;
  assign regMem_MPORT_5_data = 64'h0;
  assign regMem_MPORT_5_addr = 5'h4;
  assign regMem_MPORT_5_mask = 1'h1;
  assign regMem_MPORT_5_en = reset;
  assign regMem_MPORT_6_data = 64'h0;
  assign regMem_MPORT_6_addr = 5'h5;
  assign regMem_MPORT_6_mask = 1'h1;
  assign regMem_MPORT_6_en = reset;
  assign regMem_MPORT_7_data = 64'h0;
  assign regMem_MPORT_7_addr = 5'h6;
  assign regMem_MPORT_7_mask = 1'h1;
  assign regMem_MPORT_7_en = reset;
  assign regMem_MPORT_8_data = 64'h0;
  assign regMem_MPORT_8_addr = 5'h7;
  assign regMem_MPORT_8_mask = 1'h1;
  assign regMem_MPORT_8_en = reset;
  assign regMem_MPORT_9_data = 64'h0;
  assign regMem_MPORT_9_addr = 5'h8;
  assign regMem_MPORT_9_mask = 1'h1;
  assign regMem_MPORT_9_en = reset;
  assign regMem_MPORT_10_data = 64'h0;
  assign regMem_MPORT_10_addr = 5'h9;
  assign regMem_MPORT_10_mask = 1'h1;
  assign regMem_MPORT_10_en = reset;
  assign regMem_MPORT_11_data = 64'h0;
  assign regMem_MPORT_11_addr = 5'ha;
  assign regMem_MPORT_11_mask = 1'h1;
  assign regMem_MPORT_11_en = reset;
  assign regMem_MPORT_12_data = 64'h0;
  assign regMem_MPORT_12_addr = 5'hb;
  assign regMem_MPORT_12_mask = 1'h1;
  assign regMem_MPORT_12_en = reset;
  assign regMem_MPORT_13_data = 64'h0;
  assign regMem_MPORT_13_addr = 5'hc;
  assign regMem_MPORT_13_mask = 1'h1;
  assign regMem_MPORT_13_en = reset;
  assign regMem_MPORT_14_data = 64'h0;
  assign regMem_MPORT_14_addr = 5'hd;
  assign regMem_MPORT_14_mask = 1'h1;
  assign regMem_MPORT_14_en = reset;
  assign regMem_MPORT_15_data = 64'h0;
  assign regMem_MPORT_15_addr = 5'he;
  assign regMem_MPORT_15_mask = 1'h1;
  assign regMem_MPORT_15_en = reset;
  assign regMem_MPORT_16_data = 64'h0;
  assign regMem_MPORT_16_addr = 5'hf;
  assign regMem_MPORT_16_mask = 1'h1;
  assign regMem_MPORT_16_en = reset;
  assign regMem_MPORT_17_data = 64'h0;
  assign regMem_MPORT_17_addr = 5'h10;
  assign regMem_MPORT_17_mask = 1'h1;
  assign regMem_MPORT_17_en = reset;
  assign regMem_MPORT_18_data = 64'h0;
  assign regMem_MPORT_18_addr = 5'h11;
  assign regMem_MPORT_18_mask = 1'h1;
  assign regMem_MPORT_18_en = reset;
  assign regMem_MPORT_19_data = 64'h0;
  assign regMem_MPORT_19_addr = 5'h12;
  assign regMem_MPORT_19_mask = 1'h1;
  assign regMem_MPORT_19_en = reset;
  assign regMem_MPORT_20_data = 64'h0;
  assign regMem_MPORT_20_addr = 5'h13;
  assign regMem_MPORT_20_mask = 1'h1;
  assign regMem_MPORT_20_en = reset;
  assign regMem_MPORT_21_data = 64'h0;
  assign regMem_MPORT_21_addr = 5'h14;
  assign regMem_MPORT_21_mask = 1'h1;
  assign regMem_MPORT_21_en = reset;
  assign regMem_MPORT_22_data = 64'h0;
  assign regMem_MPORT_22_addr = 5'h15;
  assign regMem_MPORT_22_mask = 1'h1;
  assign regMem_MPORT_22_en = reset;
  assign regMem_MPORT_23_data = 64'h0;
  assign regMem_MPORT_23_addr = 5'h16;
  assign regMem_MPORT_23_mask = 1'h1;
  assign regMem_MPORT_23_en = reset;
  assign regMem_MPORT_24_data = 64'h0;
  assign regMem_MPORT_24_addr = 5'h17;
  assign regMem_MPORT_24_mask = 1'h1;
  assign regMem_MPORT_24_en = reset;
  assign regMem_MPORT_25_data = 64'h0;
  assign regMem_MPORT_25_addr = 5'h18;
  assign regMem_MPORT_25_mask = 1'h1;
  assign regMem_MPORT_25_en = reset;
  assign regMem_MPORT_26_data = 64'h0;
  assign regMem_MPORT_26_addr = 5'h19;
  assign regMem_MPORT_26_mask = 1'h1;
  assign regMem_MPORT_26_en = reset;
  assign regMem_MPORT_27_data = 64'h0;
  assign regMem_MPORT_27_addr = 5'h1a;
  assign regMem_MPORT_27_mask = 1'h1;
  assign regMem_MPORT_27_en = reset;
  assign regMem_MPORT_28_data = 64'h0;
  assign regMem_MPORT_28_addr = 5'h1b;
  assign regMem_MPORT_28_mask = 1'h1;
  assign regMem_MPORT_28_en = reset;
  assign regMem_MPORT_29_data = 64'h0;
  assign regMem_MPORT_29_addr = 5'h1c;
  assign regMem_MPORT_29_mask = 1'h1;
  assign regMem_MPORT_29_en = reset;
  assign regMem_MPORT_30_data = 64'h0;
  assign regMem_MPORT_30_addr = 5'h1d;
  assign regMem_MPORT_30_mask = 1'h1;
  assign regMem_MPORT_30_en = reset;
  assign regMem_MPORT_31_data = 64'h0;
  assign regMem_MPORT_31_addr = 5'h1e;
  assign regMem_MPORT_31_mask = 1'h1;
  assign regMem_MPORT_31_en = reset;
  assign regMem_MPORT_32_data = 64'h0;
  assign regMem_MPORT_32_addr = 5'h1f;
  assign regMem_MPORT_32_mask = 1'h1;
  assign regMem_MPORT_32_en = reset;
  assign io_r_rs1_data = io_r_rs1_addr != 5'h0 ? regMem_io_r_rs1_data_MPORT_data : 64'h0;
  assign io_r_rs2_data = io_r_rs2_addr != 5'h0 ? regMem_io_r_rs2_data_MPORT_data : 64'h0;
  always @(posedge clock) begin
    if (regMem_MPORT_en & regMem_MPORT_mask) begin
      regMem[regMem_MPORT_addr] <= regMem_MPORT_data;
    end
    if (regMem_MPORT_1_en & regMem_MPORT_1_mask) begin
      regMem[regMem_MPORT_1_addr] <= regMem_MPORT_1_data;
    end
    if (regMem_MPORT_2_en & regMem_MPORT_2_mask) begin
      regMem[regMem_MPORT_2_addr] <= regMem_MPORT_2_data;
    end
    if (regMem_MPORT_3_en & regMem_MPORT_3_mask) begin
      regMem[regMem_MPORT_3_addr] <= regMem_MPORT_3_data;
    end
    if (regMem_MPORT_4_en & regMem_MPORT_4_mask) begin
      regMem[regMem_MPORT_4_addr] <= regMem_MPORT_4_data;
    end
    if (regMem_MPORT_5_en & regMem_MPORT_5_mask) begin
      regMem[regMem_MPORT_5_addr] <= regMem_MPORT_5_data;
    end
    if (regMem_MPORT_6_en & regMem_MPORT_6_mask) begin
      regMem[regMem_MPORT_6_addr] <= regMem_MPORT_6_data;
    end
    if (regMem_MPORT_7_en & regMem_MPORT_7_mask) begin
      regMem[regMem_MPORT_7_addr] <= regMem_MPORT_7_data;
    end
    if (regMem_MPORT_8_en & regMem_MPORT_8_mask) begin
      regMem[regMem_MPORT_8_addr] <= regMem_MPORT_8_data;
    end
    if (regMem_MPORT_9_en & regMem_MPORT_9_mask) begin
      regMem[regMem_MPORT_9_addr] <= regMem_MPORT_9_data;
    end
    if (regMem_MPORT_10_en & regMem_MPORT_10_mask) begin
      regMem[regMem_MPORT_10_addr] <= regMem_MPORT_10_data;
    end
    if (regMem_MPORT_11_en & regMem_MPORT_11_mask) begin
      regMem[regMem_MPORT_11_addr] <= regMem_MPORT_11_data;
    end
    if (regMem_MPORT_12_en & regMem_MPORT_12_mask) begin
      regMem[regMem_MPORT_12_addr] <= regMem_MPORT_12_data;
    end
    if (regMem_MPORT_13_en & regMem_MPORT_13_mask) begin
      regMem[regMem_MPORT_13_addr] <= regMem_MPORT_13_data;
    end
    if (regMem_MPORT_14_en & regMem_MPORT_14_mask) begin
      regMem[regMem_MPORT_14_addr] <= regMem_MPORT_14_data;
    end
    if (regMem_MPORT_15_en & regMem_MPORT_15_mask) begin
      regMem[regMem_MPORT_15_addr] <= regMem_MPORT_15_data;
    end
    if (regMem_MPORT_16_en & regMem_MPORT_16_mask) begin
      regMem[regMem_MPORT_16_addr] <= regMem_MPORT_16_data;
    end
    if (regMem_MPORT_17_en & regMem_MPORT_17_mask) begin
      regMem[regMem_MPORT_17_addr] <= regMem_MPORT_17_data;
    end
    if (regMem_MPORT_18_en & regMem_MPORT_18_mask) begin
      regMem[regMem_MPORT_18_addr] <= regMem_MPORT_18_data;
    end
    if (regMem_MPORT_19_en & regMem_MPORT_19_mask) begin
      regMem[regMem_MPORT_19_addr] <= regMem_MPORT_19_data;
    end
    if (regMem_MPORT_20_en & regMem_MPORT_20_mask) begin
      regMem[regMem_MPORT_20_addr] <= regMem_MPORT_20_data;
    end
    if (regMem_MPORT_21_en & regMem_MPORT_21_mask) begin
      regMem[regMem_MPORT_21_addr] <= regMem_MPORT_21_data;
    end
    if (regMem_MPORT_22_en & regMem_MPORT_22_mask) begin
      regMem[regMem_MPORT_22_addr] <= regMem_MPORT_22_data;
    end
    if (regMem_MPORT_23_en & regMem_MPORT_23_mask) begin
      regMem[regMem_MPORT_23_addr] <= regMem_MPORT_23_data;
    end
    if (regMem_MPORT_24_en & regMem_MPORT_24_mask) begin
      regMem[regMem_MPORT_24_addr] <= regMem_MPORT_24_data;
    end
    if (regMem_MPORT_25_en & regMem_MPORT_25_mask) begin
      regMem[regMem_MPORT_25_addr] <= regMem_MPORT_25_data;
    end
    if (regMem_MPORT_26_en & regMem_MPORT_26_mask) begin
      regMem[regMem_MPORT_26_addr] <= regMem_MPORT_26_data;
    end
    if (regMem_MPORT_27_en & regMem_MPORT_27_mask) begin
      regMem[regMem_MPORT_27_addr] <= regMem_MPORT_27_data;
    end
    if (regMem_MPORT_28_en & regMem_MPORT_28_mask) begin
      regMem[regMem_MPORT_28_addr] <= regMem_MPORT_28_data;
    end
    if (regMem_MPORT_29_en & regMem_MPORT_29_mask) begin
      regMem[regMem_MPORT_29_addr] <= regMem_MPORT_29_data;
    end
    if (regMem_MPORT_30_en & regMem_MPORT_30_mask) begin
      regMem[regMem_MPORT_30_addr] <= regMem_MPORT_30_data;
    end
    if (regMem_MPORT_31_en & regMem_MPORT_31_mask) begin
      regMem[regMem_MPORT_31_addr] <= regMem_MPORT_31_data;
    end
    if (regMem_MPORT_32_en & regMem_MPORT_32_mask) begin
      regMem[regMem_MPORT_32_addr] <= regMem_MPORT_32_data;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regMem[initvar] = _RAND_0[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Pipeline(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_inst,
  input  [31:0] io_in_bits_pc,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [1:0]  io_dmem_req_bits_size,
  output [2:0]  io_dmem_req_bits_cmd,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [63:0] io_mmio_req_bits_wdata,
  output [1:0]  io_mmio_req_bits_size,
  output [2:0]  io_mmio_req_bits_cmd,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_redirect_valid,
  output [31:0] io_redirect_target,
  output        flushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif
  wire  decodeStage_clock;
  wire  decodeStage_reset;
  wire  decodeStage_io_flush;
  wire  decodeStage_io_in_ready;
  wire  decodeStage_io_in_valid;
  wire [31:0] decodeStage_io_in_bits_inst;
  wire [31:0] decodeStage_io_in_bits_pc;
  wire  decodeStage_io_out_ready;
  wire  decodeStage_io_out_valid;
  wire [31:0] decodeStage_io_out_bits_pc;
  wire [31:0] decodeStage_io_out_bits_inst;
  wire  decodeStage_io_out_bits_valid;
  wire  decodeStage_io_out_bits_bubble;
  wire [2:0] decodeStage_io_out_bits_opcode_type;
  wire [5:0] decodeStage_io_out_bits_opcode_func;
  wire [3:0] decodeStage_io_out_bits_br_type;
  wire  decodeStage_io_out_bits_rf_en;
  wire [4:0] decodeStage_io_out_bits_wb_addr;
  wire [1:0] decodeStage_io_out_bits_wb_stage;
  wire [63:0] decodeStage_io_out_bits_op1_data;
  wire [63:0] decodeStage_io_out_bits_op2_data;
  wire [63:0] decodeStage_io_out_bits_rs1_data;
  wire [63:0] decodeStage_io_out_bits_rs2_data;
  wire [4:0] decodeStage_io_regFile_rs1_addr;
  wire [4:0] decodeStage_io_regFile_rs2_addr;
  wire [63:0] decodeStage_io_regFile_rs1_data;
  wire [63:0] decodeStage_io_regFile_rs2_data;
  wire  decodeStage_io_bypass_0_rf_wen;
  wire [4:0] decodeStage_io_bypass_0_addr;
  wire [63:0] decodeStage_io_bypass_0_data;
  wire  decodeStage_io_bypass_1_rf_wen;
  wire [4:0] decodeStage_io_bypass_1_addr;
  wire [63:0] decodeStage_io_bypass_1_data;
  wire  executeStage_clock;
  wire  executeStage_reset;
  wire  executeStage_io_flush;
  wire  executeStage_io_in_ready;
  wire  executeStage_io_in_valid;
  wire [31:0] executeStage_io_in_bits_pc;
  wire [31:0] executeStage_io_in_bits_inst;
  wire  executeStage_io_in_bits_valid;
  wire  executeStage_io_in_bits_bubble;
  wire [2:0] executeStage_io_in_bits_opcode_type;
  wire [5:0] executeStage_io_in_bits_opcode_func;
  wire [3:0] executeStage_io_in_bits_br_type;
  wire  executeStage_io_in_bits_rf_en;
  wire [4:0] executeStage_io_in_bits_wb_addr;
  wire [1:0] executeStage_io_in_bits_wb_stage;
  wire [63:0] executeStage_io_in_bits_op1_data;
  wire [63:0] executeStage_io_in_bits_op2_data;
  wire [63:0] executeStage_io_in_bits_rs1_data;
  wire [63:0] executeStage_io_in_bits_rs2_data;
  wire  executeStage_io_dmem_req_ready;
  wire  executeStage_io_dmem_req_valid;
  wire [31:0] executeStage_io_dmem_req_bits_addr;
  wire [63:0] executeStage_io_dmem_req_bits_wdata;
  wire [1:0] executeStage_io_dmem_req_bits_size;
  wire [2:0] executeStage_io_dmem_req_bits_cmd;
  wire  executeStage_io_dmem_resp_valid;
  wire [63:0] executeStage_io_dmem_resp_bits_rdata;
  wire  executeStage_io_mmio_req_ready;
  wire  executeStage_io_mmio_req_valid;
  wire [31:0] executeStage_io_mmio_req_bits_addr;
  wire [63:0] executeStage_io_mmio_req_bits_wdata;
  wire [1:0] executeStage_io_mmio_req_bits_size;
  wire [2:0] executeStage_io_mmio_req_bits_cmd;
  wire  executeStage_io_mmio_resp_valid;
  wire [63:0] executeStage_io_mmio_resp_bits_rdata;
  wire  executeStage_io_out_ready;
  wire  executeStage_io_out_valid;
  wire  executeStage_io_out_bits_valid;
  wire  executeStage_io_out_bits_wen;
  wire [4:0] executeStage_io_out_bits_wb_addr;
  wire [63:0] executeStage_io_out_bits_wb_data;
  wire  executeStage_io_out_bits_redirect_valid;
  wire [31:0] executeStage_io_out_bits_redirect_target;
  wire  executeStage_io_bypass_rf_wen;
  wire [4:0] executeStage_io_bypass_addr;
  wire [63:0] executeStage_io_bypass_data;
  wire  executeStage_flushICache;
  wire  writeBackUnit_clock;
  wire  writeBackUnit_reset;
  wire  writeBackUnit_io_in_ready;
  wire  writeBackUnit_io_in_valid;
  wire  writeBackUnit_io_in_bits_valid;
  wire  writeBackUnit_io_in_bits_wen;
  wire [4:0] writeBackUnit_io_in_bits_wb_addr;
  wire [63:0] writeBackUnit_io_in_bits_wb_data;
  wire  writeBackUnit_io_in_bits_redirect_valid;
  wire [31:0] writeBackUnit_io_in_bits_redirect_target;
  wire  writeBackUnit_io_in_bits_flush;
  wire [4:0] writeBackUnit_io_regFile_w_addr;
  wire [63:0] writeBackUnit_io_regFile_w_data;
  wire  writeBackUnit_io_regFile_wen;
  wire  writeBackUnit_io_bypass_rf_wen;
  wire [4:0] writeBackUnit_io_bypass_addr;
  wire [63:0] writeBackUnit_io_bypass_data;
  wire  writeBackUnit_io_redirect_valid;
  wire [31:0] writeBackUnit_io_redirect_target;
  wire  regFile_clock;
  wire  regFile_reset;
  wire [4:0] regFile_io_r_rs1_addr;
  wire [4:0] regFile_io_r_rs2_addr;
  wire [63:0] regFile_io_r_rs1_data;
  wire [63:0] regFile_io_r_rs2_data;
  wire [4:0] regFile_io_w_w_addr;
  wire [63:0] regFile_io_w_w_data;
  wire  regFile_io_w_wen;
  wire  _T = executeStage_io_in_ready & executeStage_io_in_valid;
  wire  _T_1 = executeStage_io_out_ready & executeStage_io_out_valid;
  wire  _T_4 = _T & _T_1 & ~writeBackUnit_io_redirect_valid;
  wire  _T_9 = ~_T & _T_1 | writeBackUnit_io_redirect_valid;
  reg [31:0] pipelineRegs_pc;
  reg [31:0] pipelineRegs_inst;
  reg  pipelineRegs_valid;
  reg  pipelineRegs_bubble;
  reg [2:0] pipelineRegs_opcode_type;
  reg [5:0] pipelineRegs_opcode_func;
  reg [3:0] pipelineRegs_br_type;
  reg  pipelineRegs_rf_en;
  reg [4:0] pipelineRegs_wb_addr;
  reg [1:0] pipelineRegs_wb_stage;
  reg [63:0] pipelineRegs_op1_data;
  reg [63:0] pipelineRegs_op2_data;
  reg [63:0] pipelineRegs_rs1_data;
  reg [63:0] pipelineRegs_rs2_data;
  ysyx_040656_DecodeStage decodeStage (
    .clock(decodeStage_clock),
    .reset(decodeStage_reset),
    .io_flush(decodeStage_io_flush),
    .io_in_ready(decodeStage_io_in_ready),
    .io_in_valid(decodeStage_io_in_valid),
    .io_in_bits_inst(decodeStage_io_in_bits_inst),
    .io_in_bits_pc(decodeStage_io_in_bits_pc),
    .io_out_ready(decodeStage_io_out_ready),
    .io_out_valid(decodeStage_io_out_valid),
    .io_out_bits_pc(decodeStage_io_out_bits_pc),
    .io_out_bits_inst(decodeStage_io_out_bits_inst),
    .io_out_bits_valid(decodeStage_io_out_bits_valid),
    .io_out_bits_bubble(decodeStage_io_out_bits_bubble),
    .io_out_bits_opcode_type(decodeStage_io_out_bits_opcode_type),
    .io_out_bits_opcode_func(decodeStage_io_out_bits_opcode_func),
    .io_out_bits_br_type(decodeStage_io_out_bits_br_type),
    .io_out_bits_rf_en(decodeStage_io_out_bits_rf_en),
    .io_out_bits_wb_addr(decodeStage_io_out_bits_wb_addr),
    .io_out_bits_wb_stage(decodeStage_io_out_bits_wb_stage),
    .io_out_bits_op1_data(decodeStage_io_out_bits_op1_data),
    .io_out_bits_op2_data(decodeStage_io_out_bits_op2_data),
    .io_out_bits_rs1_data(decodeStage_io_out_bits_rs1_data),
    .io_out_bits_rs2_data(decodeStage_io_out_bits_rs2_data),
    .io_regFile_rs1_addr(decodeStage_io_regFile_rs1_addr),
    .io_regFile_rs2_addr(decodeStage_io_regFile_rs2_addr),
    .io_regFile_rs1_data(decodeStage_io_regFile_rs1_data),
    .io_regFile_rs2_data(decodeStage_io_regFile_rs2_data),
    .io_bypass_0_rf_wen(decodeStage_io_bypass_0_rf_wen),
    .io_bypass_0_addr(decodeStage_io_bypass_0_addr),
    .io_bypass_0_data(decodeStage_io_bypass_0_data),
    .io_bypass_1_rf_wen(decodeStage_io_bypass_1_rf_wen),
    .io_bypass_1_addr(decodeStage_io_bypass_1_addr),
    .io_bypass_1_data(decodeStage_io_bypass_1_data)
  );
  ysyx_040656_ExecuteStage executeStage (
    .clock(executeStage_clock),
    .reset(executeStage_reset),
    .io_flush(executeStage_io_flush),
    .io_in_ready(executeStage_io_in_ready),
    .io_in_valid(executeStage_io_in_valid),
    .io_in_bits_pc(executeStage_io_in_bits_pc),
    .io_in_bits_inst(executeStage_io_in_bits_inst),
    .io_in_bits_valid(executeStage_io_in_bits_valid),
    .io_in_bits_bubble(executeStage_io_in_bits_bubble),
    .io_in_bits_opcode_type(executeStage_io_in_bits_opcode_type),
    .io_in_bits_opcode_func(executeStage_io_in_bits_opcode_func),
    .io_in_bits_br_type(executeStage_io_in_bits_br_type),
    .io_in_bits_rf_en(executeStage_io_in_bits_rf_en),
    .io_in_bits_wb_addr(executeStage_io_in_bits_wb_addr),
    .io_in_bits_wb_stage(executeStage_io_in_bits_wb_stage),
    .io_in_bits_op1_data(executeStage_io_in_bits_op1_data),
    .io_in_bits_op2_data(executeStage_io_in_bits_op2_data),
    .io_in_bits_rs1_data(executeStage_io_in_bits_rs1_data),
    .io_in_bits_rs2_data(executeStage_io_in_bits_rs2_data),
    .io_dmem_req_ready(executeStage_io_dmem_req_ready),
    .io_dmem_req_valid(executeStage_io_dmem_req_valid),
    .io_dmem_req_bits_addr(executeStage_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(executeStage_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_size(executeStage_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(executeStage_io_dmem_req_bits_cmd),
    .io_dmem_resp_valid(executeStage_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(executeStage_io_dmem_resp_bits_rdata),
    .io_mmio_req_ready(executeStage_io_mmio_req_ready),
    .io_mmio_req_valid(executeStage_io_mmio_req_valid),
    .io_mmio_req_bits_addr(executeStage_io_mmio_req_bits_addr),
    .io_mmio_req_bits_wdata(executeStage_io_mmio_req_bits_wdata),
    .io_mmio_req_bits_size(executeStage_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(executeStage_io_mmio_req_bits_cmd),
    .io_mmio_resp_valid(executeStage_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(executeStage_io_mmio_resp_bits_rdata),
    .io_out_ready(executeStage_io_out_ready),
    .io_out_valid(executeStage_io_out_valid),
    .io_out_bits_valid(executeStage_io_out_bits_valid),
    .io_out_bits_wen(executeStage_io_out_bits_wen),
    .io_out_bits_wb_addr(executeStage_io_out_bits_wb_addr),
    .io_out_bits_wb_data(executeStage_io_out_bits_wb_data),
    .io_out_bits_redirect_valid(executeStage_io_out_bits_redirect_valid),
    .io_out_bits_redirect_target(executeStage_io_out_bits_redirect_target),
    .io_bypass_rf_wen(executeStage_io_bypass_rf_wen),
    .io_bypass_addr(executeStage_io_bypass_addr),
    .io_bypass_data(executeStage_io_bypass_data),
    .flushICache(executeStage_flushICache)
  );
  ysyx_040656_WriteBackUnit writeBackUnit (
    .clock(writeBackUnit_clock),
    .reset(writeBackUnit_reset),
    .io_in_ready(writeBackUnit_io_in_ready),
    .io_in_valid(writeBackUnit_io_in_valid),
    .io_in_bits_valid(writeBackUnit_io_in_bits_valid),
    .io_in_bits_wen(writeBackUnit_io_in_bits_wen),
    .io_in_bits_wb_addr(writeBackUnit_io_in_bits_wb_addr),
    .io_in_bits_wb_data(writeBackUnit_io_in_bits_wb_data),
    .io_in_bits_redirect_valid(writeBackUnit_io_in_bits_redirect_valid),
    .io_in_bits_redirect_target(writeBackUnit_io_in_bits_redirect_target),
    .io_in_bits_flush(writeBackUnit_io_in_bits_flush),
    .io_regFile_w_addr(writeBackUnit_io_regFile_w_addr),
    .io_regFile_w_data(writeBackUnit_io_regFile_w_data),
    .io_regFile_wen(writeBackUnit_io_regFile_wen),
    .io_bypass_rf_wen(writeBackUnit_io_bypass_rf_wen),
    .io_bypass_addr(writeBackUnit_io_bypass_addr),
    .io_bypass_data(writeBackUnit_io_bypass_data),
    .io_redirect_valid(writeBackUnit_io_redirect_valid),
    .io_redirect_target(writeBackUnit_io_redirect_target)
  );
  ysyx_040656_RegFile regFile (
    .clock(regFile_clock),
    .reset(regFile_reset),
    .io_r_rs1_addr(regFile_io_r_rs1_addr),
    .io_r_rs2_addr(regFile_io_r_rs2_addr),
    .io_r_rs1_data(regFile_io_r_rs1_data),
    .io_r_rs2_data(regFile_io_r_rs2_data),
    .io_w_w_addr(regFile_io_w_w_addr),
    .io_w_w_data(regFile_io_w_w_data),
    .io_w_wen(regFile_io_w_wen)
  );
  assign io_in_ready = decodeStage_io_in_ready;
  assign io_dmem_req_valid = executeStage_io_dmem_req_valid;
  assign io_dmem_req_bits_addr = executeStage_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_wdata = executeStage_io_dmem_req_bits_wdata;
  assign io_dmem_req_bits_size = executeStage_io_dmem_req_bits_size;
  assign io_dmem_req_bits_cmd = executeStage_io_dmem_req_bits_cmd;
  assign io_mmio_req_valid = executeStage_io_mmio_req_valid;
  assign io_mmio_req_bits_addr = executeStage_io_mmio_req_bits_addr;
  assign io_mmio_req_bits_wdata = executeStage_io_mmio_req_bits_wdata;
  assign io_mmio_req_bits_size = executeStage_io_mmio_req_bits_size;
  assign io_mmio_req_bits_cmd = executeStage_io_mmio_req_bits_cmd;
  assign io_redirect_valid = writeBackUnit_io_redirect_valid;
  assign io_redirect_target = writeBackUnit_io_redirect_target;
  assign flushICache = executeStage_flushICache;
  assign decodeStage_clock = clock;
  assign decodeStage_reset = reset;
  assign decodeStage_io_flush = writeBackUnit_io_redirect_valid;
  assign decodeStage_io_in_valid = io_in_valid;
  assign decodeStage_io_in_bits_inst = io_in_bits_inst;
  assign decodeStage_io_in_bits_pc = io_in_bits_pc;
  assign decodeStage_io_out_ready = executeStage_io_in_ready;
  assign decodeStage_io_regFile_rs1_data = regFile_io_r_rs1_data;
  assign decodeStage_io_regFile_rs2_data = regFile_io_r_rs2_data;
  assign decodeStage_io_bypass_0_rf_wen = executeStage_io_bypass_rf_wen;
  assign decodeStage_io_bypass_0_addr = executeStage_io_bypass_addr;
  assign decodeStage_io_bypass_0_data = executeStage_io_bypass_data;
  assign decodeStage_io_bypass_1_rf_wen = writeBackUnit_io_bypass_rf_wen;
  assign decodeStage_io_bypass_1_addr = writeBackUnit_io_bypass_addr;
  assign decodeStage_io_bypass_1_data = writeBackUnit_io_bypass_data;
  assign executeStage_clock = clock;
  assign executeStage_reset = reset;
  assign executeStage_io_flush = writeBackUnit_io_redirect_valid;
  assign executeStage_io_in_valid = 1'h1;
  assign executeStage_io_in_bits_pc = pipelineRegs_pc;
  assign executeStage_io_in_bits_inst = pipelineRegs_inst;
  assign executeStage_io_in_bits_valid = pipelineRegs_valid;
  assign executeStage_io_in_bits_bubble = pipelineRegs_bubble;
  assign executeStage_io_in_bits_opcode_type = pipelineRegs_opcode_type;
  assign executeStage_io_in_bits_opcode_func = pipelineRegs_opcode_func;
  assign executeStage_io_in_bits_br_type = pipelineRegs_br_type;
  assign executeStage_io_in_bits_rf_en = pipelineRegs_rf_en;
  assign executeStage_io_in_bits_wb_addr = pipelineRegs_wb_addr;
  assign executeStage_io_in_bits_wb_stage = pipelineRegs_wb_stage;
  assign executeStage_io_in_bits_op1_data = pipelineRegs_op1_data;
  assign executeStage_io_in_bits_op2_data = pipelineRegs_op2_data;
  assign executeStage_io_in_bits_rs1_data = pipelineRegs_rs1_data;
  assign executeStage_io_in_bits_rs2_data = pipelineRegs_rs2_data;
  assign executeStage_io_dmem_req_ready = io_dmem_req_ready;
  assign executeStage_io_dmem_resp_valid = io_dmem_resp_valid;
  assign executeStage_io_dmem_resp_bits_rdata = io_dmem_resp_bits_rdata;
  assign executeStage_io_mmio_req_ready = io_mmio_req_ready;
  assign executeStage_io_mmio_resp_valid = io_mmio_resp_valid;
  assign executeStage_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata;
  assign executeStage_io_out_ready = 1'h1;
  assign writeBackUnit_clock = clock;
  assign writeBackUnit_reset = reset;
  assign writeBackUnit_io_in_valid = executeStage_io_out_valid;
  assign writeBackUnit_io_in_bits_valid = executeStage_io_out_bits_valid;
  assign writeBackUnit_io_in_bits_wen = executeStage_io_out_bits_wen;
  assign writeBackUnit_io_in_bits_wb_addr = executeStage_io_out_bits_wb_addr;
  assign writeBackUnit_io_in_bits_wb_data = executeStage_io_out_bits_wb_data;
  assign writeBackUnit_io_in_bits_redirect_valid = executeStage_io_out_bits_redirect_valid;
  assign writeBackUnit_io_in_bits_redirect_target = executeStage_io_out_bits_redirect_target;
  assign writeBackUnit_io_in_bits_flush = writeBackUnit_io_redirect_valid;
  assign regFile_clock = clock;
  assign regFile_reset = reset;
  assign regFile_io_r_rs1_addr = decodeStage_io_regFile_rs1_addr;
  assign regFile_io_r_rs2_addr = decodeStage_io_regFile_rs2_addr;
  assign regFile_io_w_w_addr = writeBackUnit_io_regFile_w_addr;
  assign regFile_io_w_w_data = writeBackUnit_io_regFile_w_data;
  assign regFile_io_w_wen = writeBackUnit_io_regFile_wen;
  always @(posedge clock) begin
    if (reset) begin
      pipelineRegs_pc <= 32'h0;
    end else if (_T_9) begin
      pipelineRegs_pc <= 32'h0;
    end else if (_T_4) begin
      pipelineRegs_pc <= decodeStage_io_out_bits_pc;
    end
    if (reset) begin
      pipelineRegs_inst <= 32'h0;
    end else if (_T_9) begin
      pipelineRegs_inst <= 32'h0;
    end else if (_T_4) begin
      pipelineRegs_inst <= decodeStage_io_out_bits_inst;
    end
    if (reset) begin
      pipelineRegs_valid <= 1'h0;
    end else if (_T_9) begin
      pipelineRegs_valid <= 1'h0;
    end else if (_T_4) begin
      pipelineRegs_valid <= decodeStage_io_out_bits_valid;
    end
    if (reset) begin
      pipelineRegs_bubble <= 1'h0;
    end else if (_T_9) begin
      pipelineRegs_bubble <= 1'h0;
    end else if (_T_4) begin
      pipelineRegs_bubble <= decodeStage_io_out_bits_bubble;
    end
    if (reset) begin
      pipelineRegs_opcode_type <= 3'h0;
    end else if (_T_9) begin
      pipelineRegs_opcode_type <= 3'h0;
    end else if (_T_4) begin
      pipelineRegs_opcode_type <= decodeStage_io_out_bits_opcode_type;
    end
    if (reset) begin
      pipelineRegs_opcode_func <= 6'h0;
    end else if (_T_9) begin
      pipelineRegs_opcode_func <= 6'h0;
    end else if (_T_4) begin
      pipelineRegs_opcode_func <= decodeStage_io_out_bits_opcode_func;
    end
    if (reset) begin
      pipelineRegs_br_type <= 4'h0;
    end else if (_T_9) begin
      pipelineRegs_br_type <= 4'h0;
    end else if (_T_4) begin
      pipelineRegs_br_type <= decodeStage_io_out_bits_br_type;
    end
    if (reset) begin
      pipelineRegs_rf_en <= 1'h0;
    end else if (_T_9) begin
      pipelineRegs_rf_en <= 1'h0;
    end else if (_T_4) begin
      pipelineRegs_rf_en <= decodeStage_io_out_bits_rf_en;
    end
    if (reset) begin
      pipelineRegs_wb_addr <= 5'h0;
    end else if (_T_9) begin
      pipelineRegs_wb_addr <= 5'h0;
    end else if (_T_4) begin
      pipelineRegs_wb_addr <= decodeStage_io_out_bits_wb_addr;
    end
    if (reset) begin
      pipelineRegs_wb_stage <= 2'h0;
    end else if (_T_9) begin
      pipelineRegs_wb_stage <= 2'h0;
    end else if (_T_4) begin
      pipelineRegs_wb_stage <= decodeStage_io_out_bits_wb_stage;
    end
    if (reset) begin
      pipelineRegs_op1_data <= 64'h0;
    end else if (_T_9) begin
      pipelineRegs_op1_data <= 64'h0;
    end else if (_T_4) begin
      pipelineRegs_op1_data <= decodeStage_io_out_bits_op1_data;
    end
    if (reset) begin
      pipelineRegs_op2_data <= 64'h0;
    end else if (_T_9) begin
      pipelineRegs_op2_data <= 64'h0;
    end else if (_T_4) begin
      pipelineRegs_op2_data <= decodeStage_io_out_bits_op2_data;
    end
    if (reset) begin
      pipelineRegs_rs1_data <= 64'h0;
    end else if (_T_9) begin
      pipelineRegs_rs1_data <= 64'h0;
    end else if (_T_4) begin
      pipelineRegs_rs1_data <= decodeStage_io_out_bits_rs1_data;
    end
    if (reset) begin
      pipelineRegs_rs2_data <= 64'h0;
    end else if (_T_9) begin
      pipelineRegs_rs2_data <= 64'h0;
    end else if (_T_4) begin
      pipelineRegs_rs2_data <= decodeStage_io_out_bits_rs2_data;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pipelineRegs_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  pipelineRegs_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  pipelineRegs_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipelineRegs_bubble = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipelineRegs_opcode_type = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  pipelineRegs_opcode_func = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  pipelineRegs_br_type = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  pipelineRegs_rf_en = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pipelineRegs_wb_addr = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  pipelineRegs_wb_stage = _RAND_9[1:0];
  _RAND_10 = {2{`RANDOM}};
  pipelineRegs_op1_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  pipelineRegs_op2_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pipelineRegs_rs1_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pipelineRegs_rs2_data = _RAND_13[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_MyCore(
  input         clock,
  input         reset,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [1:0]  io_dmem_req_bits_size,
  output [2:0]  io_dmem_req_bits_cmd,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_imem_req_ready,
  output [31:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_dmmio_req_ready,
  output        io_dmmio_req_valid,
  output [31:0] io_dmmio_req_bits_addr,
  output [63:0] io_dmmio_req_bits_wdata,
  output [1:0]  io_dmmio_req_bits_size,
  output [2:0]  io_dmmio_req_bits_cmd,
  input         io_dmmio_resp_valid,
  input  [63:0] io_dmmio_resp_bits_rdata,
  output        flushICache
);
  wire  fetch_clock;
  wire  fetch_reset;
  wire  fetch_io_imem_req_ready;
  wire  fetch_io_imem_req_valid;
  wire [31:0] fetch_io_imem_req_bits_addr;
  wire  fetch_io_imem_resp_ready;
  wire  fetch_io_imem_resp_valid;
  wire [63:0] fetch_io_imem_resp_bits_rdata;
  wire  fetch_io_out_ready;
  wire  fetch_io_out_valid;
  wire [31:0] fetch_io_out_bits_inst;
  wire [31:0] fetch_io_out_bits_pc;
  wire  fetch_io_redirect_valid;
  wire [31:0] fetch_io_redirect_target;
  wire  pipeline_clock;
  wire  pipeline_reset;
  wire  pipeline_io_in_ready;
  wire  pipeline_io_in_valid;
  wire [31:0] pipeline_io_in_bits_inst;
  wire [31:0] pipeline_io_in_bits_pc;
  wire  pipeline_io_dmem_req_ready;
  wire  pipeline_io_dmem_req_valid;
  wire [31:0] pipeline_io_dmem_req_bits_addr;
  wire [63:0] pipeline_io_dmem_req_bits_wdata;
  wire [1:0] pipeline_io_dmem_req_bits_size;
  wire [2:0] pipeline_io_dmem_req_bits_cmd;
  wire  pipeline_io_dmem_resp_valid;
  wire [63:0] pipeline_io_dmem_resp_bits_rdata;
  wire  pipeline_io_mmio_req_ready;
  wire  pipeline_io_mmio_req_valid;
  wire [31:0] pipeline_io_mmio_req_bits_addr;
  wire [63:0] pipeline_io_mmio_req_bits_wdata;
  wire [1:0] pipeline_io_mmio_req_bits_size;
  wire [2:0] pipeline_io_mmio_req_bits_cmd;
  wire  pipeline_io_mmio_resp_valid;
  wire [63:0] pipeline_io_mmio_resp_bits_rdata;
  wire  pipeline_io_redirect_valid;
  wire [31:0] pipeline_io_redirect_target;
  wire  pipeline_flushICache;
  ysyx_040656_InstructionFetchUnit fetch (
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_imem_req_ready(fetch_io_imem_req_ready),
    .io_imem_req_valid(fetch_io_imem_req_valid),
    .io_imem_req_bits_addr(fetch_io_imem_req_bits_addr),
    .io_imem_resp_ready(fetch_io_imem_resp_ready),
    .io_imem_resp_valid(fetch_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(fetch_io_imem_resp_bits_rdata),
    .io_out_ready(fetch_io_out_ready),
    .io_out_valid(fetch_io_out_valid),
    .io_out_bits_inst(fetch_io_out_bits_inst),
    .io_out_bits_pc(fetch_io_out_bits_pc),
    .io_redirect_valid(fetch_io_redirect_valid),
    .io_redirect_target(fetch_io_redirect_target)
  );
  ysyx_040656_Pipeline pipeline (
    .clock(pipeline_clock),
    .reset(pipeline_reset),
    .io_in_ready(pipeline_io_in_ready),
    .io_in_valid(pipeline_io_in_valid),
    .io_in_bits_inst(pipeline_io_in_bits_inst),
    .io_in_bits_pc(pipeline_io_in_bits_pc),
    .io_dmem_req_ready(pipeline_io_dmem_req_ready),
    .io_dmem_req_valid(pipeline_io_dmem_req_valid),
    .io_dmem_req_bits_addr(pipeline_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(pipeline_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_size(pipeline_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(pipeline_io_dmem_req_bits_cmd),
    .io_dmem_resp_valid(pipeline_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(pipeline_io_dmem_resp_bits_rdata),
    .io_mmio_req_ready(pipeline_io_mmio_req_ready),
    .io_mmio_req_valid(pipeline_io_mmio_req_valid),
    .io_mmio_req_bits_addr(pipeline_io_mmio_req_bits_addr),
    .io_mmio_req_bits_wdata(pipeline_io_mmio_req_bits_wdata),
    .io_mmio_req_bits_size(pipeline_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(pipeline_io_mmio_req_bits_cmd),
    .io_mmio_resp_valid(pipeline_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(pipeline_io_mmio_resp_bits_rdata),
    .io_redirect_valid(pipeline_io_redirect_valid),
    .io_redirect_target(pipeline_io_redirect_target),
    .flushICache(pipeline_flushICache)
  );
  assign io_dmem_req_valid = pipeline_io_dmem_req_valid;
  assign io_dmem_req_bits_addr = pipeline_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_wdata = pipeline_io_dmem_req_bits_wdata;
  assign io_dmem_req_bits_size = pipeline_io_dmem_req_bits_size;
  assign io_dmem_req_bits_cmd = pipeline_io_dmem_req_bits_cmd;
  assign io_imem_req_bits_addr = fetch_io_imem_req_bits_addr;
  assign io_imem_resp_ready = fetch_io_imem_resp_ready;
  assign io_dmmio_req_valid = pipeline_io_mmio_req_valid;
  assign io_dmmio_req_bits_addr = pipeline_io_mmio_req_bits_addr;
  assign io_dmmio_req_bits_wdata = pipeline_io_mmio_req_bits_wdata;
  assign io_dmmio_req_bits_size = pipeline_io_mmio_req_bits_size;
  assign io_dmmio_req_bits_cmd = pipeline_io_mmio_req_bits_cmd;
  assign flushICache = pipeline_flushICache;
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_imem_req_ready = io_imem_req_ready;
  assign fetch_io_imem_resp_valid = io_imem_resp_valid;
  assign fetch_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata;
  assign fetch_io_out_ready = pipeline_io_in_ready;
  assign fetch_io_redirect_valid = pipeline_io_redirect_valid;
  assign fetch_io_redirect_target = pipeline_io_redirect_target;
  assign pipeline_clock = clock;
  assign pipeline_reset = reset;
  assign pipeline_io_in_valid = fetch_io_out_valid;
  assign pipeline_io_in_bits_inst = fetch_io_out_bits_inst;
  assign pipeline_io_in_bits_pc = fetch_io_out_bits_pc;
  assign pipeline_io_dmem_req_ready = io_dmem_req_ready;
  assign pipeline_io_dmem_resp_valid = io_dmem_resp_valid;
  assign pipeline_io_dmem_resp_bits_rdata = io_dmem_resp_bits_rdata;
  assign pipeline_io_mmio_req_ready = io_dmmio_req_ready;
  assign pipeline_io_mmio_resp_valid = io_dmmio_resp_valid;
  assign pipeline_io_mmio_resp_bits_rdata = io_dmmio_resp_bits_rdata;
endmodule
module ysyx_040656_SRAM(
  input         clock,
  input         reset,
  input  [5:0]  io_w_setIdx,
  input  [21:0] io_w_data_tag,
  input         io_w_data_valid,
  input         io_w_data_needFlush,
  input         io_w_wen,
  input  [5:0]  io_r_setIdx,
  output [21:0] io_r_data_tag,
  output        io_r_data_valid,
  output        io_r_data_needFlush,
  input         io_r_ren
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif
  reg [23:0] ram [0:63];
  wire  ram_rdata_MPORT_en;
  wire [5:0] ram_rdata_MPORT_addr;
  wire [23:0] ram_rdata_MPORT_data;
  wire [23:0] ram_MPORT_data;
  wire [5:0] ram_MPORT_addr;
  wire  ram_MPORT_mask;
  wire  ram_MPORT_en;
  wire [23:0] ram_MPORT_1_data;
  wire [5:0] ram_MPORT_1_addr;
  wire  ram_MPORT_1_mask;
  wire  ram_MPORT_1_en;
  wire [23:0] ram_MPORT_2_data;
  wire [5:0] ram_MPORT_2_addr;
  wire  ram_MPORT_2_mask;
  wire  ram_MPORT_2_en;
  wire [23:0] ram_MPORT_3_data;
  wire [5:0] ram_MPORT_3_addr;
  wire  ram_MPORT_3_mask;
  wire  ram_MPORT_3_en;
  wire [23:0] ram_MPORT_4_data;
  wire [5:0] ram_MPORT_4_addr;
  wire  ram_MPORT_4_mask;
  wire  ram_MPORT_4_en;
  wire [23:0] ram_MPORT_5_data;
  wire [5:0] ram_MPORT_5_addr;
  wire  ram_MPORT_5_mask;
  wire  ram_MPORT_5_en;
  wire [23:0] ram_MPORT_6_data;
  wire [5:0] ram_MPORT_6_addr;
  wire  ram_MPORT_6_mask;
  wire  ram_MPORT_6_en;
  wire [23:0] ram_MPORT_7_data;
  wire [5:0] ram_MPORT_7_addr;
  wire  ram_MPORT_7_mask;
  wire  ram_MPORT_7_en;
  wire [23:0] ram_MPORT_8_data;
  wire [5:0] ram_MPORT_8_addr;
  wire  ram_MPORT_8_mask;
  wire  ram_MPORT_8_en;
  wire [23:0] ram_MPORT_9_data;
  wire [5:0] ram_MPORT_9_addr;
  wire  ram_MPORT_9_mask;
  wire  ram_MPORT_9_en;
  wire [23:0] ram_MPORT_10_data;
  wire [5:0] ram_MPORT_10_addr;
  wire  ram_MPORT_10_mask;
  wire  ram_MPORT_10_en;
  wire [23:0] ram_MPORT_11_data;
  wire [5:0] ram_MPORT_11_addr;
  wire  ram_MPORT_11_mask;
  wire  ram_MPORT_11_en;
  wire [23:0] ram_MPORT_12_data;
  wire [5:0] ram_MPORT_12_addr;
  wire  ram_MPORT_12_mask;
  wire  ram_MPORT_12_en;
  wire [23:0] ram_MPORT_13_data;
  wire [5:0] ram_MPORT_13_addr;
  wire  ram_MPORT_13_mask;
  wire  ram_MPORT_13_en;
  wire [23:0] ram_MPORT_14_data;
  wire [5:0] ram_MPORT_14_addr;
  wire  ram_MPORT_14_mask;
  wire  ram_MPORT_14_en;
  wire [23:0] ram_MPORT_15_data;
  wire [5:0] ram_MPORT_15_addr;
  wire  ram_MPORT_15_mask;
  wire  ram_MPORT_15_en;
  wire [23:0] ram_MPORT_16_data;
  wire [5:0] ram_MPORT_16_addr;
  wire  ram_MPORT_16_mask;
  wire  ram_MPORT_16_en;
  wire [23:0] ram_MPORT_17_data;
  wire [5:0] ram_MPORT_17_addr;
  wire  ram_MPORT_17_mask;
  wire  ram_MPORT_17_en;
  wire [23:0] ram_MPORT_18_data;
  wire [5:0] ram_MPORT_18_addr;
  wire  ram_MPORT_18_mask;
  wire  ram_MPORT_18_en;
  wire [23:0] ram_MPORT_19_data;
  wire [5:0] ram_MPORT_19_addr;
  wire  ram_MPORT_19_mask;
  wire  ram_MPORT_19_en;
  wire [23:0] ram_MPORT_20_data;
  wire [5:0] ram_MPORT_20_addr;
  wire  ram_MPORT_20_mask;
  wire  ram_MPORT_20_en;
  wire [23:0] ram_MPORT_21_data;
  wire [5:0] ram_MPORT_21_addr;
  wire  ram_MPORT_21_mask;
  wire  ram_MPORT_21_en;
  wire [23:0] ram_MPORT_22_data;
  wire [5:0] ram_MPORT_22_addr;
  wire  ram_MPORT_22_mask;
  wire  ram_MPORT_22_en;
  wire [23:0] ram_MPORT_23_data;
  wire [5:0] ram_MPORT_23_addr;
  wire  ram_MPORT_23_mask;
  wire  ram_MPORT_23_en;
  wire [23:0] ram_MPORT_24_data;
  wire [5:0] ram_MPORT_24_addr;
  wire  ram_MPORT_24_mask;
  wire  ram_MPORT_24_en;
  wire [23:0] ram_MPORT_25_data;
  wire [5:0] ram_MPORT_25_addr;
  wire  ram_MPORT_25_mask;
  wire  ram_MPORT_25_en;
  wire [23:0] ram_MPORT_26_data;
  wire [5:0] ram_MPORT_26_addr;
  wire  ram_MPORT_26_mask;
  wire  ram_MPORT_26_en;
  wire [23:0] ram_MPORT_27_data;
  wire [5:0] ram_MPORT_27_addr;
  wire  ram_MPORT_27_mask;
  wire  ram_MPORT_27_en;
  wire [23:0] ram_MPORT_28_data;
  wire [5:0] ram_MPORT_28_addr;
  wire  ram_MPORT_28_mask;
  wire  ram_MPORT_28_en;
  wire [23:0] ram_MPORT_29_data;
  wire [5:0] ram_MPORT_29_addr;
  wire  ram_MPORT_29_mask;
  wire  ram_MPORT_29_en;
  wire [23:0] ram_MPORT_30_data;
  wire [5:0] ram_MPORT_30_addr;
  wire  ram_MPORT_30_mask;
  wire  ram_MPORT_30_en;
  wire [23:0] ram_MPORT_31_data;
  wire [5:0] ram_MPORT_31_addr;
  wire  ram_MPORT_31_mask;
  wire  ram_MPORT_31_en;
  wire [23:0] ram_MPORT_32_data;
  wire [5:0] ram_MPORT_32_addr;
  wire  ram_MPORT_32_mask;
  wire  ram_MPORT_32_en;
  wire [23:0] ram_MPORT_33_data;
  wire [5:0] ram_MPORT_33_addr;
  wire  ram_MPORT_33_mask;
  wire  ram_MPORT_33_en;
  wire [23:0] ram_MPORT_34_data;
  wire [5:0] ram_MPORT_34_addr;
  wire  ram_MPORT_34_mask;
  wire  ram_MPORT_34_en;
  wire [23:0] ram_MPORT_35_data;
  wire [5:0] ram_MPORT_35_addr;
  wire  ram_MPORT_35_mask;
  wire  ram_MPORT_35_en;
  wire [23:0] ram_MPORT_36_data;
  wire [5:0] ram_MPORT_36_addr;
  wire  ram_MPORT_36_mask;
  wire  ram_MPORT_36_en;
  wire [23:0] ram_MPORT_37_data;
  wire [5:0] ram_MPORT_37_addr;
  wire  ram_MPORT_37_mask;
  wire  ram_MPORT_37_en;
  wire [23:0] ram_MPORT_38_data;
  wire [5:0] ram_MPORT_38_addr;
  wire  ram_MPORT_38_mask;
  wire  ram_MPORT_38_en;
  wire [23:0] ram_MPORT_39_data;
  wire [5:0] ram_MPORT_39_addr;
  wire  ram_MPORT_39_mask;
  wire  ram_MPORT_39_en;
  wire [23:0] ram_MPORT_40_data;
  wire [5:0] ram_MPORT_40_addr;
  wire  ram_MPORT_40_mask;
  wire  ram_MPORT_40_en;
  wire [23:0] ram_MPORT_41_data;
  wire [5:0] ram_MPORT_41_addr;
  wire  ram_MPORT_41_mask;
  wire  ram_MPORT_41_en;
  wire [23:0] ram_MPORT_42_data;
  wire [5:0] ram_MPORT_42_addr;
  wire  ram_MPORT_42_mask;
  wire  ram_MPORT_42_en;
  wire [23:0] ram_MPORT_43_data;
  wire [5:0] ram_MPORT_43_addr;
  wire  ram_MPORT_43_mask;
  wire  ram_MPORT_43_en;
  wire [23:0] ram_MPORT_44_data;
  wire [5:0] ram_MPORT_44_addr;
  wire  ram_MPORT_44_mask;
  wire  ram_MPORT_44_en;
  wire [23:0] ram_MPORT_45_data;
  wire [5:0] ram_MPORT_45_addr;
  wire  ram_MPORT_45_mask;
  wire  ram_MPORT_45_en;
  wire [23:0] ram_MPORT_46_data;
  wire [5:0] ram_MPORT_46_addr;
  wire  ram_MPORT_46_mask;
  wire  ram_MPORT_46_en;
  wire [23:0] ram_MPORT_47_data;
  wire [5:0] ram_MPORT_47_addr;
  wire  ram_MPORT_47_mask;
  wire  ram_MPORT_47_en;
  wire [23:0] ram_MPORT_48_data;
  wire [5:0] ram_MPORT_48_addr;
  wire  ram_MPORT_48_mask;
  wire  ram_MPORT_48_en;
  wire [23:0] ram_MPORT_49_data;
  wire [5:0] ram_MPORT_49_addr;
  wire  ram_MPORT_49_mask;
  wire  ram_MPORT_49_en;
  wire [23:0] ram_MPORT_50_data;
  wire [5:0] ram_MPORT_50_addr;
  wire  ram_MPORT_50_mask;
  wire  ram_MPORT_50_en;
  wire [23:0] ram_MPORT_51_data;
  wire [5:0] ram_MPORT_51_addr;
  wire  ram_MPORT_51_mask;
  wire  ram_MPORT_51_en;
  wire [23:0] ram_MPORT_52_data;
  wire [5:0] ram_MPORT_52_addr;
  wire  ram_MPORT_52_mask;
  wire  ram_MPORT_52_en;
  wire [23:0] ram_MPORT_53_data;
  wire [5:0] ram_MPORT_53_addr;
  wire  ram_MPORT_53_mask;
  wire  ram_MPORT_53_en;
  wire [23:0] ram_MPORT_54_data;
  wire [5:0] ram_MPORT_54_addr;
  wire  ram_MPORT_54_mask;
  wire  ram_MPORT_54_en;
  wire [23:0] ram_MPORT_55_data;
  wire [5:0] ram_MPORT_55_addr;
  wire  ram_MPORT_55_mask;
  wire  ram_MPORT_55_en;
  wire [23:0] ram_MPORT_56_data;
  wire [5:0] ram_MPORT_56_addr;
  wire  ram_MPORT_56_mask;
  wire  ram_MPORT_56_en;
  wire [23:0] ram_MPORT_57_data;
  wire [5:0] ram_MPORT_57_addr;
  wire  ram_MPORT_57_mask;
  wire  ram_MPORT_57_en;
  wire [23:0] ram_MPORT_58_data;
  wire [5:0] ram_MPORT_58_addr;
  wire  ram_MPORT_58_mask;
  wire  ram_MPORT_58_en;
  wire [23:0] ram_MPORT_59_data;
  wire [5:0] ram_MPORT_59_addr;
  wire  ram_MPORT_59_mask;
  wire  ram_MPORT_59_en;
  wire [23:0] ram_MPORT_60_data;
  wire [5:0] ram_MPORT_60_addr;
  wire  ram_MPORT_60_mask;
  wire  ram_MPORT_60_en;
  wire [23:0] ram_MPORT_61_data;
  wire [5:0] ram_MPORT_61_addr;
  wire  ram_MPORT_61_mask;
  wire  ram_MPORT_61_en;
  wire [23:0] ram_MPORT_62_data;
  wire [5:0] ram_MPORT_62_addr;
  wire  ram_MPORT_62_mask;
  wire  ram_MPORT_62_en;
  wire [23:0] ram_MPORT_63_data;
  wire [5:0] ram_MPORT_63_addr;
  wire  ram_MPORT_63_mask;
  wire  ram_MPORT_63_en;
  wire [23:0] ram_MPORT_64_data;
  wire [5:0] ram_MPORT_64_addr;
  wire  ram_MPORT_64_mask;
  wire  ram_MPORT_64_en;
  reg  ram_rdata_MPORT_en_pipe_0;
  reg [5:0] ram_rdata_MPORT_addr_pipe_0;
  wire  _realRen_T = ~io_w_wen;
  wire [22:0] wdata_hi = {io_w_data_tag,io_w_data_valid};
  reg  rdata_REG;
  reg [23:0] rdata_r;
  wire [23:0] _GEN_9 = rdata_REG ? ram_rdata_MPORT_data : rdata_r;
  assign ram_rdata_MPORT_en = ram_rdata_MPORT_en_pipe_0;
  assign ram_rdata_MPORT_addr = ram_rdata_MPORT_addr_pipe_0;
  assign ram_rdata_MPORT_data = ram[ram_rdata_MPORT_addr];
  assign ram_MPORT_data = {wdata_hi,io_w_data_needFlush};
  assign ram_MPORT_addr = io_w_setIdx;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_w_wen;
  assign ram_MPORT_1_data = 24'h0;
  assign ram_MPORT_1_addr = 6'h0;
  assign ram_MPORT_1_mask = 1'h1;
  assign ram_MPORT_1_en = reset;
  assign ram_MPORT_2_data = 24'h0;
  assign ram_MPORT_2_addr = 6'h1;
  assign ram_MPORT_2_mask = 1'h1;
  assign ram_MPORT_2_en = reset;
  assign ram_MPORT_3_data = 24'h0;
  assign ram_MPORT_3_addr = 6'h2;
  assign ram_MPORT_3_mask = 1'h1;
  assign ram_MPORT_3_en = reset;
  assign ram_MPORT_4_data = 24'h0;
  assign ram_MPORT_4_addr = 6'h3;
  assign ram_MPORT_4_mask = 1'h1;
  assign ram_MPORT_4_en = reset;
  assign ram_MPORT_5_data = 24'h0;
  assign ram_MPORT_5_addr = 6'h4;
  assign ram_MPORT_5_mask = 1'h1;
  assign ram_MPORT_5_en = reset;
  assign ram_MPORT_6_data = 24'h0;
  assign ram_MPORT_6_addr = 6'h5;
  assign ram_MPORT_6_mask = 1'h1;
  assign ram_MPORT_6_en = reset;
  assign ram_MPORT_7_data = 24'h0;
  assign ram_MPORT_7_addr = 6'h6;
  assign ram_MPORT_7_mask = 1'h1;
  assign ram_MPORT_7_en = reset;
  assign ram_MPORT_8_data = 24'h0;
  assign ram_MPORT_8_addr = 6'h7;
  assign ram_MPORT_8_mask = 1'h1;
  assign ram_MPORT_8_en = reset;
  assign ram_MPORT_9_data = 24'h0;
  assign ram_MPORT_9_addr = 6'h8;
  assign ram_MPORT_9_mask = 1'h1;
  assign ram_MPORT_9_en = reset;
  assign ram_MPORT_10_data = 24'h0;
  assign ram_MPORT_10_addr = 6'h9;
  assign ram_MPORT_10_mask = 1'h1;
  assign ram_MPORT_10_en = reset;
  assign ram_MPORT_11_data = 24'h0;
  assign ram_MPORT_11_addr = 6'ha;
  assign ram_MPORT_11_mask = 1'h1;
  assign ram_MPORT_11_en = reset;
  assign ram_MPORT_12_data = 24'h0;
  assign ram_MPORT_12_addr = 6'hb;
  assign ram_MPORT_12_mask = 1'h1;
  assign ram_MPORT_12_en = reset;
  assign ram_MPORT_13_data = 24'h0;
  assign ram_MPORT_13_addr = 6'hc;
  assign ram_MPORT_13_mask = 1'h1;
  assign ram_MPORT_13_en = reset;
  assign ram_MPORT_14_data = 24'h0;
  assign ram_MPORT_14_addr = 6'hd;
  assign ram_MPORT_14_mask = 1'h1;
  assign ram_MPORT_14_en = reset;
  assign ram_MPORT_15_data = 24'h0;
  assign ram_MPORT_15_addr = 6'he;
  assign ram_MPORT_15_mask = 1'h1;
  assign ram_MPORT_15_en = reset;
  assign ram_MPORT_16_data = 24'h0;
  assign ram_MPORT_16_addr = 6'hf;
  assign ram_MPORT_16_mask = 1'h1;
  assign ram_MPORT_16_en = reset;
  assign ram_MPORT_17_data = 24'h0;
  assign ram_MPORT_17_addr = 6'h10;
  assign ram_MPORT_17_mask = 1'h1;
  assign ram_MPORT_17_en = reset;
  assign ram_MPORT_18_data = 24'h0;
  assign ram_MPORT_18_addr = 6'h11;
  assign ram_MPORT_18_mask = 1'h1;
  assign ram_MPORT_18_en = reset;
  assign ram_MPORT_19_data = 24'h0;
  assign ram_MPORT_19_addr = 6'h12;
  assign ram_MPORT_19_mask = 1'h1;
  assign ram_MPORT_19_en = reset;
  assign ram_MPORT_20_data = 24'h0;
  assign ram_MPORT_20_addr = 6'h13;
  assign ram_MPORT_20_mask = 1'h1;
  assign ram_MPORT_20_en = reset;
  assign ram_MPORT_21_data = 24'h0;
  assign ram_MPORT_21_addr = 6'h14;
  assign ram_MPORT_21_mask = 1'h1;
  assign ram_MPORT_21_en = reset;
  assign ram_MPORT_22_data = 24'h0;
  assign ram_MPORT_22_addr = 6'h15;
  assign ram_MPORT_22_mask = 1'h1;
  assign ram_MPORT_22_en = reset;
  assign ram_MPORT_23_data = 24'h0;
  assign ram_MPORT_23_addr = 6'h16;
  assign ram_MPORT_23_mask = 1'h1;
  assign ram_MPORT_23_en = reset;
  assign ram_MPORT_24_data = 24'h0;
  assign ram_MPORT_24_addr = 6'h17;
  assign ram_MPORT_24_mask = 1'h1;
  assign ram_MPORT_24_en = reset;
  assign ram_MPORT_25_data = 24'h0;
  assign ram_MPORT_25_addr = 6'h18;
  assign ram_MPORT_25_mask = 1'h1;
  assign ram_MPORT_25_en = reset;
  assign ram_MPORT_26_data = 24'h0;
  assign ram_MPORT_26_addr = 6'h19;
  assign ram_MPORT_26_mask = 1'h1;
  assign ram_MPORT_26_en = reset;
  assign ram_MPORT_27_data = 24'h0;
  assign ram_MPORT_27_addr = 6'h1a;
  assign ram_MPORT_27_mask = 1'h1;
  assign ram_MPORT_27_en = reset;
  assign ram_MPORT_28_data = 24'h0;
  assign ram_MPORT_28_addr = 6'h1b;
  assign ram_MPORT_28_mask = 1'h1;
  assign ram_MPORT_28_en = reset;
  assign ram_MPORT_29_data = 24'h0;
  assign ram_MPORT_29_addr = 6'h1c;
  assign ram_MPORT_29_mask = 1'h1;
  assign ram_MPORT_29_en = reset;
  assign ram_MPORT_30_data = 24'h0;
  assign ram_MPORT_30_addr = 6'h1d;
  assign ram_MPORT_30_mask = 1'h1;
  assign ram_MPORT_30_en = reset;
  assign ram_MPORT_31_data = 24'h0;
  assign ram_MPORT_31_addr = 6'h1e;
  assign ram_MPORT_31_mask = 1'h1;
  assign ram_MPORT_31_en = reset;
  assign ram_MPORT_32_data = 24'h0;
  assign ram_MPORT_32_addr = 6'h1f;
  assign ram_MPORT_32_mask = 1'h1;
  assign ram_MPORT_32_en = reset;
  assign ram_MPORT_33_data = 24'h0;
  assign ram_MPORT_33_addr = 6'h20;
  assign ram_MPORT_33_mask = 1'h1;
  assign ram_MPORT_33_en = reset;
  assign ram_MPORT_34_data = 24'h0;
  assign ram_MPORT_34_addr = 6'h21;
  assign ram_MPORT_34_mask = 1'h1;
  assign ram_MPORT_34_en = reset;
  assign ram_MPORT_35_data = 24'h0;
  assign ram_MPORT_35_addr = 6'h22;
  assign ram_MPORT_35_mask = 1'h1;
  assign ram_MPORT_35_en = reset;
  assign ram_MPORT_36_data = 24'h0;
  assign ram_MPORT_36_addr = 6'h23;
  assign ram_MPORT_36_mask = 1'h1;
  assign ram_MPORT_36_en = reset;
  assign ram_MPORT_37_data = 24'h0;
  assign ram_MPORT_37_addr = 6'h24;
  assign ram_MPORT_37_mask = 1'h1;
  assign ram_MPORT_37_en = reset;
  assign ram_MPORT_38_data = 24'h0;
  assign ram_MPORT_38_addr = 6'h25;
  assign ram_MPORT_38_mask = 1'h1;
  assign ram_MPORT_38_en = reset;
  assign ram_MPORT_39_data = 24'h0;
  assign ram_MPORT_39_addr = 6'h26;
  assign ram_MPORT_39_mask = 1'h1;
  assign ram_MPORT_39_en = reset;
  assign ram_MPORT_40_data = 24'h0;
  assign ram_MPORT_40_addr = 6'h27;
  assign ram_MPORT_40_mask = 1'h1;
  assign ram_MPORT_40_en = reset;
  assign ram_MPORT_41_data = 24'h0;
  assign ram_MPORT_41_addr = 6'h28;
  assign ram_MPORT_41_mask = 1'h1;
  assign ram_MPORT_41_en = reset;
  assign ram_MPORT_42_data = 24'h0;
  assign ram_MPORT_42_addr = 6'h29;
  assign ram_MPORT_42_mask = 1'h1;
  assign ram_MPORT_42_en = reset;
  assign ram_MPORT_43_data = 24'h0;
  assign ram_MPORT_43_addr = 6'h2a;
  assign ram_MPORT_43_mask = 1'h1;
  assign ram_MPORT_43_en = reset;
  assign ram_MPORT_44_data = 24'h0;
  assign ram_MPORT_44_addr = 6'h2b;
  assign ram_MPORT_44_mask = 1'h1;
  assign ram_MPORT_44_en = reset;
  assign ram_MPORT_45_data = 24'h0;
  assign ram_MPORT_45_addr = 6'h2c;
  assign ram_MPORT_45_mask = 1'h1;
  assign ram_MPORT_45_en = reset;
  assign ram_MPORT_46_data = 24'h0;
  assign ram_MPORT_46_addr = 6'h2d;
  assign ram_MPORT_46_mask = 1'h1;
  assign ram_MPORT_46_en = reset;
  assign ram_MPORT_47_data = 24'h0;
  assign ram_MPORT_47_addr = 6'h2e;
  assign ram_MPORT_47_mask = 1'h1;
  assign ram_MPORT_47_en = reset;
  assign ram_MPORT_48_data = 24'h0;
  assign ram_MPORT_48_addr = 6'h2f;
  assign ram_MPORT_48_mask = 1'h1;
  assign ram_MPORT_48_en = reset;
  assign ram_MPORT_49_data = 24'h0;
  assign ram_MPORT_49_addr = 6'h30;
  assign ram_MPORT_49_mask = 1'h1;
  assign ram_MPORT_49_en = reset;
  assign ram_MPORT_50_data = 24'h0;
  assign ram_MPORT_50_addr = 6'h31;
  assign ram_MPORT_50_mask = 1'h1;
  assign ram_MPORT_50_en = reset;
  assign ram_MPORT_51_data = 24'h0;
  assign ram_MPORT_51_addr = 6'h32;
  assign ram_MPORT_51_mask = 1'h1;
  assign ram_MPORT_51_en = reset;
  assign ram_MPORT_52_data = 24'h0;
  assign ram_MPORT_52_addr = 6'h33;
  assign ram_MPORT_52_mask = 1'h1;
  assign ram_MPORT_52_en = reset;
  assign ram_MPORT_53_data = 24'h0;
  assign ram_MPORT_53_addr = 6'h34;
  assign ram_MPORT_53_mask = 1'h1;
  assign ram_MPORT_53_en = reset;
  assign ram_MPORT_54_data = 24'h0;
  assign ram_MPORT_54_addr = 6'h35;
  assign ram_MPORT_54_mask = 1'h1;
  assign ram_MPORT_54_en = reset;
  assign ram_MPORT_55_data = 24'h0;
  assign ram_MPORT_55_addr = 6'h36;
  assign ram_MPORT_55_mask = 1'h1;
  assign ram_MPORT_55_en = reset;
  assign ram_MPORT_56_data = 24'h0;
  assign ram_MPORT_56_addr = 6'h37;
  assign ram_MPORT_56_mask = 1'h1;
  assign ram_MPORT_56_en = reset;
  assign ram_MPORT_57_data = 24'h0;
  assign ram_MPORT_57_addr = 6'h38;
  assign ram_MPORT_57_mask = 1'h1;
  assign ram_MPORT_57_en = reset;
  assign ram_MPORT_58_data = 24'h0;
  assign ram_MPORT_58_addr = 6'h39;
  assign ram_MPORT_58_mask = 1'h1;
  assign ram_MPORT_58_en = reset;
  assign ram_MPORT_59_data = 24'h0;
  assign ram_MPORT_59_addr = 6'h3a;
  assign ram_MPORT_59_mask = 1'h1;
  assign ram_MPORT_59_en = reset;
  assign ram_MPORT_60_data = 24'h0;
  assign ram_MPORT_60_addr = 6'h3b;
  assign ram_MPORT_60_mask = 1'h1;
  assign ram_MPORT_60_en = reset;
  assign ram_MPORT_61_data = 24'h0;
  assign ram_MPORT_61_addr = 6'h3c;
  assign ram_MPORT_61_mask = 1'h1;
  assign ram_MPORT_61_en = reset;
  assign ram_MPORT_62_data = 24'h0;
  assign ram_MPORT_62_addr = 6'h3d;
  assign ram_MPORT_62_mask = 1'h1;
  assign ram_MPORT_62_en = reset;
  assign ram_MPORT_63_data = 24'h0;
  assign ram_MPORT_63_addr = 6'h3e;
  assign ram_MPORT_63_mask = 1'h1;
  assign ram_MPORT_63_en = reset;
  assign ram_MPORT_64_data = 24'h0;
  assign ram_MPORT_64_addr = 6'h3f;
  assign ram_MPORT_64_mask = 1'h1;
  assign ram_MPORT_64_en = reset;
  assign io_r_data_tag = _GEN_9[23:2];
  assign io_r_data_valid = _GEN_9[1];
  assign io_r_data_needFlush = _GEN_9[0];
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data;
    end
    if (ram_MPORT_1_en & ram_MPORT_1_mask) begin
      ram[ram_MPORT_1_addr] <= ram_MPORT_1_data;
    end
    if (ram_MPORT_2_en & ram_MPORT_2_mask) begin
      ram[ram_MPORT_2_addr] <= ram_MPORT_2_data;
    end
    if (ram_MPORT_3_en & ram_MPORT_3_mask) begin
      ram[ram_MPORT_3_addr] <= ram_MPORT_3_data;
    end
    if (ram_MPORT_4_en & ram_MPORT_4_mask) begin
      ram[ram_MPORT_4_addr] <= ram_MPORT_4_data;
    end
    if (ram_MPORT_5_en & ram_MPORT_5_mask) begin
      ram[ram_MPORT_5_addr] <= ram_MPORT_5_data;
    end
    if (ram_MPORT_6_en & ram_MPORT_6_mask) begin
      ram[ram_MPORT_6_addr] <= ram_MPORT_6_data;
    end
    if (ram_MPORT_7_en & ram_MPORT_7_mask) begin
      ram[ram_MPORT_7_addr] <= ram_MPORT_7_data;
    end
    if (ram_MPORT_8_en & ram_MPORT_8_mask) begin
      ram[ram_MPORT_8_addr] <= ram_MPORT_8_data;
    end
    if (ram_MPORT_9_en & ram_MPORT_9_mask) begin
      ram[ram_MPORT_9_addr] <= ram_MPORT_9_data;
    end
    if (ram_MPORT_10_en & ram_MPORT_10_mask) begin
      ram[ram_MPORT_10_addr] <= ram_MPORT_10_data;
    end
    if (ram_MPORT_11_en & ram_MPORT_11_mask) begin
      ram[ram_MPORT_11_addr] <= ram_MPORT_11_data;
    end
    if (ram_MPORT_12_en & ram_MPORT_12_mask) begin
      ram[ram_MPORT_12_addr] <= ram_MPORT_12_data;
    end
    if (ram_MPORT_13_en & ram_MPORT_13_mask) begin
      ram[ram_MPORT_13_addr] <= ram_MPORT_13_data;
    end
    if (ram_MPORT_14_en & ram_MPORT_14_mask) begin
      ram[ram_MPORT_14_addr] <= ram_MPORT_14_data;
    end
    if (ram_MPORT_15_en & ram_MPORT_15_mask) begin
      ram[ram_MPORT_15_addr] <= ram_MPORT_15_data;
    end
    if (ram_MPORT_16_en & ram_MPORT_16_mask) begin
      ram[ram_MPORT_16_addr] <= ram_MPORT_16_data;
    end
    if (ram_MPORT_17_en & ram_MPORT_17_mask) begin
      ram[ram_MPORT_17_addr] <= ram_MPORT_17_data;
    end
    if (ram_MPORT_18_en & ram_MPORT_18_mask) begin
      ram[ram_MPORT_18_addr] <= ram_MPORT_18_data;
    end
    if (ram_MPORT_19_en & ram_MPORT_19_mask) begin
      ram[ram_MPORT_19_addr] <= ram_MPORT_19_data;
    end
    if (ram_MPORT_20_en & ram_MPORT_20_mask) begin
      ram[ram_MPORT_20_addr] <= ram_MPORT_20_data;
    end
    if (ram_MPORT_21_en & ram_MPORT_21_mask) begin
      ram[ram_MPORT_21_addr] <= ram_MPORT_21_data;
    end
    if (ram_MPORT_22_en & ram_MPORT_22_mask) begin
      ram[ram_MPORT_22_addr] <= ram_MPORT_22_data;
    end
    if (ram_MPORT_23_en & ram_MPORT_23_mask) begin
      ram[ram_MPORT_23_addr] <= ram_MPORT_23_data;
    end
    if (ram_MPORT_24_en & ram_MPORT_24_mask) begin
      ram[ram_MPORT_24_addr] <= ram_MPORT_24_data;
    end
    if (ram_MPORT_25_en & ram_MPORT_25_mask) begin
      ram[ram_MPORT_25_addr] <= ram_MPORT_25_data;
    end
    if (ram_MPORT_26_en & ram_MPORT_26_mask) begin
      ram[ram_MPORT_26_addr] <= ram_MPORT_26_data;
    end
    if (ram_MPORT_27_en & ram_MPORT_27_mask) begin
      ram[ram_MPORT_27_addr] <= ram_MPORT_27_data;
    end
    if (ram_MPORT_28_en & ram_MPORT_28_mask) begin
      ram[ram_MPORT_28_addr] <= ram_MPORT_28_data;
    end
    if (ram_MPORT_29_en & ram_MPORT_29_mask) begin
      ram[ram_MPORT_29_addr] <= ram_MPORT_29_data;
    end
    if (ram_MPORT_30_en & ram_MPORT_30_mask) begin
      ram[ram_MPORT_30_addr] <= ram_MPORT_30_data;
    end
    if (ram_MPORT_31_en & ram_MPORT_31_mask) begin
      ram[ram_MPORT_31_addr] <= ram_MPORT_31_data;
    end
    if (ram_MPORT_32_en & ram_MPORT_32_mask) begin
      ram[ram_MPORT_32_addr] <= ram_MPORT_32_data;
    end
    if (ram_MPORT_33_en & ram_MPORT_33_mask) begin
      ram[ram_MPORT_33_addr] <= ram_MPORT_33_data;
    end
    if (ram_MPORT_34_en & ram_MPORT_34_mask) begin
      ram[ram_MPORT_34_addr] <= ram_MPORT_34_data;
    end
    if (ram_MPORT_35_en & ram_MPORT_35_mask) begin
      ram[ram_MPORT_35_addr] <= ram_MPORT_35_data;
    end
    if (ram_MPORT_36_en & ram_MPORT_36_mask) begin
      ram[ram_MPORT_36_addr] <= ram_MPORT_36_data;
    end
    if (ram_MPORT_37_en & ram_MPORT_37_mask) begin
      ram[ram_MPORT_37_addr] <= ram_MPORT_37_data;
    end
    if (ram_MPORT_38_en & ram_MPORT_38_mask) begin
      ram[ram_MPORT_38_addr] <= ram_MPORT_38_data;
    end
    if (ram_MPORT_39_en & ram_MPORT_39_mask) begin
      ram[ram_MPORT_39_addr] <= ram_MPORT_39_data;
    end
    if (ram_MPORT_40_en & ram_MPORT_40_mask) begin
      ram[ram_MPORT_40_addr] <= ram_MPORT_40_data;
    end
    if (ram_MPORT_41_en & ram_MPORT_41_mask) begin
      ram[ram_MPORT_41_addr] <= ram_MPORT_41_data;
    end
    if (ram_MPORT_42_en & ram_MPORT_42_mask) begin
      ram[ram_MPORT_42_addr] <= ram_MPORT_42_data;
    end
    if (ram_MPORT_43_en & ram_MPORT_43_mask) begin
      ram[ram_MPORT_43_addr] <= ram_MPORT_43_data;
    end
    if (ram_MPORT_44_en & ram_MPORT_44_mask) begin
      ram[ram_MPORT_44_addr] <= ram_MPORT_44_data;
    end
    if (ram_MPORT_45_en & ram_MPORT_45_mask) begin
      ram[ram_MPORT_45_addr] <= ram_MPORT_45_data;
    end
    if (ram_MPORT_46_en & ram_MPORT_46_mask) begin
      ram[ram_MPORT_46_addr] <= ram_MPORT_46_data;
    end
    if (ram_MPORT_47_en & ram_MPORT_47_mask) begin
      ram[ram_MPORT_47_addr] <= ram_MPORT_47_data;
    end
    if (ram_MPORT_48_en & ram_MPORT_48_mask) begin
      ram[ram_MPORT_48_addr] <= ram_MPORT_48_data;
    end
    if (ram_MPORT_49_en & ram_MPORT_49_mask) begin
      ram[ram_MPORT_49_addr] <= ram_MPORT_49_data;
    end
    if (ram_MPORT_50_en & ram_MPORT_50_mask) begin
      ram[ram_MPORT_50_addr] <= ram_MPORT_50_data;
    end
    if (ram_MPORT_51_en & ram_MPORT_51_mask) begin
      ram[ram_MPORT_51_addr] <= ram_MPORT_51_data;
    end
    if (ram_MPORT_52_en & ram_MPORT_52_mask) begin
      ram[ram_MPORT_52_addr] <= ram_MPORT_52_data;
    end
    if (ram_MPORT_53_en & ram_MPORT_53_mask) begin
      ram[ram_MPORT_53_addr] <= ram_MPORT_53_data;
    end
    if (ram_MPORT_54_en & ram_MPORT_54_mask) begin
      ram[ram_MPORT_54_addr] <= ram_MPORT_54_data;
    end
    if (ram_MPORT_55_en & ram_MPORT_55_mask) begin
      ram[ram_MPORT_55_addr] <= ram_MPORT_55_data;
    end
    if (ram_MPORT_56_en & ram_MPORT_56_mask) begin
      ram[ram_MPORT_56_addr] <= ram_MPORT_56_data;
    end
    if (ram_MPORT_57_en & ram_MPORT_57_mask) begin
      ram[ram_MPORT_57_addr] <= ram_MPORT_57_data;
    end
    if (ram_MPORT_58_en & ram_MPORT_58_mask) begin
      ram[ram_MPORT_58_addr] <= ram_MPORT_58_data;
    end
    if (ram_MPORT_59_en & ram_MPORT_59_mask) begin
      ram[ram_MPORT_59_addr] <= ram_MPORT_59_data;
    end
    if (ram_MPORT_60_en & ram_MPORT_60_mask) begin
      ram[ram_MPORT_60_addr] <= ram_MPORT_60_data;
    end
    if (ram_MPORT_61_en & ram_MPORT_61_mask) begin
      ram[ram_MPORT_61_addr] <= ram_MPORT_61_data;
    end
    if (ram_MPORT_62_en & ram_MPORT_62_mask) begin
      ram[ram_MPORT_62_addr] <= ram_MPORT_62_data;
    end
    if (ram_MPORT_63_en & ram_MPORT_63_mask) begin
      ram[ram_MPORT_63_addr] <= ram_MPORT_63_data;
    end
    if (ram_MPORT_64_en & ram_MPORT_64_mask) begin
      ram[ram_MPORT_64_addr] <= ram_MPORT_64_data;
    end
    ram_rdata_MPORT_en_pipe_0 <= io_r_ren & _realRen_T;
    if (io_r_ren & _realRen_T) begin
      ram_rdata_MPORT_addr_pipe_0 <= io_r_setIdx;
    end
    rdata_REG <= io_r_ren & ~io_w_wen;
    if (reset) begin
      rdata_r <= 24'h0;
    end else if (rdata_REG) begin
      rdata_r <= ram_rdata_MPORT_data;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[23:0];
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_rdata_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  rdata_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rdata_r = _RAND_4[23:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_findingBlock(
  input        io_inWayValid_0,
  input        io_inWayValid_1,
  input  [1:0] io_inIdx_0,
  input  [1:0] io_inIdx_1,
  input  [1:0] io_inValue_0,
  input  [1:0] io_inValue_1,
  output       io_outWayValid,
  output [1:0] io_outIdx,
  output [1:0] io_outValue
);
  wire  _available_T = ~io_inWayValid_0;
  wire  available = ~io_inWayValid_0 | ~io_inWayValid_1;
  wire  compare = io_inValue_0 > io_inValue_1;
  wire [1:0] idxCompare = compare ? io_inIdx_0 : io_inIdx_1;
  wire [1:0] _io_outIdx_T_1 = _available_T ? io_inIdx_0 : io_inIdx_1;
  assign io_outWayValid = ~available;
  assign io_outIdx = available ? _io_outIdx_T_1 : idxCompare;
  assign io_outValue = compare ? io_inValue_0 : io_inValue_1;
endmodule
module ysyx_040656_LRU(
  input        io_inWayValid_0,
  input        io_inWayValid_1,
  input        io_inWayValid_2,
  input        io_inWayValid_3,
  input  [1:0] io_inValue_0,
  input  [1:0] io_inValue_1,
  input  [1:0] io_inValue_2,
  input  [1:0] io_inValue_3,
  output [1:0] io_outIdx
);
  wire  Lut_0_0_io_inWayValid_0;
  wire  Lut_0_0_io_inWayValid_1;
  wire [1:0] Lut_0_0_io_inIdx_0;
  wire [1:0] Lut_0_0_io_inIdx_1;
  wire [1:0] Lut_0_0_io_inValue_0;
  wire [1:0] Lut_0_0_io_inValue_1;
  wire  Lut_0_0_io_outWayValid;
  wire [1:0] Lut_0_0_io_outIdx;
  wire [1:0] Lut_0_0_io_outValue;
  wire  Lut_1_0_io_inWayValid_0;
  wire  Lut_1_0_io_inWayValid_1;
  wire [1:0] Lut_1_0_io_inIdx_0;
  wire [1:0] Lut_1_0_io_inIdx_1;
  wire [1:0] Lut_1_0_io_inValue_0;
  wire [1:0] Lut_1_0_io_inValue_1;
  wire  Lut_1_0_io_outWayValid;
  wire [1:0] Lut_1_0_io_outIdx;
  wire [1:0] Lut_1_0_io_outValue;
  wire  Lut_1_1_io_inWayValid_0;
  wire  Lut_1_1_io_inWayValid_1;
  wire [1:0] Lut_1_1_io_inIdx_0;
  wire [1:0] Lut_1_1_io_inIdx_1;
  wire [1:0] Lut_1_1_io_inValue_0;
  wire [1:0] Lut_1_1_io_inValue_1;
  wire  Lut_1_1_io_outWayValid;
  wire [1:0] Lut_1_1_io_outIdx;
  wire [1:0] Lut_1_1_io_outValue;
  ysyx_040656_findingBlock Lut_0_0 (
    .io_inWayValid_0(Lut_0_0_io_inWayValid_0),
    .io_inWayValid_1(Lut_0_0_io_inWayValid_1),
    .io_inIdx_0(Lut_0_0_io_inIdx_0),
    .io_inIdx_1(Lut_0_0_io_inIdx_1),
    .io_inValue_0(Lut_0_0_io_inValue_0),
    .io_inValue_1(Lut_0_0_io_inValue_1),
    .io_outWayValid(Lut_0_0_io_outWayValid),
    .io_outIdx(Lut_0_0_io_outIdx),
    .io_outValue(Lut_0_0_io_outValue)
  );
  ysyx_040656_findingBlock Lut_1_0 (
    .io_inWayValid_0(Lut_1_0_io_inWayValid_0),
    .io_inWayValid_1(Lut_1_0_io_inWayValid_1),
    .io_inIdx_0(Lut_1_0_io_inIdx_0),
    .io_inIdx_1(Lut_1_0_io_inIdx_1),
    .io_inValue_0(Lut_1_0_io_inValue_0),
    .io_inValue_1(Lut_1_0_io_inValue_1),
    .io_outWayValid(Lut_1_0_io_outWayValid),
    .io_outIdx(Lut_1_0_io_outIdx),
    .io_outValue(Lut_1_0_io_outValue)
  );
  ysyx_040656_findingBlock Lut_1_1 (
    .io_inWayValid_0(Lut_1_1_io_inWayValid_0),
    .io_inWayValid_1(Lut_1_1_io_inWayValid_1),
    .io_inIdx_0(Lut_1_1_io_inIdx_0),
    .io_inIdx_1(Lut_1_1_io_inIdx_1),
    .io_inValue_0(Lut_1_1_io_inValue_0),
    .io_inValue_1(Lut_1_1_io_inValue_1),
    .io_outWayValid(Lut_1_1_io_outWayValid),
    .io_outIdx(Lut_1_1_io_outIdx),
    .io_outValue(Lut_1_1_io_outValue)
  );
  assign io_outIdx = Lut_0_0_io_outIdx;
  assign Lut_0_0_io_inWayValid_0 = Lut_1_0_io_outWayValid;
  assign Lut_0_0_io_inWayValid_1 = Lut_1_1_io_outWayValid;
  assign Lut_0_0_io_inIdx_0 = Lut_1_0_io_outIdx;
  assign Lut_0_0_io_inIdx_1 = Lut_1_1_io_outIdx;
  assign Lut_0_0_io_inValue_0 = Lut_1_0_io_outValue;
  assign Lut_0_0_io_inValue_1 = Lut_1_1_io_outValue;
  assign Lut_1_0_io_inWayValid_0 = io_inWayValid_0;
  assign Lut_1_0_io_inWayValid_1 = io_inWayValid_1;
  assign Lut_1_0_io_inIdx_0 = 2'h0;
  assign Lut_1_0_io_inIdx_1 = 2'h1;
  assign Lut_1_0_io_inValue_0 = io_inValue_0;
  assign Lut_1_0_io_inValue_1 = io_inValue_1;
  assign Lut_1_1_io_inWayValid_0 = io_inWayValid_2;
  assign Lut_1_1_io_inWayValid_1 = io_inWayValid_3;
  assign Lut_1_1_io_inIdx_0 = 2'h2;
  assign Lut_1_1_io_inIdx_1 = 2'h3;
  assign Lut_1_1_io_inValue_0 = io_inValue_2;
  assign Lut_1_1_io_inValue_1 = io_inValue_3;
endmodule
module ysyx_040656_ICache(
  input          clock,
  input          reset,
  output         io_in_req_ready,
  input  [31:0]  io_in_req_bits_addr,
  input          io_in_resp_ready,
  output         io_in_resp_valid,
  output [31:0]  io_in_resp_bits_rdata,
  input          io_out_req_ready,
  output         io_out_req_valid,
  output [31:0]  io_out_req_bits_addr,
  output [127:0] io_out_req_bits_wdata,
  output [2:0]   io_out_req_bits_cmd,
  output         io_out_resp_ready,
  input          io_out_resp_valid,
  input  [127:0] io_out_resp_bits_rdata,
  input          io_mmio_req_ready,
  output         io_mmio_req_valid,
  output [31:0]  io_mmio_req_bits_addr,
  output [1:0]   io_mmio_req_bits_size,
  output         io_mmio_resp_ready,
  input          io_mmio_resp_valid,
  input  [63:0]  io_mmio_resp_bits_rdata,
  input  [127:0] io_dataArray_0_rdata,
  output         io_dataArray_0_wen,
  output [5:0]   io_dataArray_0_addr,
  output [127:0] io_dataArray_0_wdata,
  input  [127:0] io_dataArray_1_rdata,
  output         io_dataArray_1_wen,
  output [5:0]   io_dataArray_1_addr,
  output [127:0] io_dataArray_1_wdata,
  input  [127:0] io_dataArray_2_rdata,
  output         io_dataArray_2_wen,
  output [5:0]   io_dataArray_2_addr,
  output [127:0] io_dataArray_2_wdata,
  input  [127:0] io_dataArray_3_rdata,
  output         io_dataArray_3_wen,
  output [5:0]   io_dataArray_3_addr,
  output [127:0] io_dataArray_3_wdata,
  input          difftestFENCEI
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [63:0] _RAND_261;
`endif
  wire  metaArray_0_clock;
  wire  metaArray_0_reset;
  wire [5:0] metaArray_0_io_w_setIdx;
  wire [21:0] metaArray_0_io_w_data_tag;
  wire  metaArray_0_io_w_data_valid;
  wire  metaArray_0_io_w_data_needFlush;
  wire  metaArray_0_io_w_wen;
  wire [5:0] metaArray_0_io_r_setIdx;
  wire [21:0] metaArray_0_io_r_data_tag;
  wire  metaArray_0_io_r_data_valid;
  wire  metaArray_0_io_r_data_needFlush;
  wire  metaArray_0_io_r_ren;
  wire  metaArray_1_clock;
  wire  metaArray_1_reset;
  wire [5:0] metaArray_1_io_w_setIdx;
  wire [21:0] metaArray_1_io_w_data_tag;
  wire  metaArray_1_io_w_data_valid;
  wire  metaArray_1_io_w_data_needFlush;
  wire  metaArray_1_io_w_wen;
  wire [5:0] metaArray_1_io_r_setIdx;
  wire [21:0] metaArray_1_io_r_data_tag;
  wire  metaArray_1_io_r_data_valid;
  wire  metaArray_1_io_r_data_needFlush;
  wire  metaArray_1_io_r_ren;
  wire  metaArray_2_clock;
  wire  metaArray_2_reset;
  wire [5:0] metaArray_2_io_w_setIdx;
  wire [21:0] metaArray_2_io_w_data_tag;
  wire  metaArray_2_io_w_data_valid;
  wire  metaArray_2_io_w_data_needFlush;
  wire  metaArray_2_io_w_wen;
  wire [5:0] metaArray_2_io_r_setIdx;
  wire [21:0] metaArray_2_io_r_data_tag;
  wire  metaArray_2_io_r_data_valid;
  wire  metaArray_2_io_r_data_needFlush;
  wire  metaArray_2_io_r_ren;
  wire  metaArray_3_clock;
  wire  metaArray_3_reset;
  wire [5:0] metaArray_3_io_w_setIdx;
  wire [21:0] metaArray_3_io_w_data_tag;
  wire  metaArray_3_io_w_data_valid;
  wire  metaArray_3_io_w_data_needFlush;
  wire  metaArray_3_io_w_wen;
  wire [5:0] metaArray_3_io_r_setIdx;
  wire [21:0] metaArray_3_io_r_data_tag;
  wire  metaArray_3_io_r_data_valid;
  wire  metaArray_3_io_r_data_needFlush;
  wire  metaArray_3_io_r_ren;
  wire  selTree_io_inWayValid_0;
  wire  selTree_io_inWayValid_1;
  wire  selTree_io_inWayValid_2;
  wire  selTree_io_inWayValid_3;
  wire [1:0] selTree_io_inValue_0;
  wire [1:0] selTree_io_inValue_1;
  wire [1:0] selTree_io_inValue_2;
  wire [1:0] selTree_io_inValue_3;
  wire [1:0] selTree_io_outIdx;
  reg [2:0] icache_status;
  reg [1:0] regCount_0_0;
  reg [1:0] regCount_0_1;
  reg [1:0] regCount_0_2;
  reg [1:0] regCount_0_3;
  reg [1:0] regCount_1_0;
  reg [1:0] regCount_1_1;
  reg [1:0] regCount_1_2;
  reg [1:0] regCount_1_3;
  reg [1:0] regCount_2_0;
  reg [1:0] regCount_2_1;
  reg [1:0] regCount_2_2;
  reg [1:0] regCount_2_3;
  reg [1:0] regCount_3_0;
  reg [1:0] regCount_3_1;
  reg [1:0] regCount_3_2;
  reg [1:0] regCount_3_3;
  reg [1:0] regCount_4_0;
  reg [1:0] regCount_4_1;
  reg [1:0] regCount_4_2;
  reg [1:0] regCount_4_3;
  reg [1:0] regCount_5_0;
  reg [1:0] regCount_5_1;
  reg [1:0] regCount_5_2;
  reg [1:0] regCount_5_3;
  reg [1:0] regCount_6_0;
  reg [1:0] regCount_6_1;
  reg [1:0] regCount_6_2;
  reg [1:0] regCount_6_3;
  reg [1:0] regCount_7_0;
  reg [1:0] regCount_7_1;
  reg [1:0] regCount_7_2;
  reg [1:0] regCount_7_3;
  reg [1:0] regCount_8_0;
  reg [1:0] regCount_8_1;
  reg [1:0] regCount_8_2;
  reg [1:0] regCount_8_3;
  reg [1:0] regCount_9_0;
  reg [1:0] regCount_9_1;
  reg [1:0] regCount_9_2;
  reg [1:0] regCount_9_3;
  reg [1:0] regCount_10_0;
  reg [1:0] regCount_10_1;
  reg [1:0] regCount_10_2;
  reg [1:0] regCount_10_3;
  reg [1:0] regCount_11_0;
  reg [1:0] regCount_11_1;
  reg [1:0] regCount_11_2;
  reg [1:0] regCount_11_3;
  reg [1:0] regCount_12_0;
  reg [1:0] regCount_12_1;
  reg [1:0] regCount_12_2;
  reg [1:0] regCount_12_3;
  reg [1:0] regCount_13_0;
  reg [1:0] regCount_13_1;
  reg [1:0] regCount_13_2;
  reg [1:0] regCount_13_3;
  reg [1:0] regCount_14_0;
  reg [1:0] regCount_14_1;
  reg [1:0] regCount_14_2;
  reg [1:0] regCount_14_3;
  reg [1:0] regCount_15_0;
  reg [1:0] regCount_15_1;
  reg [1:0] regCount_15_2;
  reg [1:0] regCount_15_3;
  reg [1:0] regCount_16_0;
  reg [1:0] regCount_16_1;
  reg [1:0] regCount_16_2;
  reg [1:0] regCount_16_3;
  reg [1:0] regCount_17_0;
  reg [1:0] regCount_17_1;
  reg [1:0] regCount_17_2;
  reg [1:0] regCount_17_3;
  reg [1:0] regCount_18_0;
  reg [1:0] regCount_18_1;
  reg [1:0] regCount_18_2;
  reg [1:0] regCount_18_3;
  reg [1:0] regCount_19_0;
  reg [1:0] regCount_19_1;
  reg [1:0] regCount_19_2;
  reg [1:0] regCount_19_3;
  reg [1:0] regCount_20_0;
  reg [1:0] regCount_20_1;
  reg [1:0] regCount_20_2;
  reg [1:0] regCount_20_3;
  reg [1:0] regCount_21_0;
  reg [1:0] regCount_21_1;
  reg [1:0] regCount_21_2;
  reg [1:0] regCount_21_3;
  reg [1:0] regCount_22_0;
  reg [1:0] regCount_22_1;
  reg [1:0] regCount_22_2;
  reg [1:0] regCount_22_3;
  reg [1:0] regCount_23_0;
  reg [1:0] regCount_23_1;
  reg [1:0] regCount_23_2;
  reg [1:0] regCount_23_3;
  reg [1:0] regCount_24_0;
  reg [1:0] regCount_24_1;
  reg [1:0] regCount_24_2;
  reg [1:0] regCount_24_3;
  reg [1:0] regCount_25_0;
  reg [1:0] regCount_25_1;
  reg [1:0] regCount_25_2;
  reg [1:0] regCount_25_3;
  reg [1:0] regCount_26_0;
  reg [1:0] regCount_26_1;
  reg [1:0] regCount_26_2;
  reg [1:0] regCount_26_3;
  reg [1:0] regCount_27_0;
  reg [1:0] regCount_27_1;
  reg [1:0] regCount_27_2;
  reg [1:0] regCount_27_3;
  reg [1:0] regCount_28_0;
  reg [1:0] regCount_28_1;
  reg [1:0] regCount_28_2;
  reg [1:0] regCount_28_3;
  reg [1:0] regCount_29_0;
  reg [1:0] regCount_29_1;
  reg [1:0] regCount_29_2;
  reg [1:0] regCount_29_3;
  reg [1:0] regCount_30_0;
  reg [1:0] regCount_30_1;
  reg [1:0] regCount_30_2;
  reg [1:0] regCount_30_3;
  reg [1:0] regCount_31_0;
  reg [1:0] regCount_31_1;
  reg [1:0] regCount_31_2;
  reg [1:0] regCount_31_3;
  reg [1:0] regCount_32_0;
  reg [1:0] regCount_32_1;
  reg [1:0] regCount_32_2;
  reg [1:0] regCount_32_3;
  reg [1:0] regCount_33_0;
  reg [1:0] regCount_33_1;
  reg [1:0] regCount_33_2;
  reg [1:0] regCount_33_3;
  reg [1:0] regCount_34_0;
  reg [1:0] regCount_34_1;
  reg [1:0] regCount_34_2;
  reg [1:0] regCount_34_3;
  reg [1:0] regCount_35_0;
  reg [1:0] regCount_35_1;
  reg [1:0] regCount_35_2;
  reg [1:0] regCount_35_3;
  reg [1:0] regCount_36_0;
  reg [1:0] regCount_36_1;
  reg [1:0] regCount_36_2;
  reg [1:0] regCount_36_3;
  reg [1:0] regCount_37_0;
  reg [1:0] regCount_37_1;
  reg [1:0] regCount_37_2;
  reg [1:0] regCount_37_3;
  reg [1:0] regCount_38_0;
  reg [1:0] regCount_38_1;
  reg [1:0] regCount_38_2;
  reg [1:0] regCount_38_3;
  reg [1:0] regCount_39_0;
  reg [1:0] regCount_39_1;
  reg [1:0] regCount_39_2;
  reg [1:0] regCount_39_3;
  reg [1:0] regCount_40_0;
  reg [1:0] regCount_40_1;
  reg [1:0] regCount_40_2;
  reg [1:0] regCount_40_3;
  reg [1:0] regCount_41_0;
  reg [1:0] regCount_41_1;
  reg [1:0] regCount_41_2;
  reg [1:0] regCount_41_3;
  reg [1:0] regCount_42_0;
  reg [1:0] regCount_42_1;
  reg [1:0] regCount_42_2;
  reg [1:0] regCount_42_3;
  reg [1:0] regCount_43_0;
  reg [1:0] regCount_43_1;
  reg [1:0] regCount_43_2;
  reg [1:0] regCount_43_3;
  reg [1:0] regCount_44_0;
  reg [1:0] regCount_44_1;
  reg [1:0] regCount_44_2;
  reg [1:0] regCount_44_3;
  reg [1:0] regCount_45_0;
  reg [1:0] regCount_45_1;
  reg [1:0] regCount_45_2;
  reg [1:0] regCount_45_3;
  reg [1:0] regCount_46_0;
  reg [1:0] regCount_46_1;
  reg [1:0] regCount_46_2;
  reg [1:0] regCount_46_3;
  reg [1:0] regCount_47_0;
  reg [1:0] regCount_47_1;
  reg [1:0] regCount_47_2;
  reg [1:0] regCount_47_3;
  reg [1:0] regCount_48_0;
  reg [1:0] regCount_48_1;
  reg [1:0] regCount_48_2;
  reg [1:0] regCount_48_3;
  reg [1:0] regCount_49_0;
  reg [1:0] regCount_49_1;
  reg [1:0] regCount_49_2;
  reg [1:0] regCount_49_3;
  reg [1:0] regCount_50_0;
  reg [1:0] regCount_50_1;
  reg [1:0] regCount_50_2;
  reg [1:0] regCount_50_3;
  reg [1:0] regCount_51_0;
  reg [1:0] regCount_51_1;
  reg [1:0] regCount_51_2;
  reg [1:0] regCount_51_3;
  reg [1:0] regCount_52_0;
  reg [1:0] regCount_52_1;
  reg [1:0] regCount_52_2;
  reg [1:0] regCount_52_3;
  reg [1:0] regCount_53_0;
  reg [1:0] regCount_53_1;
  reg [1:0] regCount_53_2;
  reg [1:0] regCount_53_3;
  reg [1:0] regCount_54_0;
  reg [1:0] regCount_54_1;
  reg [1:0] regCount_54_2;
  reg [1:0] regCount_54_3;
  reg [1:0] regCount_55_0;
  reg [1:0] regCount_55_1;
  reg [1:0] regCount_55_2;
  reg [1:0] regCount_55_3;
  reg [1:0] regCount_56_0;
  reg [1:0] regCount_56_1;
  reg [1:0] regCount_56_2;
  reg [1:0] regCount_56_3;
  reg [1:0] regCount_57_0;
  reg [1:0] regCount_57_1;
  reg [1:0] regCount_57_2;
  reg [1:0] regCount_57_3;
  reg [1:0] regCount_58_0;
  reg [1:0] regCount_58_1;
  reg [1:0] regCount_58_2;
  reg [1:0] regCount_58_3;
  reg [1:0] regCount_59_0;
  reg [1:0] regCount_59_1;
  reg [1:0] regCount_59_2;
  reg [1:0] regCount_59_3;
  reg [1:0] regCount_60_0;
  reg [1:0] regCount_60_1;
  reg [1:0] regCount_60_2;
  reg [1:0] regCount_60_3;
  reg [1:0] regCount_61_0;
  reg [1:0] regCount_61_1;
  reg [1:0] regCount_61_2;
  reg [1:0] regCount_61_3;
  reg [1:0] regCount_62_0;
  reg [1:0] regCount_62_1;
  reg [1:0] regCount_62_2;
  reg [1:0] regCount_62_3;
  reg [1:0] regCount_63_0;
  reg [1:0] regCount_63_1;
  reg [1:0] regCount_63_2;
  reg [1:0] regCount_63_3;
  wire  s1_isMMIO_selVec_0 = io_in_req_bits_addr <= 32'h1ffffff;
  wire  s1_isMMIO_selVec_1 = io_in_req_bits_addr >= 32'h2000000 & io_in_req_bits_addr <= 32'h200ffff;
  wire  s1_isMMIO_selVec_2 = io_in_req_bits_addr >= 32'h2010000 & io_in_req_bits_addr <= 32'h7fffffff;
  wire  s1_isMMIO_selVec_3 = io_in_req_bits_addr >= 32'hfc000000;
  wire [3:0] _s1_isMMIO_hit_T = {s1_isMMIO_selVec_3,s1_isMMIO_selVec_2,s1_isMMIO_selVec_1,s1_isMMIO_selVec_0};
  wire  s1_isMMIO_hit = |_s1_isMMIO_hit_T;
  wire [63:0] dataWays_0_0 = io_dataArray_0_rdata[63:0];
  wire [63:0] dataWays_0_1 = io_dataArray_0_rdata[127:64];
  wire [63:0] dataWays_1_0 = io_dataArray_1_rdata[63:0];
  wire [63:0] dataWays_1_1 = io_dataArray_1_rdata[127:64];
  wire [63:0] dataWays_2_0 = io_dataArray_2_rdata[63:0];
  wire [63:0] dataWays_2_1 = io_dataArray_2_rdata[127:64];
  wire [63:0] dataWays_3_0 = io_dataArray_3_rdata[63:0];
  wire [63:0] dataWays_3_1 = io_dataArray_3_rdata[127:64];
  reg  s2_pipeline_valid;
  reg [31:0] s2_pipeline_addr;
  reg [1:0] s2_pipeline_size;
  reg  s2_pipeline_isMMIO;
  wire  _s2_stall_T = io_in_resp_ready & io_in_resp_valid;
  wire  s2_stall = s2_pipeline_valid & ~_s2_stall_T;
  wire  _T_15 = ~s2_stall;
  wire  _GEN_4 = ~s2_stall | s2_pipeline_valid;
  wire [21:0] metaWays_0_tag = metaArray_0_io_r_data_tag;
  wire  metaWays_0_valid = metaArray_0_io_r_data_valid;
  wire  hitVec_0 = metaWays_0_valid & metaWays_0_tag == s2_pipeline_addr[31:10];
  wire [1:0] _GEN_9 = 6'h1 == s2_pipeline_addr[9:4] ? regCount_1_0 : regCount_0_0;
  wire [1:0] _GEN_10 = 6'h2 == s2_pipeline_addr[9:4] ? regCount_2_0 : _GEN_9;
  wire [1:0] _GEN_11 = 6'h3 == s2_pipeline_addr[9:4] ? regCount_3_0 : _GEN_10;
  wire [1:0] _GEN_12 = 6'h4 == s2_pipeline_addr[9:4] ? regCount_4_0 : _GEN_11;
  wire [1:0] _GEN_13 = 6'h5 == s2_pipeline_addr[9:4] ? regCount_5_0 : _GEN_12;
  wire [1:0] _GEN_14 = 6'h6 == s2_pipeline_addr[9:4] ? regCount_6_0 : _GEN_13;
  wire [1:0] _GEN_15 = 6'h7 == s2_pipeline_addr[9:4] ? regCount_7_0 : _GEN_14;
  wire [1:0] _GEN_16 = 6'h8 == s2_pipeline_addr[9:4] ? regCount_8_0 : _GEN_15;
  wire [1:0] _GEN_17 = 6'h9 == s2_pipeline_addr[9:4] ? regCount_9_0 : _GEN_16;
  wire [1:0] _GEN_18 = 6'ha == s2_pipeline_addr[9:4] ? regCount_10_0 : _GEN_17;
  wire [1:0] _GEN_19 = 6'hb == s2_pipeline_addr[9:4] ? regCount_11_0 : _GEN_18;
  wire [1:0] _GEN_20 = 6'hc == s2_pipeline_addr[9:4] ? regCount_12_0 : _GEN_19;
  wire [1:0] _GEN_21 = 6'hd == s2_pipeline_addr[9:4] ? regCount_13_0 : _GEN_20;
  wire [1:0] _GEN_22 = 6'he == s2_pipeline_addr[9:4] ? regCount_14_0 : _GEN_21;
  wire [1:0] _GEN_23 = 6'hf == s2_pipeline_addr[9:4] ? regCount_15_0 : _GEN_22;
  wire [1:0] _GEN_24 = 6'h10 == s2_pipeline_addr[9:4] ? regCount_16_0 : _GEN_23;
  wire [1:0] _GEN_25 = 6'h11 == s2_pipeline_addr[9:4] ? regCount_17_0 : _GEN_24;
  wire [1:0] _GEN_26 = 6'h12 == s2_pipeline_addr[9:4] ? regCount_18_0 : _GEN_25;
  wire [1:0] _GEN_27 = 6'h13 == s2_pipeline_addr[9:4] ? regCount_19_0 : _GEN_26;
  wire [1:0] _GEN_28 = 6'h14 == s2_pipeline_addr[9:4] ? regCount_20_0 : _GEN_27;
  wire [1:0] _GEN_29 = 6'h15 == s2_pipeline_addr[9:4] ? regCount_21_0 : _GEN_28;
  wire [1:0] _GEN_30 = 6'h16 == s2_pipeline_addr[9:4] ? regCount_22_0 : _GEN_29;
  wire [1:0] _GEN_31 = 6'h17 == s2_pipeline_addr[9:4] ? regCount_23_0 : _GEN_30;
  wire [1:0] _GEN_32 = 6'h18 == s2_pipeline_addr[9:4] ? regCount_24_0 : _GEN_31;
  wire [1:0] _GEN_33 = 6'h19 == s2_pipeline_addr[9:4] ? regCount_25_0 : _GEN_32;
  wire [1:0] _GEN_34 = 6'h1a == s2_pipeline_addr[9:4] ? regCount_26_0 : _GEN_33;
  wire [1:0] _GEN_35 = 6'h1b == s2_pipeline_addr[9:4] ? regCount_27_0 : _GEN_34;
  wire [1:0] _GEN_36 = 6'h1c == s2_pipeline_addr[9:4] ? regCount_28_0 : _GEN_35;
  wire [1:0] _GEN_37 = 6'h1d == s2_pipeline_addr[9:4] ? regCount_29_0 : _GEN_36;
  wire [1:0] _GEN_38 = 6'h1e == s2_pipeline_addr[9:4] ? regCount_30_0 : _GEN_37;
  wire [1:0] _GEN_39 = 6'h1f == s2_pipeline_addr[9:4] ? regCount_31_0 : _GEN_38;
  wire [1:0] _GEN_40 = 6'h20 == s2_pipeline_addr[9:4] ? regCount_32_0 : _GEN_39;
  wire [1:0] _GEN_41 = 6'h21 == s2_pipeline_addr[9:4] ? regCount_33_0 : _GEN_40;
  wire [1:0] _GEN_42 = 6'h22 == s2_pipeline_addr[9:4] ? regCount_34_0 : _GEN_41;
  wire [1:0] _GEN_43 = 6'h23 == s2_pipeline_addr[9:4] ? regCount_35_0 : _GEN_42;
  wire [1:0] _GEN_44 = 6'h24 == s2_pipeline_addr[9:4] ? regCount_36_0 : _GEN_43;
  wire [1:0] _GEN_45 = 6'h25 == s2_pipeline_addr[9:4] ? regCount_37_0 : _GEN_44;
  wire [1:0] _GEN_46 = 6'h26 == s2_pipeline_addr[9:4] ? regCount_38_0 : _GEN_45;
  wire [1:0] _GEN_47 = 6'h27 == s2_pipeline_addr[9:4] ? regCount_39_0 : _GEN_46;
  wire [1:0] _GEN_48 = 6'h28 == s2_pipeline_addr[9:4] ? regCount_40_0 : _GEN_47;
  wire [1:0] _GEN_49 = 6'h29 == s2_pipeline_addr[9:4] ? regCount_41_0 : _GEN_48;
  wire [1:0] _GEN_50 = 6'h2a == s2_pipeline_addr[9:4] ? regCount_42_0 : _GEN_49;
  wire [1:0] _GEN_51 = 6'h2b == s2_pipeline_addr[9:4] ? regCount_43_0 : _GEN_50;
  wire [1:0] _GEN_52 = 6'h2c == s2_pipeline_addr[9:4] ? regCount_44_0 : _GEN_51;
  wire [1:0] _GEN_53 = 6'h2d == s2_pipeline_addr[9:4] ? regCount_45_0 : _GEN_52;
  wire [1:0] _GEN_54 = 6'h2e == s2_pipeline_addr[9:4] ? regCount_46_0 : _GEN_53;
  wire [1:0] _GEN_55 = 6'h2f == s2_pipeline_addr[9:4] ? regCount_47_0 : _GEN_54;
  wire [1:0] _GEN_56 = 6'h30 == s2_pipeline_addr[9:4] ? regCount_48_0 : _GEN_55;
  wire [1:0] _GEN_57 = 6'h31 == s2_pipeline_addr[9:4] ? regCount_49_0 : _GEN_56;
  wire [1:0] _GEN_58 = 6'h32 == s2_pipeline_addr[9:4] ? regCount_50_0 : _GEN_57;
  wire [1:0] _GEN_59 = 6'h33 == s2_pipeline_addr[9:4] ? regCount_51_0 : _GEN_58;
  wire [1:0] _GEN_60 = 6'h34 == s2_pipeline_addr[9:4] ? regCount_52_0 : _GEN_59;
  wire [1:0] _GEN_61 = 6'h35 == s2_pipeline_addr[9:4] ? regCount_53_0 : _GEN_60;
  wire [1:0] _GEN_62 = 6'h36 == s2_pipeline_addr[9:4] ? regCount_54_0 : _GEN_61;
  wire [1:0] _GEN_63 = 6'h37 == s2_pipeline_addr[9:4] ? regCount_55_0 : _GEN_62;
  wire [1:0] _GEN_64 = 6'h38 == s2_pipeline_addr[9:4] ? regCount_56_0 : _GEN_63;
  wire [1:0] _GEN_65 = 6'h39 == s2_pipeline_addr[9:4] ? regCount_57_0 : _GEN_64;
  wire [1:0] _GEN_66 = 6'h3a == s2_pipeline_addr[9:4] ? regCount_58_0 : _GEN_65;
  wire [1:0] _GEN_67 = 6'h3b == s2_pipeline_addr[9:4] ? regCount_59_0 : _GEN_66;
  wire [1:0] _GEN_68 = 6'h3c == s2_pipeline_addr[9:4] ? regCount_60_0 : _GEN_67;
  wire [1:0] _GEN_69 = 6'h3d == s2_pipeline_addr[9:4] ? regCount_61_0 : _GEN_68;
  wire [1:0] _GEN_70 = 6'h3e == s2_pipeline_addr[9:4] ? regCount_62_0 : _GEN_69;
  wire [1:0] _GEN_71 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_0 : _GEN_70;
  wire [21:0] metaWays_1_tag = metaArray_1_io_r_data_tag;
  wire  metaWays_1_valid = metaArray_1_io_r_data_valid;
  wire  hitVec_1 = metaWays_1_valid & metaWays_1_tag == s2_pipeline_addr[31:10];
  wire [1:0] _GEN_73 = 6'h1 == s2_pipeline_addr[9:4] ? regCount_1_1 : regCount_0_1;
  wire [1:0] _GEN_74 = 6'h2 == s2_pipeline_addr[9:4] ? regCount_2_1 : _GEN_73;
  wire [1:0] _GEN_75 = 6'h3 == s2_pipeline_addr[9:4] ? regCount_3_1 : _GEN_74;
  wire [1:0] _GEN_76 = 6'h4 == s2_pipeline_addr[9:4] ? regCount_4_1 : _GEN_75;
  wire [1:0] _GEN_77 = 6'h5 == s2_pipeline_addr[9:4] ? regCount_5_1 : _GEN_76;
  wire [1:0] _GEN_78 = 6'h6 == s2_pipeline_addr[9:4] ? regCount_6_1 : _GEN_77;
  wire [1:0] _GEN_79 = 6'h7 == s2_pipeline_addr[9:4] ? regCount_7_1 : _GEN_78;
  wire [1:0] _GEN_80 = 6'h8 == s2_pipeline_addr[9:4] ? regCount_8_1 : _GEN_79;
  wire [1:0] _GEN_81 = 6'h9 == s2_pipeline_addr[9:4] ? regCount_9_1 : _GEN_80;
  wire [1:0] _GEN_82 = 6'ha == s2_pipeline_addr[9:4] ? regCount_10_1 : _GEN_81;
  wire [1:0] _GEN_83 = 6'hb == s2_pipeline_addr[9:4] ? regCount_11_1 : _GEN_82;
  wire [1:0] _GEN_84 = 6'hc == s2_pipeline_addr[9:4] ? regCount_12_1 : _GEN_83;
  wire [1:0] _GEN_85 = 6'hd == s2_pipeline_addr[9:4] ? regCount_13_1 : _GEN_84;
  wire [1:0] _GEN_86 = 6'he == s2_pipeline_addr[9:4] ? regCount_14_1 : _GEN_85;
  wire [1:0] _GEN_87 = 6'hf == s2_pipeline_addr[9:4] ? regCount_15_1 : _GEN_86;
  wire [1:0] _GEN_88 = 6'h10 == s2_pipeline_addr[9:4] ? regCount_16_1 : _GEN_87;
  wire [1:0] _GEN_89 = 6'h11 == s2_pipeline_addr[9:4] ? regCount_17_1 : _GEN_88;
  wire [1:0] _GEN_90 = 6'h12 == s2_pipeline_addr[9:4] ? regCount_18_1 : _GEN_89;
  wire [1:0] _GEN_91 = 6'h13 == s2_pipeline_addr[9:4] ? regCount_19_1 : _GEN_90;
  wire [1:0] _GEN_92 = 6'h14 == s2_pipeline_addr[9:4] ? regCount_20_1 : _GEN_91;
  wire [1:0] _GEN_93 = 6'h15 == s2_pipeline_addr[9:4] ? regCount_21_1 : _GEN_92;
  wire [1:0] _GEN_94 = 6'h16 == s2_pipeline_addr[9:4] ? regCount_22_1 : _GEN_93;
  wire [1:0] _GEN_95 = 6'h17 == s2_pipeline_addr[9:4] ? regCount_23_1 : _GEN_94;
  wire [1:0] _GEN_96 = 6'h18 == s2_pipeline_addr[9:4] ? regCount_24_1 : _GEN_95;
  wire [1:0] _GEN_97 = 6'h19 == s2_pipeline_addr[9:4] ? regCount_25_1 : _GEN_96;
  wire [1:0] _GEN_98 = 6'h1a == s2_pipeline_addr[9:4] ? regCount_26_1 : _GEN_97;
  wire [1:0] _GEN_99 = 6'h1b == s2_pipeline_addr[9:4] ? regCount_27_1 : _GEN_98;
  wire [1:0] _GEN_100 = 6'h1c == s2_pipeline_addr[9:4] ? regCount_28_1 : _GEN_99;
  wire [1:0] _GEN_101 = 6'h1d == s2_pipeline_addr[9:4] ? regCount_29_1 : _GEN_100;
  wire [1:0] _GEN_102 = 6'h1e == s2_pipeline_addr[9:4] ? regCount_30_1 : _GEN_101;
  wire [1:0] _GEN_103 = 6'h1f == s2_pipeline_addr[9:4] ? regCount_31_1 : _GEN_102;
  wire [1:0] _GEN_104 = 6'h20 == s2_pipeline_addr[9:4] ? regCount_32_1 : _GEN_103;
  wire [1:0] _GEN_105 = 6'h21 == s2_pipeline_addr[9:4] ? regCount_33_1 : _GEN_104;
  wire [1:0] _GEN_106 = 6'h22 == s2_pipeline_addr[9:4] ? regCount_34_1 : _GEN_105;
  wire [1:0] _GEN_107 = 6'h23 == s2_pipeline_addr[9:4] ? regCount_35_1 : _GEN_106;
  wire [1:0] _GEN_108 = 6'h24 == s2_pipeline_addr[9:4] ? regCount_36_1 : _GEN_107;
  wire [1:0] _GEN_109 = 6'h25 == s2_pipeline_addr[9:4] ? regCount_37_1 : _GEN_108;
  wire [1:0] _GEN_110 = 6'h26 == s2_pipeline_addr[9:4] ? regCount_38_1 : _GEN_109;
  wire [1:0] _GEN_111 = 6'h27 == s2_pipeline_addr[9:4] ? regCount_39_1 : _GEN_110;
  wire [1:0] _GEN_112 = 6'h28 == s2_pipeline_addr[9:4] ? regCount_40_1 : _GEN_111;
  wire [1:0] _GEN_113 = 6'h29 == s2_pipeline_addr[9:4] ? regCount_41_1 : _GEN_112;
  wire [1:0] _GEN_114 = 6'h2a == s2_pipeline_addr[9:4] ? regCount_42_1 : _GEN_113;
  wire [1:0] _GEN_115 = 6'h2b == s2_pipeline_addr[9:4] ? regCount_43_1 : _GEN_114;
  wire [1:0] _GEN_116 = 6'h2c == s2_pipeline_addr[9:4] ? regCount_44_1 : _GEN_115;
  wire [1:0] _GEN_117 = 6'h2d == s2_pipeline_addr[9:4] ? regCount_45_1 : _GEN_116;
  wire [1:0] _GEN_118 = 6'h2e == s2_pipeline_addr[9:4] ? regCount_46_1 : _GEN_117;
  wire [1:0] _GEN_119 = 6'h2f == s2_pipeline_addr[9:4] ? regCount_47_1 : _GEN_118;
  wire [1:0] _GEN_120 = 6'h30 == s2_pipeline_addr[9:4] ? regCount_48_1 : _GEN_119;
  wire [1:0] _GEN_121 = 6'h31 == s2_pipeline_addr[9:4] ? regCount_49_1 : _GEN_120;
  wire [1:0] _GEN_122 = 6'h32 == s2_pipeline_addr[9:4] ? regCount_50_1 : _GEN_121;
  wire [1:0] _GEN_123 = 6'h33 == s2_pipeline_addr[9:4] ? regCount_51_1 : _GEN_122;
  wire [1:0] _GEN_124 = 6'h34 == s2_pipeline_addr[9:4] ? regCount_52_1 : _GEN_123;
  wire [1:0] _GEN_125 = 6'h35 == s2_pipeline_addr[9:4] ? regCount_53_1 : _GEN_124;
  wire [1:0] _GEN_126 = 6'h36 == s2_pipeline_addr[9:4] ? regCount_54_1 : _GEN_125;
  wire [1:0] _GEN_127 = 6'h37 == s2_pipeline_addr[9:4] ? regCount_55_1 : _GEN_126;
  wire [1:0] _GEN_128 = 6'h38 == s2_pipeline_addr[9:4] ? regCount_56_1 : _GEN_127;
  wire [1:0] _GEN_129 = 6'h39 == s2_pipeline_addr[9:4] ? regCount_57_1 : _GEN_128;
  wire [1:0] _GEN_130 = 6'h3a == s2_pipeline_addr[9:4] ? regCount_58_1 : _GEN_129;
  wire [1:0] _GEN_131 = 6'h3b == s2_pipeline_addr[9:4] ? regCount_59_1 : _GEN_130;
  wire [1:0] _GEN_132 = 6'h3c == s2_pipeline_addr[9:4] ? regCount_60_1 : _GEN_131;
  wire [1:0] _GEN_133 = 6'h3d == s2_pipeline_addr[9:4] ? regCount_61_1 : _GEN_132;
  wire [1:0] _GEN_134 = 6'h3e == s2_pipeline_addr[9:4] ? regCount_62_1 : _GEN_133;
  wire [1:0] _GEN_135 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_1 : _GEN_134;
  wire [21:0] metaWays_2_tag = metaArray_2_io_r_data_tag;
  wire  metaWays_2_valid = metaArray_2_io_r_data_valid;
  wire  hitVec_2 = metaWays_2_valid & metaWays_2_tag == s2_pipeline_addr[31:10];
  wire [1:0] _GEN_137 = 6'h1 == s2_pipeline_addr[9:4] ? regCount_1_2 : regCount_0_2;
  wire [1:0] _GEN_138 = 6'h2 == s2_pipeline_addr[9:4] ? regCount_2_2 : _GEN_137;
  wire [1:0] _GEN_139 = 6'h3 == s2_pipeline_addr[9:4] ? regCount_3_2 : _GEN_138;
  wire [1:0] _GEN_140 = 6'h4 == s2_pipeline_addr[9:4] ? regCount_4_2 : _GEN_139;
  wire [1:0] _GEN_141 = 6'h5 == s2_pipeline_addr[9:4] ? regCount_5_2 : _GEN_140;
  wire [1:0] _GEN_142 = 6'h6 == s2_pipeline_addr[9:4] ? regCount_6_2 : _GEN_141;
  wire [1:0] _GEN_143 = 6'h7 == s2_pipeline_addr[9:4] ? regCount_7_2 : _GEN_142;
  wire [1:0] _GEN_144 = 6'h8 == s2_pipeline_addr[9:4] ? regCount_8_2 : _GEN_143;
  wire [1:0] _GEN_145 = 6'h9 == s2_pipeline_addr[9:4] ? regCount_9_2 : _GEN_144;
  wire [1:0] _GEN_146 = 6'ha == s2_pipeline_addr[9:4] ? regCount_10_2 : _GEN_145;
  wire [1:0] _GEN_147 = 6'hb == s2_pipeline_addr[9:4] ? regCount_11_2 : _GEN_146;
  wire [1:0] _GEN_148 = 6'hc == s2_pipeline_addr[9:4] ? regCount_12_2 : _GEN_147;
  wire [1:0] _GEN_149 = 6'hd == s2_pipeline_addr[9:4] ? regCount_13_2 : _GEN_148;
  wire [1:0] _GEN_150 = 6'he == s2_pipeline_addr[9:4] ? regCount_14_2 : _GEN_149;
  wire [1:0] _GEN_151 = 6'hf == s2_pipeline_addr[9:4] ? regCount_15_2 : _GEN_150;
  wire [1:0] _GEN_152 = 6'h10 == s2_pipeline_addr[9:4] ? regCount_16_2 : _GEN_151;
  wire [1:0] _GEN_153 = 6'h11 == s2_pipeline_addr[9:4] ? regCount_17_2 : _GEN_152;
  wire [1:0] _GEN_154 = 6'h12 == s2_pipeline_addr[9:4] ? regCount_18_2 : _GEN_153;
  wire [1:0] _GEN_155 = 6'h13 == s2_pipeline_addr[9:4] ? regCount_19_2 : _GEN_154;
  wire [1:0] _GEN_156 = 6'h14 == s2_pipeline_addr[9:4] ? regCount_20_2 : _GEN_155;
  wire [1:0] _GEN_157 = 6'h15 == s2_pipeline_addr[9:4] ? regCount_21_2 : _GEN_156;
  wire [1:0] _GEN_158 = 6'h16 == s2_pipeline_addr[9:4] ? regCount_22_2 : _GEN_157;
  wire [1:0] _GEN_159 = 6'h17 == s2_pipeline_addr[9:4] ? regCount_23_2 : _GEN_158;
  wire [1:0] _GEN_160 = 6'h18 == s2_pipeline_addr[9:4] ? regCount_24_2 : _GEN_159;
  wire [1:0] _GEN_161 = 6'h19 == s2_pipeline_addr[9:4] ? regCount_25_2 : _GEN_160;
  wire [1:0] _GEN_162 = 6'h1a == s2_pipeline_addr[9:4] ? regCount_26_2 : _GEN_161;
  wire [1:0] _GEN_163 = 6'h1b == s2_pipeline_addr[9:4] ? regCount_27_2 : _GEN_162;
  wire [1:0] _GEN_164 = 6'h1c == s2_pipeline_addr[9:4] ? regCount_28_2 : _GEN_163;
  wire [1:0] _GEN_165 = 6'h1d == s2_pipeline_addr[9:4] ? regCount_29_2 : _GEN_164;
  wire [1:0] _GEN_166 = 6'h1e == s2_pipeline_addr[9:4] ? regCount_30_2 : _GEN_165;
  wire [1:0] _GEN_167 = 6'h1f == s2_pipeline_addr[9:4] ? regCount_31_2 : _GEN_166;
  wire [1:0] _GEN_168 = 6'h20 == s2_pipeline_addr[9:4] ? regCount_32_2 : _GEN_167;
  wire [1:0] _GEN_169 = 6'h21 == s2_pipeline_addr[9:4] ? regCount_33_2 : _GEN_168;
  wire [1:0] _GEN_170 = 6'h22 == s2_pipeline_addr[9:4] ? regCount_34_2 : _GEN_169;
  wire [1:0] _GEN_171 = 6'h23 == s2_pipeline_addr[9:4] ? regCount_35_2 : _GEN_170;
  wire [1:0] _GEN_172 = 6'h24 == s2_pipeline_addr[9:4] ? regCount_36_2 : _GEN_171;
  wire [1:0] _GEN_173 = 6'h25 == s2_pipeline_addr[9:4] ? regCount_37_2 : _GEN_172;
  wire [1:0] _GEN_174 = 6'h26 == s2_pipeline_addr[9:4] ? regCount_38_2 : _GEN_173;
  wire [1:0] _GEN_175 = 6'h27 == s2_pipeline_addr[9:4] ? regCount_39_2 : _GEN_174;
  wire [1:0] _GEN_176 = 6'h28 == s2_pipeline_addr[9:4] ? regCount_40_2 : _GEN_175;
  wire [1:0] _GEN_177 = 6'h29 == s2_pipeline_addr[9:4] ? regCount_41_2 : _GEN_176;
  wire [1:0] _GEN_178 = 6'h2a == s2_pipeline_addr[9:4] ? regCount_42_2 : _GEN_177;
  wire [1:0] _GEN_179 = 6'h2b == s2_pipeline_addr[9:4] ? regCount_43_2 : _GEN_178;
  wire [1:0] _GEN_180 = 6'h2c == s2_pipeline_addr[9:4] ? regCount_44_2 : _GEN_179;
  wire [1:0] _GEN_181 = 6'h2d == s2_pipeline_addr[9:4] ? regCount_45_2 : _GEN_180;
  wire [1:0] _GEN_182 = 6'h2e == s2_pipeline_addr[9:4] ? regCount_46_2 : _GEN_181;
  wire [1:0] _GEN_183 = 6'h2f == s2_pipeline_addr[9:4] ? regCount_47_2 : _GEN_182;
  wire [1:0] _GEN_184 = 6'h30 == s2_pipeline_addr[9:4] ? regCount_48_2 : _GEN_183;
  wire [1:0] _GEN_185 = 6'h31 == s2_pipeline_addr[9:4] ? regCount_49_2 : _GEN_184;
  wire [1:0] _GEN_186 = 6'h32 == s2_pipeline_addr[9:4] ? regCount_50_2 : _GEN_185;
  wire [1:0] _GEN_187 = 6'h33 == s2_pipeline_addr[9:4] ? regCount_51_2 : _GEN_186;
  wire [1:0] _GEN_188 = 6'h34 == s2_pipeline_addr[9:4] ? regCount_52_2 : _GEN_187;
  wire [1:0] _GEN_189 = 6'h35 == s2_pipeline_addr[9:4] ? regCount_53_2 : _GEN_188;
  wire [1:0] _GEN_190 = 6'h36 == s2_pipeline_addr[9:4] ? regCount_54_2 : _GEN_189;
  wire [1:0] _GEN_191 = 6'h37 == s2_pipeline_addr[9:4] ? regCount_55_2 : _GEN_190;
  wire [1:0] _GEN_192 = 6'h38 == s2_pipeline_addr[9:4] ? regCount_56_2 : _GEN_191;
  wire [1:0] _GEN_193 = 6'h39 == s2_pipeline_addr[9:4] ? regCount_57_2 : _GEN_192;
  wire [1:0] _GEN_194 = 6'h3a == s2_pipeline_addr[9:4] ? regCount_58_2 : _GEN_193;
  wire [1:0] _GEN_195 = 6'h3b == s2_pipeline_addr[9:4] ? regCount_59_2 : _GEN_194;
  wire [1:0] _GEN_196 = 6'h3c == s2_pipeline_addr[9:4] ? regCount_60_2 : _GEN_195;
  wire [1:0] _GEN_197 = 6'h3d == s2_pipeline_addr[9:4] ? regCount_61_2 : _GEN_196;
  wire [1:0] _GEN_198 = 6'h3e == s2_pipeline_addr[9:4] ? regCount_62_2 : _GEN_197;
  wire [1:0] _GEN_199 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_2 : _GEN_198;
  wire [21:0] metaWays_3_tag = metaArray_3_io_r_data_tag;
  wire  metaWays_3_valid = metaArray_3_io_r_data_valid;
  wire  hitVec_3 = metaWays_3_valid & metaWays_3_tag == s2_pipeline_addr[31:10];
  wire [1:0] _GEN_201 = 6'h1 == s2_pipeline_addr[9:4] ? regCount_1_3 : regCount_0_3;
  wire [1:0] _GEN_202 = 6'h2 == s2_pipeline_addr[9:4] ? regCount_2_3 : _GEN_201;
  wire [1:0] _GEN_203 = 6'h3 == s2_pipeline_addr[9:4] ? regCount_3_3 : _GEN_202;
  wire [1:0] _GEN_204 = 6'h4 == s2_pipeline_addr[9:4] ? regCount_4_3 : _GEN_203;
  wire [1:0] _GEN_205 = 6'h5 == s2_pipeline_addr[9:4] ? regCount_5_3 : _GEN_204;
  wire [1:0] _GEN_206 = 6'h6 == s2_pipeline_addr[9:4] ? regCount_6_3 : _GEN_205;
  wire [1:0] _GEN_207 = 6'h7 == s2_pipeline_addr[9:4] ? regCount_7_3 : _GEN_206;
  wire [1:0] _GEN_208 = 6'h8 == s2_pipeline_addr[9:4] ? regCount_8_3 : _GEN_207;
  wire [1:0] _GEN_209 = 6'h9 == s2_pipeline_addr[9:4] ? regCount_9_3 : _GEN_208;
  wire [1:0] _GEN_210 = 6'ha == s2_pipeline_addr[9:4] ? regCount_10_3 : _GEN_209;
  wire [1:0] _GEN_211 = 6'hb == s2_pipeline_addr[9:4] ? regCount_11_3 : _GEN_210;
  wire [1:0] _GEN_212 = 6'hc == s2_pipeline_addr[9:4] ? regCount_12_3 : _GEN_211;
  wire [1:0] _GEN_213 = 6'hd == s2_pipeline_addr[9:4] ? regCount_13_3 : _GEN_212;
  wire [1:0] _GEN_214 = 6'he == s2_pipeline_addr[9:4] ? regCount_14_3 : _GEN_213;
  wire [1:0] _GEN_215 = 6'hf == s2_pipeline_addr[9:4] ? regCount_15_3 : _GEN_214;
  wire [1:0] _GEN_216 = 6'h10 == s2_pipeline_addr[9:4] ? regCount_16_3 : _GEN_215;
  wire [1:0] _GEN_217 = 6'h11 == s2_pipeline_addr[9:4] ? regCount_17_3 : _GEN_216;
  wire [1:0] _GEN_218 = 6'h12 == s2_pipeline_addr[9:4] ? regCount_18_3 : _GEN_217;
  wire [1:0] _GEN_219 = 6'h13 == s2_pipeline_addr[9:4] ? regCount_19_3 : _GEN_218;
  wire [1:0] _GEN_220 = 6'h14 == s2_pipeline_addr[9:4] ? regCount_20_3 : _GEN_219;
  wire [1:0] _GEN_221 = 6'h15 == s2_pipeline_addr[9:4] ? regCount_21_3 : _GEN_220;
  wire [1:0] _GEN_222 = 6'h16 == s2_pipeline_addr[9:4] ? regCount_22_3 : _GEN_221;
  wire [1:0] _GEN_223 = 6'h17 == s2_pipeline_addr[9:4] ? regCount_23_3 : _GEN_222;
  wire [1:0] _GEN_224 = 6'h18 == s2_pipeline_addr[9:4] ? regCount_24_3 : _GEN_223;
  wire [1:0] _GEN_225 = 6'h19 == s2_pipeline_addr[9:4] ? regCount_25_3 : _GEN_224;
  wire [1:0] _GEN_226 = 6'h1a == s2_pipeline_addr[9:4] ? regCount_26_3 : _GEN_225;
  wire [1:0] _GEN_227 = 6'h1b == s2_pipeline_addr[9:4] ? regCount_27_3 : _GEN_226;
  wire [1:0] _GEN_228 = 6'h1c == s2_pipeline_addr[9:4] ? regCount_28_3 : _GEN_227;
  wire [1:0] _GEN_229 = 6'h1d == s2_pipeline_addr[9:4] ? regCount_29_3 : _GEN_228;
  wire [1:0] _GEN_230 = 6'h1e == s2_pipeline_addr[9:4] ? regCount_30_3 : _GEN_229;
  wire [1:0] _GEN_231 = 6'h1f == s2_pipeline_addr[9:4] ? regCount_31_3 : _GEN_230;
  wire [1:0] _GEN_232 = 6'h20 == s2_pipeline_addr[9:4] ? regCount_32_3 : _GEN_231;
  wire [1:0] _GEN_233 = 6'h21 == s2_pipeline_addr[9:4] ? regCount_33_3 : _GEN_232;
  wire [1:0] _GEN_234 = 6'h22 == s2_pipeline_addr[9:4] ? regCount_34_3 : _GEN_233;
  wire [1:0] _GEN_235 = 6'h23 == s2_pipeline_addr[9:4] ? regCount_35_3 : _GEN_234;
  wire [1:0] _GEN_236 = 6'h24 == s2_pipeline_addr[9:4] ? regCount_36_3 : _GEN_235;
  wire [1:0] _GEN_237 = 6'h25 == s2_pipeline_addr[9:4] ? regCount_37_3 : _GEN_236;
  wire [1:0] _GEN_238 = 6'h26 == s2_pipeline_addr[9:4] ? regCount_38_3 : _GEN_237;
  wire [1:0] _GEN_239 = 6'h27 == s2_pipeline_addr[9:4] ? regCount_39_3 : _GEN_238;
  wire [1:0] _GEN_240 = 6'h28 == s2_pipeline_addr[9:4] ? regCount_40_3 : _GEN_239;
  wire [1:0] _GEN_241 = 6'h29 == s2_pipeline_addr[9:4] ? regCount_41_3 : _GEN_240;
  wire [1:0] _GEN_242 = 6'h2a == s2_pipeline_addr[9:4] ? regCount_42_3 : _GEN_241;
  wire [1:0] _GEN_243 = 6'h2b == s2_pipeline_addr[9:4] ? regCount_43_3 : _GEN_242;
  wire [1:0] _GEN_244 = 6'h2c == s2_pipeline_addr[9:4] ? regCount_44_3 : _GEN_243;
  wire [1:0] _GEN_245 = 6'h2d == s2_pipeline_addr[9:4] ? regCount_45_3 : _GEN_244;
  wire [1:0] _GEN_246 = 6'h2e == s2_pipeline_addr[9:4] ? regCount_46_3 : _GEN_245;
  wire [1:0] _GEN_247 = 6'h2f == s2_pipeline_addr[9:4] ? regCount_47_3 : _GEN_246;
  wire [1:0] _GEN_248 = 6'h30 == s2_pipeline_addr[9:4] ? regCount_48_3 : _GEN_247;
  wire [1:0] _GEN_249 = 6'h31 == s2_pipeline_addr[9:4] ? regCount_49_3 : _GEN_248;
  wire [1:0] _GEN_250 = 6'h32 == s2_pipeline_addr[9:4] ? regCount_50_3 : _GEN_249;
  wire [1:0] _GEN_251 = 6'h33 == s2_pipeline_addr[9:4] ? regCount_51_3 : _GEN_250;
  wire [1:0] _GEN_252 = 6'h34 == s2_pipeline_addr[9:4] ? regCount_52_3 : _GEN_251;
  wire [1:0] _GEN_253 = 6'h35 == s2_pipeline_addr[9:4] ? regCount_53_3 : _GEN_252;
  wire [1:0] _GEN_254 = 6'h36 == s2_pipeline_addr[9:4] ? regCount_54_3 : _GEN_253;
  wire [1:0] _GEN_255 = 6'h37 == s2_pipeline_addr[9:4] ? regCount_55_3 : _GEN_254;
  wire [1:0] _GEN_256 = 6'h38 == s2_pipeline_addr[9:4] ? regCount_56_3 : _GEN_255;
  wire [1:0] _GEN_257 = 6'h39 == s2_pipeline_addr[9:4] ? regCount_57_3 : _GEN_256;
  wire [1:0] _GEN_258 = 6'h3a == s2_pipeline_addr[9:4] ? regCount_58_3 : _GEN_257;
  wire [1:0] _GEN_259 = 6'h3b == s2_pipeline_addr[9:4] ? regCount_59_3 : _GEN_258;
  wire [1:0] _GEN_260 = 6'h3c == s2_pipeline_addr[9:4] ? regCount_60_3 : _GEN_259;
  wire [1:0] _GEN_261 = 6'h3d == s2_pipeline_addr[9:4] ? regCount_61_3 : _GEN_260;
  wire [1:0] _GEN_262 = 6'h3e == s2_pipeline_addr[9:4] ? regCount_62_3 : _GEN_261;
  wire [1:0] _GEN_263 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_3 : _GEN_262;
  wire [3:0] _s2_idxWayHit_T = {hitVec_3,hitVec_2,hitVec_1,hitVec_0};
  wire [1:0] s2_idxWayHit_hi_1 = _s2_idxWayHit_T[3:2];
  wire [1:0] s2_idxWayHit_lo_1 = _s2_idxWayHit_T[1:0];
  wire  _s2_idxWayHit_T_1 = |s2_idxWayHit_hi_1;
  wire [1:0] _s2_idxWayHit_T_2 = s2_idxWayHit_hi_1 | s2_idxWayHit_lo_1;
  wire [1:0] s2_idxWayHit = {_s2_idxWayHit_T_1,_s2_idxWayHit_T_2[1]};
  wire [1:0] s2_wordsMask = 2'h1 << s2_pipeline_addr[3];
  wire  s2_hit = s2_pipeline_valid & |_s2_idxWayHit_T;
  wire [63:0] _s2_dataBlockHit_T = hitVec_0 ? dataWays_0_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_1 = hitVec_1 ? dataWays_1_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_2 = hitVec_2 ? dataWays_2_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_3 = hitVec_3 ? dataWays_3_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_4 = _s2_dataBlockHit_T | _s2_dataBlockHit_T_1;
  wire [63:0] _s2_dataBlockHit_T_5 = _s2_dataBlockHit_T_4 | _s2_dataBlockHit_T_2;
  wire [63:0] s2_dataBlockHit_0 = _s2_dataBlockHit_T_5 | _s2_dataBlockHit_T_3;
  wire [63:0] _s2_dataBlockHit_T_7 = hitVec_0 ? dataWays_0_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_8 = hitVec_1 ? dataWays_1_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_9 = hitVec_2 ? dataWays_2_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_10 = hitVec_3 ? dataWays_3_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_11 = _s2_dataBlockHit_T_7 | _s2_dataBlockHit_T_8;
  wire [63:0] _s2_dataBlockHit_T_12 = _s2_dataBlockHit_T_11 | _s2_dataBlockHit_T_9;
  wire [63:0] s2_dataBlockHit_1 = _s2_dataBlockHit_T_12 | _s2_dataBlockHit_T_10;
  wire [63:0] _s2_hitWord_T_2 = s2_wordsMask[0] ? s2_dataBlockHit_0 : 64'h0;
  wire [63:0] _s2_hitWord_T_3 = s2_wordsMask[1] ? s2_dataBlockHit_1 : 64'h0;
  wire [63:0] s2_hitWord = _s2_hitWord_T_2 | _s2_hitWord_T_3;
  wire  s2_isMMIO = s2_pipeline_valid & s2_pipeline_isMMIO;
  wire  s2_miss = s2_pipeline_valid & ~s2_hit;
  wire  metaWays_0_needFlush = metaArray_0_io_r_data_needFlush;
  wire  metaWays_1_needFlush = metaArray_1_io_r_data_needFlush;
  wire  _GEN_265 = 2'h1 == selTree_io_outIdx ? metaWays_1_needFlush : metaWays_0_needFlush;
  wire  metaWays_2_needFlush = metaArray_2_io_r_data_needFlush;
  wire  _GEN_266 = 2'h2 == selTree_io_outIdx ? metaWays_2_needFlush : _GEN_265;
  wire  metaWays_3_needFlush = metaArray_3_io_r_data_needFlush;
  wire  _GEN_267 = 2'h3 == selTree_io_outIdx ? metaWays_3_needFlush : _GEN_266;
  wire [2:0] _GEN_268 = _GEN_267 ? 3'h3 : 3'h1;
  wire  _T_23 = io_out_req_ready & io_out_req_valid;
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid;
  wire [2:0] _GEN_272 = _T_25 ? 3'h7 : icache_status;
  wire [2:0] _GEN_273 = _T_23 ? 3'h4 : icache_status;
  wire [2:0] _GEN_274 = _T_25 ? 3'h1 : icache_status;
  wire  _T_31 = io_mmio_req_ready & io_mmio_req_valid;
  wire [2:0] _GEN_275 = _T_31 ? 3'h6 : icache_status;
  wire  _T_33 = io_mmio_resp_ready & io_mmio_resp_valid;
  wire [2:0] _GEN_276 = _T_33 ? 3'h7 : icache_status;
  wire [2:0] _GEN_277 = _s2_stall_T ? 3'h0 : icache_status;
  wire [2:0] _GEN_278 = 3'h7 == icache_status ? _GEN_277 : icache_status;
  wire [2:0] _GEN_279 = 3'h6 == icache_status ? _GEN_276 : _GEN_278;
  wire [2:0] _GEN_280 = 3'h5 == icache_status ? _GEN_275 : _GEN_279;
  wire [2:0] _GEN_281 = 3'h4 == icache_status ? _GEN_274 : _GEN_280;
  wire [2:0] _GEN_282 = 3'h3 == icache_status ? _GEN_273 : _GEN_281;
  wire  cacheUpdate = icache_status == 3'h2 & _T_25;
  wire  _hitUpdate_T = icache_status == 3'h0;
  wire  hitUpdate = icache_status == 3'h0 & s2_hit;
  wire  _metaArray_0_io_w_wen_T = 2'h0 == selTree_io_outIdx;
  wire  _metaArray_0_io_w_wen_T_1 = cacheUpdate & 2'h0 == selTree_io_outIdx;
  wire  _metaArray_1_io_w_wen_T = 2'h1 == selTree_io_outIdx;
  wire  _metaArray_1_io_w_wen_T_1 = cacheUpdate & 2'h1 == selTree_io_outIdx;
  wire  _metaArray_2_io_w_wen_T = 2'h2 == selTree_io_outIdx;
  wire  _metaArray_2_io_w_wen_T_1 = cacheUpdate & 2'h2 == selTree_io_outIdx;
  wire  _metaArray_3_io_w_wen_T = 2'h3 == selTree_io_outIdx;
  wire  _metaArray_3_io_w_wen_T_1 = cacheUpdate & 2'h3 == selTree_io_outIdx;
  wire [63:0] dataRefill_0 = io_out_resp_bits_rdata[63:0];
  wire [63:0] dataRefill_1 = io_out_resp_bits_rdata[127:64];
  wire [127:0] _io_dataArray_0_wdata_T_1 = {dataRefill_1,dataRefill_0};
  wire [1:0] _GEN_863 = 6'h0 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_0_1 : regCount_0_0;
  wire [1:0] _GEN_864 = 6'h0 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_0_2 : _GEN_863;
  wire [1:0] _GEN_865 = 6'h0 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_0_3 : _GEN_864;
  wire [1:0] _GEN_866 = 6'h1 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_1_0 : _GEN_865;
  wire [1:0] _GEN_867 = 6'h1 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_1_1 : _GEN_866;
  wire [1:0] _GEN_868 = 6'h1 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_1_2 : _GEN_867;
  wire [1:0] _GEN_869 = 6'h1 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_1_3 : _GEN_868;
  wire [1:0] _GEN_870 = 6'h2 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_2_0 : _GEN_869;
  wire [1:0] _GEN_871 = 6'h2 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_2_1 : _GEN_870;
  wire [1:0] _GEN_872 = 6'h2 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_2_2 : _GEN_871;
  wire [1:0] _GEN_873 = 6'h2 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_2_3 : _GEN_872;
  wire [1:0] _GEN_874 = 6'h3 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_3_0 : _GEN_873;
  wire [1:0] _GEN_875 = 6'h3 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_3_1 : _GEN_874;
  wire [1:0] _GEN_876 = 6'h3 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_3_2 : _GEN_875;
  wire [1:0] _GEN_877 = 6'h3 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_3_3 : _GEN_876;
  wire [1:0] _GEN_878 = 6'h4 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_4_0 : _GEN_877;
  wire [1:0] _GEN_879 = 6'h4 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_4_1 : _GEN_878;
  wire [1:0] _GEN_880 = 6'h4 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_4_2 : _GEN_879;
  wire [1:0] _GEN_881 = 6'h4 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_4_3 : _GEN_880;
  wire [1:0] _GEN_882 = 6'h5 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_5_0 : _GEN_881;
  wire [1:0] _GEN_883 = 6'h5 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_5_1 : _GEN_882;
  wire [1:0] _GEN_884 = 6'h5 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_5_2 : _GEN_883;
  wire [1:0] _GEN_885 = 6'h5 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_5_3 : _GEN_884;
  wire [1:0] _GEN_886 = 6'h6 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_6_0 : _GEN_885;
  wire [1:0] _GEN_887 = 6'h6 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_6_1 : _GEN_886;
  wire [1:0] _GEN_888 = 6'h6 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_6_2 : _GEN_887;
  wire [1:0] _GEN_889 = 6'h6 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_6_3 : _GEN_888;
  wire [1:0] _GEN_890 = 6'h7 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_7_0 : _GEN_889;
  wire [1:0] _GEN_891 = 6'h7 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_7_1 : _GEN_890;
  wire [1:0] _GEN_892 = 6'h7 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_7_2 : _GEN_891;
  wire [1:0] _GEN_893 = 6'h7 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_7_3 : _GEN_892;
  wire [1:0] _GEN_894 = 6'h8 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_8_0 : _GEN_893;
  wire [1:0] _GEN_895 = 6'h8 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_8_1 : _GEN_894;
  wire [1:0] _GEN_896 = 6'h8 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_8_2 : _GEN_895;
  wire [1:0] _GEN_897 = 6'h8 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_8_3 : _GEN_896;
  wire [1:0] _GEN_898 = 6'h9 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_9_0 : _GEN_897;
  wire [1:0] _GEN_899 = 6'h9 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_9_1 : _GEN_898;
  wire [1:0] _GEN_900 = 6'h9 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_9_2 : _GEN_899;
  wire [1:0] _GEN_901 = 6'h9 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_9_3 : _GEN_900;
  wire [1:0] _GEN_902 = 6'ha == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_10_0 : _GEN_901;
  wire [1:0] _GEN_903 = 6'ha == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_10_1 : _GEN_902;
  wire [1:0] _GEN_904 = 6'ha == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_10_2 : _GEN_903;
  wire [1:0] _GEN_905 = 6'ha == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_10_3 : _GEN_904;
  wire [1:0] _GEN_906 = 6'hb == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_11_0 : _GEN_905;
  wire [1:0] _GEN_907 = 6'hb == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_11_1 : _GEN_906;
  wire [1:0] _GEN_908 = 6'hb == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_11_2 : _GEN_907;
  wire [1:0] _GEN_909 = 6'hb == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_11_3 : _GEN_908;
  wire [1:0] _GEN_910 = 6'hc == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_12_0 : _GEN_909;
  wire [1:0] _GEN_911 = 6'hc == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_12_1 : _GEN_910;
  wire [1:0] _GEN_912 = 6'hc == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_12_2 : _GEN_911;
  wire [1:0] _GEN_913 = 6'hc == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_12_3 : _GEN_912;
  wire [1:0] _GEN_914 = 6'hd == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_13_0 : _GEN_913;
  wire [1:0] _GEN_915 = 6'hd == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_13_1 : _GEN_914;
  wire [1:0] _GEN_916 = 6'hd == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_13_2 : _GEN_915;
  wire [1:0] _GEN_917 = 6'hd == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_13_3 : _GEN_916;
  wire [1:0] _GEN_918 = 6'he == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_14_0 : _GEN_917;
  wire [1:0] _GEN_919 = 6'he == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_14_1 : _GEN_918;
  wire [1:0] _GEN_920 = 6'he == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_14_2 : _GEN_919;
  wire [1:0] _GEN_921 = 6'he == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_14_3 : _GEN_920;
  wire [1:0] _GEN_922 = 6'hf == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_15_0 : _GEN_921;
  wire [1:0] _GEN_923 = 6'hf == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_15_1 : _GEN_922;
  wire [1:0] _GEN_924 = 6'hf == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_15_2 : _GEN_923;
  wire [1:0] _GEN_925 = 6'hf == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_15_3 : _GEN_924;
  wire [1:0] _GEN_926 = 6'h10 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_16_0 : _GEN_925;
  wire [1:0] _GEN_927 = 6'h10 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_16_1 : _GEN_926;
  wire [1:0] _GEN_928 = 6'h10 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_16_2 : _GEN_927;
  wire [1:0] _GEN_929 = 6'h10 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_16_3 : _GEN_928;
  wire [1:0] _GEN_930 = 6'h11 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_17_0 : _GEN_929;
  wire [1:0] _GEN_931 = 6'h11 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_17_1 : _GEN_930;
  wire [1:0] _GEN_932 = 6'h11 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_17_2 : _GEN_931;
  wire [1:0] _GEN_933 = 6'h11 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_17_3 : _GEN_932;
  wire [1:0] _GEN_934 = 6'h12 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_18_0 : _GEN_933;
  wire [1:0] _GEN_935 = 6'h12 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_18_1 : _GEN_934;
  wire [1:0] _GEN_936 = 6'h12 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_18_2 : _GEN_935;
  wire [1:0] _GEN_937 = 6'h12 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_18_3 : _GEN_936;
  wire [1:0] _GEN_938 = 6'h13 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_19_0 : _GEN_937;
  wire [1:0] _GEN_939 = 6'h13 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_19_1 : _GEN_938;
  wire [1:0] _GEN_940 = 6'h13 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_19_2 : _GEN_939;
  wire [1:0] _GEN_941 = 6'h13 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_19_3 : _GEN_940;
  wire [1:0] _GEN_942 = 6'h14 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_20_0 : _GEN_941;
  wire [1:0] _GEN_943 = 6'h14 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_20_1 : _GEN_942;
  wire [1:0] _GEN_944 = 6'h14 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_20_2 : _GEN_943;
  wire [1:0] _GEN_945 = 6'h14 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_20_3 : _GEN_944;
  wire [1:0] _GEN_946 = 6'h15 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_21_0 : _GEN_945;
  wire [1:0] _GEN_947 = 6'h15 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_21_1 : _GEN_946;
  wire [1:0] _GEN_948 = 6'h15 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_21_2 : _GEN_947;
  wire [1:0] _GEN_949 = 6'h15 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_21_3 : _GEN_948;
  wire [1:0] _GEN_950 = 6'h16 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_22_0 : _GEN_949;
  wire [1:0] _GEN_951 = 6'h16 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_22_1 : _GEN_950;
  wire [1:0] _GEN_952 = 6'h16 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_22_2 : _GEN_951;
  wire [1:0] _GEN_953 = 6'h16 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_22_3 : _GEN_952;
  wire [1:0] _GEN_954 = 6'h17 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_23_0 : _GEN_953;
  wire [1:0] _GEN_955 = 6'h17 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_23_1 : _GEN_954;
  wire [1:0] _GEN_956 = 6'h17 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_23_2 : _GEN_955;
  wire [1:0] _GEN_957 = 6'h17 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_23_3 : _GEN_956;
  wire [1:0] _GEN_958 = 6'h18 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_24_0 : _GEN_957;
  wire [1:0] _GEN_959 = 6'h18 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_24_1 : _GEN_958;
  wire [1:0] _GEN_960 = 6'h18 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_24_2 : _GEN_959;
  wire [1:0] _GEN_961 = 6'h18 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_24_3 : _GEN_960;
  wire [1:0] _GEN_962 = 6'h19 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_25_0 : _GEN_961;
  wire [1:0] _GEN_963 = 6'h19 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_25_1 : _GEN_962;
  wire [1:0] _GEN_964 = 6'h19 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_25_2 : _GEN_963;
  wire [1:0] _GEN_965 = 6'h19 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_25_3 : _GEN_964;
  wire [1:0] _GEN_966 = 6'h1a == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_26_0 : _GEN_965;
  wire [1:0] _GEN_967 = 6'h1a == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_26_1 : _GEN_966;
  wire [1:0] _GEN_968 = 6'h1a == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_26_2 : _GEN_967;
  wire [1:0] _GEN_969 = 6'h1a == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_26_3 : _GEN_968;
  wire [1:0] _GEN_970 = 6'h1b == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_27_0 : _GEN_969;
  wire [1:0] _GEN_971 = 6'h1b == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_27_1 : _GEN_970;
  wire [1:0] _GEN_972 = 6'h1b == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_27_2 : _GEN_971;
  wire [1:0] _GEN_973 = 6'h1b == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_27_3 : _GEN_972;
  wire [1:0] _GEN_974 = 6'h1c == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_28_0 : _GEN_973;
  wire [1:0] _GEN_975 = 6'h1c == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_28_1 : _GEN_974;
  wire [1:0] _GEN_976 = 6'h1c == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_28_2 : _GEN_975;
  wire [1:0] _GEN_977 = 6'h1c == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_28_3 : _GEN_976;
  wire [1:0] _GEN_978 = 6'h1d == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_29_0 : _GEN_977;
  wire [1:0] _GEN_979 = 6'h1d == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_29_1 : _GEN_978;
  wire [1:0] _GEN_980 = 6'h1d == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_29_2 : _GEN_979;
  wire [1:0] _GEN_981 = 6'h1d == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_29_3 : _GEN_980;
  wire [1:0] _GEN_982 = 6'h1e == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_30_0 : _GEN_981;
  wire [1:0] _GEN_983 = 6'h1e == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_30_1 : _GEN_982;
  wire [1:0] _GEN_984 = 6'h1e == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_30_2 : _GEN_983;
  wire [1:0] _GEN_985 = 6'h1e == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_30_3 : _GEN_984;
  wire [1:0] _GEN_986 = 6'h1f == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_31_0 : _GEN_985;
  wire [1:0] _GEN_987 = 6'h1f == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_31_1 : _GEN_986;
  wire [1:0] _GEN_988 = 6'h1f == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_31_2 : _GEN_987;
  wire [1:0] _GEN_989 = 6'h1f == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_31_3 : _GEN_988;
  wire [1:0] _GEN_990 = 6'h20 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_32_0 : _GEN_989;
  wire [1:0] _GEN_991 = 6'h20 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_32_1 : _GEN_990;
  wire [1:0] _GEN_992 = 6'h20 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_32_2 : _GEN_991;
  wire [1:0] _GEN_993 = 6'h20 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_32_3 : _GEN_992;
  wire [1:0] _GEN_994 = 6'h21 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_33_0 : _GEN_993;
  wire [1:0] _GEN_995 = 6'h21 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_33_1 : _GEN_994;
  wire [1:0] _GEN_996 = 6'h21 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_33_2 : _GEN_995;
  wire [1:0] _GEN_997 = 6'h21 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_33_3 : _GEN_996;
  wire [1:0] _GEN_998 = 6'h22 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_34_0 : _GEN_997;
  wire [1:0] _GEN_999 = 6'h22 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_34_1 : _GEN_998;
  wire [1:0] _GEN_1000 = 6'h22 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_34_2 : _GEN_999;
  wire [1:0] _GEN_1001 = 6'h22 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_34_3 : _GEN_1000;
  wire [1:0] _GEN_1002 = 6'h23 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_35_0 : _GEN_1001;
  wire [1:0] _GEN_1003 = 6'h23 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_35_1 : _GEN_1002;
  wire [1:0] _GEN_1004 = 6'h23 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_35_2 : _GEN_1003;
  wire [1:0] _GEN_1005 = 6'h23 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_35_3 : _GEN_1004;
  wire [1:0] _GEN_1006 = 6'h24 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_36_0 : _GEN_1005;
  wire [1:0] _GEN_1007 = 6'h24 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_36_1 : _GEN_1006;
  wire [1:0] _GEN_1008 = 6'h24 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_36_2 : _GEN_1007;
  wire [1:0] _GEN_1009 = 6'h24 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_36_3 : _GEN_1008;
  wire [1:0] _GEN_1010 = 6'h25 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_37_0 : _GEN_1009;
  wire [1:0] _GEN_1011 = 6'h25 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_37_1 : _GEN_1010;
  wire [1:0] _GEN_1012 = 6'h25 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_37_2 : _GEN_1011;
  wire [1:0] _GEN_1013 = 6'h25 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_37_3 : _GEN_1012;
  wire [1:0] _GEN_1014 = 6'h26 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_38_0 : _GEN_1013;
  wire [1:0] _GEN_1015 = 6'h26 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_38_1 : _GEN_1014;
  wire [1:0] _GEN_1016 = 6'h26 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_38_2 : _GEN_1015;
  wire [1:0] _GEN_1017 = 6'h26 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_38_3 : _GEN_1016;
  wire [1:0] _GEN_1018 = 6'h27 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_39_0 : _GEN_1017;
  wire [1:0] _GEN_1019 = 6'h27 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_39_1 : _GEN_1018;
  wire [1:0] _GEN_1020 = 6'h27 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_39_2 : _GEN_1019;
  wire [1:0] _GEN_1021 = 6'h27 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_39_3 : _GEN_1020;
  wire [1:0] _GEN_1022 = 6'h28 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_40_0 : _GEN_1021;
  wire [1:0] _GEN_1023 = 6'h28 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_40_1 : _GEN_1022;
  wire [1:0] _GEN_1024 = 6'h28 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_40_2 : _GEN_1023;
  wire [1:0] _GEN_1025 = 6'h28 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_40_3 : _GEN_1024;
  wire [1:0] _GEN_1026 = 6'h29 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_41_0 : _GEN_1025;
  wire [1:0] _GEN_1027 = 6'h29 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_41_1 : _GEN_1026;
  wire [1:0] _GEN_1028 = 6'h29 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_41_2 : _GEN_1027;
  wire [1:0] _GEN_1029 = 6'h29 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_41_3 : _GEN_1028;
  wire [1:0] _GEN_1030 = 6'h2a == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_42_0 : _GEN_1029;
  wire [1:0] _GEN_1031 = 6'h2a == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_42_1 : _GEN_1030;
  wire [1:0] _GEN_1032 = 6'h2a == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_42_2 : _GEN_1031;
  wire [1:0] _GEN_1033 = 6'h2a == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_42_3 : _GEN_1032;
  wire [1:0] _GEN_1034 = 6'h2b == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_43_0 : _GEN_1033;
  wire [1:0] _GEN_1035 = 6'h2b == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_43_1 : _GEN_1034;
  wire [1:0] _GEN_1036 = 6'h2b == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_43_2 : _GEN_1035;
  wire [1:0] _GEN_1037 = 6'h2b == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_43_3 : _GEN_1036;
  wire [1:0] _GEN_1038 = 6'h2c == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_44_0 : _GEN_1037;
  wire [1:0] _GEN_1039 = 6'h2c == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_44_1 : _GEN_1038;
  wire [1:0] _GEN_1040 = 6'h2c == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_44_2 : _GEN_1039;
  wire [1:0] _GEN_1041 = 6'h2c == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_44_3 : _GEN_1040;
  wire [1:0] _GEN_1042 = 6'h2d == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_45_0 : _GEN_1041;
  wire [1:0] _GEN_1043 = 6'h2d == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_45_1 : _GEN_1042;
  wire [1:0] _GEN_1044 = 6'h2d == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_45_2 : _GEN_1043;
  wire [1:0] _GEN_1045 = 6'h2d == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_45_3 : _GEN_1044;
  wire [1:0] _GEN_1046 = 6'h2e == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_46_0 : _GEN_1045;
  wire [1:0] _GEN_1047 = 6'h2e == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_46_1 : _GEN_1046;
  wire [1:0] _GEN_1048 = 6'h2e == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_46_2 : _GEN_1047;
  wire [1:0] _GEN_1049 = 6'h2e == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_46_3 : _GEN_1048;
  wire [1:0] _GEN_1050 = 6'h2f == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_47_0 : _GEN_1049;
  wire [1:0] _GEN_1051 = 6'h2f == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_47_1 : _GEN_1050;
  wire [1:0] _GEN_1052 = 6'h2f == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_47_2 : _GEN_1051;
  wire [1:0] _GEN_1053 = 6'h2f == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_47_3 : _GEN_1052;
  wire [1:0] _GEN_1054 = 6'h30 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_48_0 : _GEN_1053;
  wire [1:0] _GEN_1055 = 6'h30 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_48_1 : _GEN_1054;
  wire [1:0] _GEN_1056 = 6'h30 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_48_2 : _GEN_1055;
  wire [1:0] _GEN_1057 = 6'h30 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_48_3 : _GEN_1056;
  wire [1:0] _GEN_1058 = 6'h31 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_49_0 : _GEN_1057;
  wire [1:0] _GEN_1059 = 6'h31 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_49_1 : _GEN_1058;
  wire [1:0] _GEN_1060 = 6'h31 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_49_2 : _GEN_1059;
  wire [1:0] _GEN_1061 = 6'h31 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_49_3 : _GEN_1060;
  wire [1:0] _GEN_1062 = 6'h32 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_50_0 : _GEN_1061;
  wire [1:0] _GEN_1063 = 6'h32 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_50_1 : _GEN_1062;
  wire [1:0] _GEN_1064 = 6'h32 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_50_2 : _GEN_1063;
  wire [1:0] _GEN_1065 = 6'h32 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_50_3 : _GEN_1064;
  wire [1:0] _GEN_1066 = 6'h33 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_51_0 : _GEN_1065;
  wire [1:0] _GEN_1067 = 6'h33 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_51_1 : _GEN_1066;
  wire [1:0] _GEN_1068 = 6'h33 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_51_2 : _GEN_1067;
  wire [1:0] _GEN_1069 = 6'h33 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_51_3 : _GEN_1068;
  wire [1:0] _GEN_1070 = 6'h34 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_52_0 : _GEN_1069;
  wire [1:0] _GEN_1071 = 6'h34 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_52_1 : _GEN_1070;
  wire [1:0] _GEN_1072 = 6'h34 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_52_2 : _GEN_1071;
  wire [1:0] _GEN_1073 = 6'h34 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_52_3 : _GEN_1072;
  wire [1:0] _GEN_1074 = 6'h35 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_53_0 : _GEN_1073;
  wire [1:0] _GEN_1075 = 6'h35 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_53_1 : _GEN_1074;
  wire [1:0] _GEN_1076 = 6'h35 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_53_2 : _GEN_1075;
  wire [1:0] _GEN_1077 = 6'h35 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_53_3 : _GEN_1076;
  wire [1:0] _GEN_1078 = 6'h36 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_54_0 : _GEN_1077;
  wire [1:0] _GEN_1079 = 6'h36 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_54_1 : _GEN_1078;
  wire [1:0] _GEN_1080 = 6'h36 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_54_2 : _GEN_1079;
  wire [1:0] _GEN_1081 = 6'h36 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_54_3 : _GEN_1080;
  wire [1:0] _GEN_1082 = 6'h37 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_55_0 : _GEN_1081;
  wire [1:0] _GEN_1083 = 6'h37 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_55_1 : _GEN_1082;
  wire [1:0] _GEN_1084 = 6'h37 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_55_2 : _GEN_1083;
  wire [1:0] _GEN_1085 = 6'h37 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_55_3 : _GEN_1084;
  wire [1:0] _GEN_1086 = 6'h38 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_56_0 : _GEN_1085;
  wire [1:0] _GEN_1087 = 6'h38 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_56_1 : _GEN_1086;
  wire [1:0] _GEN_1088 = 6'h38 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_56_2 : _GEN_1087;
  wire [1:0] _GEN_1089 = 6'h38 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_56_3 : _GEN_1088;
  wire [1:0] _GEN_1090 = 6'h39 == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_57_0 : _GEN_1089;
  wire [1:0] _GEN_1091 = 6'h39 == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_57_1 : _GEN_1090;
  wire [1:0] _GEN_1092 = 6'h39 == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_57_2 : _GEN_1091;
  wire [1:0] _GEN_1093 = 6'h39 == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_57_3 : _GEN_1092;
  wire [1:0] _GEN_1094 = 6'h3a == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_58_0 : _GEN_1093;
  wire [1:0] _GEN_1095 = 6'h3a == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_58_1 : _GEN_1094;
  wire [1:0] _GEN_1096 = 6'h3a == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_58_2 : _GEN_1095;
  wire [1:0] _GEN_1097 = 6'h3a == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_58_3 : _GEN_1096;
  wire [1:0] _GEN_1098 = 6'h3b == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_59_0 : _GEN_1097;
  wire [1:0] _GEN_1099 = 6'h3b == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_59_1 : _GEN_1098;
  wire [1:0] _GEN_1100 = 6'h3b == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_59_2 : _GEN_1099;
  wire [1:0] _GEN_1101 = 6'h3b == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_59_3 : _GEN_1100;
  wire [1:0] _GEN_1102 = 6'h3c == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_60_0 : _GEN_1101;
  wire [1:0] _GEN_1103 = 6'h3c == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_60_1 : _GEN_1102;
  wire [1:0] _GEN_1104 = 6'h3c == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_60_2 : _GEN_1103;
  wire [1:0] _GEN_1105 = 6'h3c == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_60_3 : _GEN_1104;
  wire [1:0] _GEN_1106 = 6'h3d == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_61_0 : _GEN_1105;
  wire [1:0] _GEN_1107 = 6'h3d == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_61_1 : _GEN_1106;
  wire [1:0] _GEN_1108 = 6'h3d == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_61_2 : _GEN_1107;
  wire [1:0] _GEN_1109 = 6'h3d == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_61_3 : _GEN_1108;
  wire [1:0] _GEN_1110 = 6'h3e == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_62_0 : _GEN_1109;
  wire [1:0] _GEN_1111 = 6'h3e == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_62_1 : _GEN_1110;
  wire [1:0] _GEN_1112 = 6'h3e == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_62_2 : _GEN_1111;
  wire [1:0] _GEN_1113 = 6'h3e == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_62_3 : _GEN_1112;
  wire [1:0] _GEN_1114 = 6'h3f == s2_pipeline_addr[9:4] & 2'h0 == s2_idxWayHit ? regCount_63_0 : _GEN_1113;
  wire [1:0] _GEN_1115 = 6'h3f == s2_pipeline_addr[9:4] & 2'h1 == s2_idxWayHit ? regCount_63_1 : _GEN_1114;
  wire [1:0] _GEN_1116 = 6'h3f == s2_pipeline_addr[9:4] & 2'h2 == s2_idxWayHit ? regCount_63_2 : _GEN_1115;
  wire [1:0] _GEN_1117 = 6'h3f == s2_pipeline_addr[9:4] & 2'h3 == s2_idxWayHit ? regCount_63_3 : _GEN_1116;
  wire [1:0] _newCountHit_0_T_5 = _GEN_71 + 2'h1;
  wire [1:0] _GEN_1246 = _GEN_71 < _GEN_1117 ? _newCountHit_0_T_5 : _GEN_71;
  wire [1:0] newCountHit_0 = 2'h0 != s2_idxWayHit ? _GEN_1246 : 2'h0;
  wire [1:0] _newCountHit_1_T_5 = _GEN_135 + 2'h1;
  wire [1:0] _GEN_1696 = _GEN_135 < _GEN_1117 ? _newCountHit_1_T_5 : _GEN_135;
  wire [1:0] newCountHit_1 = 2'h1 != s2_idxWayHit ? _GEN_1696 : 2'h0;
  wire [1:0] _newCountHit_2_T_5 = _GEN_199 + 2'h1;
  wire [1:0] _GEN_2146 = _GEN_199 < _GEN_1117 ? _newCountHit_2_T_5 : _GEN_199;
  wire [1:0] newCountHit_2 = 2'h2 != s2_idxWayHit ? _GEN_2146 : 2'h0;
  wire [1:0] _newCountHit_3_T_5 = _GEN_263 + 2'h1;
  wire [1:0] _GEN_2596 = _GEN_263 < _GEN_1117 ? _newCountHit_3_T_5 : _GEN_263;
  wire [1:0] newCountHit_3 = 2'h3 != s2_idxWayHit ? _GEN_2596 : 2'h0;
  wire [1:0] _GEN_2726 = metaWays_0_valid ? _newCountHit_0_T_5 : _GEN_71;
  wire [1:0] newCountRefill_0 = _metaArray_0_io_w_wen_T ? 2'h0 : _GEN_2726;
  wire [1:0] _GEN_2856 = metaWays_1_valid ? _newCountHit_1_T_5 : _GEN_135;
  wire [1:0] newCountRefill_1 = _metaArray_1_io_w_wen_T ? 2'h0 : _GEN_2856;
  wire [1:0] _GEN_2986 = metaWays_2_valid ? _newCountHit_2_T_5 : _GEN_199;
  wire [1:0] newCountRefill_2 = _metaArray_2_io_w_wen_T ? 2'h0 : _GEN_2986;
  wire [1:0] _GEN_3116 = metaWays_3_valid ? _newCountHit_3_T_5 : _GEN_263;
  wire [1:0] newCountRefill_3 = _metaArray_3_io_w_wen_T ? 2'h0 : _GEN_3116;
  wire  countUpdate = hitUpdate | cacheUpdate;
  reg [63:0] mmioRespData;
  wire [63:0] rdata = s2_pipeline_isMMIO ? mmioRespData : s2_hitWord;
  wire  _mmioResp_T = icache_status == 3'h7;
  wire  mmioResp = icache_status == 3'h7 & s2_pipeline_isMMIO;
  wire  _cacheResp_T_2 = _hitUpdate_T | _mmioResp_T;
  wire  cacheResp = (_hitUpdate_T | _mmioResp_T) & s2_hit & ~s2_pipeline_isMMIO;
  wire [21:0] _GEN_3632 = 2'h1 == selTree_io_outIdx ? metaWays_1_tag : metaWays_0_tag;
  wire [21:0] _GEN_3633 = 2'h2 == selTree_io_outIdx ? metaWays_2_tag : _GEN_3632;
  wire [21:0] _GEN_3634 = 2'h3 == selTree_io_outIdx ? metaWays_3_tag : _GEN_3633;
  wire [31:0] writeBackAddr = {_GEN_3634,s2_pipeline_addr[9:4],4'h0};
  wire  _x5_T = icache_status == 3'h3;
  wire [63:0] _GEN_3636 = 2'h1 == selTree_io_outIdx ? dataWays_1_1 : dataWays_0_1;
  wire [63:0] _GEN_3637 = 2'h2 == selTree_io_outIdx ? dataWays_2_1 : _GEN_3636;
  wire [63:0] _GEN_3638 = 2'h3 == selTree_io_outIdx ? dataWays_3_1 : _GEN_3637;
  wire [63:0] _GEN_3640 = 2'h1 == selTree_io_outIdx ? dataWays_1_0 : dataWays_0_0;
  wire [63:0] _GEN_3641 = 2'h2 == selTree_io_outIdx ? dataWays_2_0 : _GEN_3640;
  wire [63:0] _GEN_3642 = 2'h3 == selTree_io_outIdx ? dataWays_3_0 : _GEN_3641;
  wire [127:0] _x6_T_1 = {_GEN_3638,_GEN_3642};
  ysyx_040656_SRAM metaArray_0 (
    .clock(metaArray_0_clock),
    .reset(metaArray_0_reset),
    .io_w_setIdx(metaArray_0_io_w_setIdx),
    .io_w_data_tag(metaArray_0_io_w_data_tag),
    .io_w_data_valid(metaArray_0_io_w_data_valid),
    .io_w_data_needFlush(metaArray_0_io_w_data_needFlush),
    .io_w_wen(metaArray_0_io_w_wen),
    .io_r_setIdx(metaArray_0_io_r_setIdx),
    .io_r_data_tag(metaArray_0_io_r_data_tag),
    .io_r_data_valid(metaArray_0_io_r_data_valid),
    .io_r_data_needFlush(metaArray_0_io_r_data_needFlush),
    .io_r_ren(metaArray_0_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_1 (
    .clock(metaArray_1_clock),
    .reset(metaArray_1_reset),
    .io_w_setIdx(metaArray_1_io_w_setIdx),
    .io_w_data_tag(metaArray_1_io_w_data_tag),
    .io_w_data_valid(metaArray_1_io_w_data_valid),
    .io_w_data_needFlush(metaArray_1_io_w_data_needFlush),
    .io_w_wen(metaArray_1_io_w_wen),
    .io_r_setIdx(metaArray_1_io_r_setIdx),
    .io_r_data_tag(metaArray_1_io_r_data_tag),
    .io_r_data_valid(metaArray_1_io_r_data_valid),
    .io_r_data_needFlush(metaArray_1_io_r_data_needFlush),
    .io_r_ren(metaArray_1_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_2 (
    .clock(metaArray_2_clock),
    .reset(metaArray_2_reset),
    .io_w_setIdx(metaArray_2_io_w_setIdx),
    .io_w_data_tag(metaArray_2_io_w_data_tag),
    .io_w_data_valid(metaArray_2_io_w_data_valid),
    .io_w_data_needFlush(metaArray_2_io_w_data_needFlush),
    .io_w_wen(metaArray_2_io_w_wen),
    .io_r_setIdx(metaArray_2_io_r_setIdx),
    .io_r_data_tag(metaArray_2_io_r_data_tag),
    .io_r_data_valid(metaArray_2_io_r_data_valid),
    .io_r_data_needFlush(metaArray_2_io_r_data_needFlush),
    .io_r_ren(metaArray_2_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_3 (
    .clock(metaArray_3_clock),
    .reset(metaArray_3_reset),
    .io_w_setIdx(metaArray_3_io_w_setIdx),
    .io_w_data_tag(metaArray_3_io_w_data_tag),
    .io_w_data_valid(metaArray_3_io_w_data_valid),
    .io_w_data_needFlush(metaArray_3_io_w_data_needFlush),
    .io_w_wen(metaArray_3_io_w_wen),
    .io_r_setIdx(metaArray_3_io_r_setIdx),
    .io_r_data_tag(metaArray_3_io_r_data_tag),
    .io_r_data_valid(metaArray_3_io_r_data_valid),
    .io_r_data_needFlush(metaArray_3_io_r_data_needFlush),
    .io_r_ren(metaArray_3_io_r_ren)
  );
  ysyx_040656_LRU selTree (
    .io_inWayValid_0(selTree_io_inWayValid_0),
    .io_inWayValid_1(selTree_io_inWayValid_1),
    .io_inWayValid_2(selTree_io_inWayValid_2),
    .io_inWayValid_3(selTree_io_inWayValid_3),
    .io_inValue_0(selTree_io_inValue_0),
    .io_inValue_1(selTree_io_inValue_1),
    .io_inValue_2(selTree_io_inValue_2),
    .io_inValue_3(selTree_io_inValue_3),
    .io_outIdx(selTree_io_outIdx)
  );
  assign io_in_req_ready = _cacheResp_T_2 & _T_15;
  assign io_in_resp_valid = mmioResp | cacheResp;
  assign io_in_resp_bits_rdata = s2_pipeline_addr[2:0] == 3'h4 ? rdata[63:32] : rdata[31:0];
  assign io_out_req_valid = icache_status == 3'h1 | _x5_T;
  assign io_out_req_bits_addr = icache_status == 3'h3 ? writeBackAddr : s2_pipeline_addr;
  assign io_out_req_bits_wdata = icache_status == 3'h3 ? _x6_T_1 : 128'h0;
  assign io_out_req_bits_cmd = {{2'd0}, _x5_T};
  assign io_out_resp_ready = 1'h1;
  assign io_mmio_req_valid = icache_status == 3'h5;
  assign io_mmio_req_bits_addr = s2_pipeline_addr;
  assign io_mmio_req_bits_size = s2_pipeline_size;
  assign io_mmio_resp_ready = 1'h1;
  assign io_dataArray_0_wen = ~(reset | _metaArray_0_io_w_wen_T_1);
  assign io_dataArray_0_addr = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign io_dataArray_0_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_1_wen = ~(reset | _metaArray_1_io_w_wen_T_1);
  assign io_dataArray_1_addr = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign io_dataArray_1_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_2_wen = ~(reset | _metaArray_2_io_w_wen_T_1);
  assign io_dataArray_2_addr = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign io_dataArray_2_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_3_wen = ~(reset | _metaArray_3_io_w_wen_T_1);
  assign io_dataArray_3_addr = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign io_dataArray_3_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign metaArray_0_clock = clock;
  assign metaArray_0_reset = reset | difftestFENCEI;
  assign metaArray_0_io_w_setIdx = s2_pipeline_addr[9:4];
  assign metaArray_0_io_w_data_tag = s2_pipeline_addr[31:10];
  assign metaArray_0_io_w_data_valid = 1'h1;
  assign metaArray_0_io_w_data_needFlush = 1'h0;
  assign metaArray_0_io_w_wen = cacheUpdate & 2'h0 == selTree_io_outIdx;
  assign metaArray_0_io_r_setIdx = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign metaArray_0_io_r_ren = ~cacheUpdate;
  assign metaArray_1_clock = clock;
  assign metaArray_1_reset = reset | difftestFENCEI;
  assign metaArray_1_io_w_setIdx = s2_pipeline_addr[9:4];
  assign metaArray_1_io_w_data_tag = s2_pipeline_addr[31:10];
  assign metaArray_1_io_w_data_valid = 1'h1;
  assign metaArray_1_io_w_data_needFlush = 1'h0;
  assign metaArray_1_io_w_wen = cacheUpdate & 2'h1 == selTree_io_outIdx;
  assign metaArray_1_io_r_setIdx = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign metaArray_1_io_r_ren = ~cacheUpdate;
  assign metaArray_2_clock = clock;
  assign metaArray_2_reset = reset | difftestFENCEI;
  assign metaArray_2_io_w_setIdx = s2_pipeline_addr[9:4];
  assign metaArray_2_io_w_data_tag = s2_pipeline_addr[31:10];
  assign metaArray_2_io_w_data_valid = 1'h1;
  assign metaArray_2_io_w_data_needFlush = 1'h0;
  assign metaArray_2_io_w_wen = cacheUpdate & 2'h2 == selTree_io_outIdx;
  assign metaArray_2_io_r_setIdx = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign metaArray_2_io_r_ren = ~cacheUpdate;
  assign metaArray_3_clock = clock;
  assign metaArray_3_reset = reset | difftestFENCEI;
  assign metaArray_3_io_w_setIdx = s2_pipeline_addr[9:4];
  assign metaArray_3_io_w_data_tag = s2_pipeline_addr[31:10];
  assign metaArray_3_io_w_data_valid = 1'h1;
  assign metaArray_3_io_w_data_needFlush = 1'h0;
  assign metaArray_3_io_w_wen = cacheUpdate & 2'h3 == selTree_io_outIdx;
  assign metaArray_3_io_r_setIdx = s2_stall ? s2_pipeline_addr[9:4] : io_in_req_bits_addr[9:4];
  assign metaArray_3_io_r_ren = ~cacheUpdate;
  assign selTree_io_inWayValid_0 = metaArray_0_io_r_data_valid;
  assign selTree_io_inWayValid_1 = metaArray_1_io_r_data_valid;
  assign selTree_io_inWayValid_2 = metaArray_2_io_r_data_valid;
  assign selTree_io_inWayValid_3 = metaArray_3_io_r_data_valid;
  assign selTree_io_inValue_0 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_0 : _GEN_70;
  assign selTree_io_inValue_1 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_1 : _GEN_134;
  assign selTree_io_inValue_2 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_2 : _GEN_198;
  assign selTree_io_inValue_3 = 6'h3f == s2_pipeline_addr[9:4] ? regCount_63_3 : _GEN_262;
  always @(posedge clock) begin
    if (reset) begin
      icache_status <= 3'h0;
    end else if (3'h0 == icache_status) begin
      if (s2_isMMIO) begin
        icache_status <= 3'h5;
      end else if (s2_miss) begin
        icache_status <= _GEN_268;
      end
    end else if (3'h1 == icache_status) begin
      if (_T_23) begin
        icache_status <= 3'h2;
      end
    end else if (3'h2 == icache_status) begin
      icache_status <= _GEN_272;
    end else begin
      icache_status <= _GEN_282;
    end
    if (reset) begin
      regCount_0_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_0_0 <= newCountRefill_0;
        end else begin
          regCount_0_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_0_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_0_1 <= newCountRefill_1;
        end else begin
          regCount_0_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_0_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_0_2 <= newCountRefill_2;
        end else begin
          regCount_0_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_0_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_0_3 <= newCountRefill_3;
        end else begin
          regCount_0_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_1_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_1_0 <= newCountRefill_0;
        end else begin
          regCount_1_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_1_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_1_1 <= newCountRefill_1;
        end else begin
          regCount_1_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_1_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_1_2 <= newCountRefill_2;
        end else begin
          regCount_1_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_1_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_1_3 <= newCountRefill_3;
        end else begin
          regCount_1_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_2_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_2_0 <= newCountRefill_0;
        end else begin
          regCount_2_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_2_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_2_1 <= newCountRefill_1;
        end else begin
          regCount_2_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_2_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_2_2 <= newCountRefill_2;
        end else begin
          regCount_2_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_2_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_2_3 <= newCountRefill_3;
        end else begin
          regCount_2_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_3_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_3_0 <= newCountRefill_0;
        end else begin
          regCount_3_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_3_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_3_1 <= newCountRefill_1;
        end else begin
          regCount_3_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_3_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_3_2 <= newCountRefill_2;
        end else begin
          regCount_3_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_3_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_3_3 <= newCountRefill_3;
        end else begin
          regCount_3_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_4_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_4_0 <= newCountRefill_0;
        end else begin
          regCount_4_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_4_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_4_1 <= newCountRefill_1;
        end else begin
          regCount_4_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_4_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_4_2 <= newCountRefill_2;
        end else begin
          regCount_4_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_4_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_4_3 <= newCountRefill_3;
        end else begin
          regCount_4_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_5_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_5_0 <= newCountRefill_0;
        end else begin
          regCount_5_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_5_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_5_1 <= newCountRefill_1;
        end else begin
          regCount_5_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_5_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_5_2 <= newCountRefill_2;
        end else begin
          regCount_5_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_5_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_5_3 <= newCountRefill_3;
        end else begin
          regCount_5_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_6_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_6_0 <= newCountRefill_0;
        end else begin
          regCount_6_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_6_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_6_1 <= newCountRefill_1;
        end else begin
          regCount_6_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_6_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_6_2 <= newCountRefill_2;
        end else begin
          regCount_6_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_6_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_6_3 <= newCountRefill_3;
        end else begin
          regCount_6_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_7_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_7_0 <= newCountRefill_0;
        end else begin
          regCount_7_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_7_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_7_1 <= newCountRefill_1;
        end else begin
          regCount_7_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_7_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_7_2 <= newCountRefill_2;
        end else begin
          regCount_7_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_7_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_7_3 <= newCountRefill_3;
        end else begin
          regCount_7_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_8_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_8_0 <= newCountRefill_0;
        end else begin
          regCount_8_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_8_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_8_1 <= newCountRefill_1;
        end else begin
          regCount_8_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_8_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_8_2 <= newCountRefill_2;
        end else begin
          regCount_8_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_8_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_8_3 <= newCountRefill_3;
        end else begin
          regCount_8_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_9_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_9_0 <= newCountRefill_0;
        end else begin
          regCount_9_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_9_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_9_1 <= newCountRefill_1;
        end else begin
          regCount_9_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_9_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_9_2 <= newCountRefill_2;
        end else begin
          regCount_9_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_9_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_9_3 <= newCountRefill_3;
        end else begin
          regCount_9_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_10_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_10_0 <= newCountRefill_0;
        end else begin
          regCount_10_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_10_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_10_1 <= newCountRefill_1;
        end else begin
          regCount_10_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_10_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_10_2 <= newCountRefill_2;
        end else begin
          regCount_10_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_10_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_10_3 <= newCountRefill_3;
        end else begin
          regCount_10_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_11_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_11_0 <= newCountRefill_0;
        end else begin
          regCount_11_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_11_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_11_1 <= newCountRefill_1;
        end else begin
          regCount_11_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_11_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_11_2 <= newCountRefill_2;
        end else begin
          regCount_11_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_11_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_11_3 <= newCountRefill_3;
        end else begin
          regCount_11_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_12_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_12_0 <= newCountRefill_0;
        end else begin
          regCount_12_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_12_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_12_1 <= newCountRefill_1;
        end else begin
          regCount_12_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_12_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_12_2 <= newCountRefill_2;
        end else begin
          regCount_12_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_12_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_12_3 <= newCountRefill_3;
        end else begin
          regCount_12_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_13_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_13_0 <= newCountRefill_0;
        end else begin
          regCount_13_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_13_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_13_1 <= newCountRefill_1;
        end else begin
          regCount_13_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_13_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_13_2 <= newCountRefill_2;
        end else begin
          regCount_13_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_13_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_13_3 <= newCountRefill_3;
        end else begin
          regCount_13_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_14_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_14_0 <= newCountRefill_0;
        end else begin
          regCount_14_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_14_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_14_1 <= newCountRefill_1;
        end else begin
          regCount_14_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_14_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_14_2 <= newCountRefill_2;
        end else begin
          regCount_14_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_14_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_14_3 <= newCountRefill_3;
        end else begin
          regCount_14_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_15_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_15_0 <= newCountRefill_0;
        end else begin
          regCount_15_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_15_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_15_1 <= newCountRefill_1;
        end else begin
          regCount_15_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_15_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_15_2 <= newCountRefill_2;
        end else begin
          regCount_15_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_15_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_15_3 <= newCountRefill_3;
        end else begin
          regCount_15_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_16_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_16_0 <= newCountRefill_0;
        end else begin
          regCount_16_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_16_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_16_1 <= newCountRefill_1;
        end else begin
          regCount_16_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_16_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_16_2 <= newCountRefill_2;
        end else begin
          regCount_16_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_16_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_16_3 <= newCountRefill_3;
        end else begin
          regCount_16_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_17_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_17_0 <= newCountRefill_0;
        end else begin
          regCount_17_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_17_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_17_1 <= newCountRefill_1;
        end else begin
          regCount_17_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_17_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_17_2 <= newCountRefill_2;
        end else begin
          regCount_17_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_17_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_17_3 <= newCountRefill_3;
        end else begin
          regCount_17_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_18_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_18_0 <= newCountRefill_0;
        end else begin
          regCount_18_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_18_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_18_1 <= newCountRefill_1;
        end else begin
          regCount_18_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_18_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_18_2 <= newCountRefill_2;
        end else begin
          regCount_18_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_18_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_18_3 <= newCountRefill_3;
        end else begin
          regCount_18_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_19_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_19_0 <= newCountRefill_0;
        end else begin
          regCount_19_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_19_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_19_1 <= newCountRefill_1;
        end else begin
          regCount_19_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_19_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_19_2 <= newCountRefill_2;
        end else begin
          regCount_19_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_19_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_19_3 <= newCountRefill_3;
        end else begin
          regCount_19_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_20_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_20_0 <= newCountRefill_0;
        end else begin
          regCount_20_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_20_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_20_1 <= newCountRefill_1;
        end else begin
          regCount_20_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_20_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_20_2 <= newCountRefill_2;
        end else begin
          regCount_20_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_20_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_20_3 <= newCountRefill_3;
        end else begin
          regCount_20_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_21_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_21_0 <= newCountRefill_0;
        end else begin
          regCount_21_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_21_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_21_1 <= newCountRefill_1;
        end else begin
          regCount_21_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_21_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_21_2 <= newCountRefill_2;
        end else begin
          regCount_21_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_21_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_21_3 <= newCountRefill_3;
        end else begin
          regCount_21_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_22_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_22_0 <= newCountRefill_0;
        end else begin
          regCount_22_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_22_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_22_1 <= newCountRefill_1;
        end else begin
          regCount_22_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_22_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_22_2 <= newCountRefill_2;
        end else begin
          regCount_22_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_22_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_22_3 <= newCountRefill_3;
        end else begin
          regCount_22_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_23_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_23_0 <= newCountRefill_0;
        end else begin
          regCount_23_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_23_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_23_1 <= newCountRefill_1;
        end else begin
          regCount_23_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_23_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_23_2 <= newCountRefill_2;
        end else begin
          regCount_23_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_23_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_23_3 <= newCountRefill_3;
        end else begin
          regCount_23_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_24_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_24_0 <= newCountRefill_0;
        end else begin
          regCount_24_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_24_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_24_1 <= newCountRefill_1;
        end else begin
          regCount_24_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_24_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_24_2 <= newCountRefill_2;
        end else begin
          regCount_24_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_24_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_24_3 <= newCountRefill_3;
        end else begin
          regCount_24_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_25_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_25_0 <= newCountRefill_0;
        end else begin
          regCount_25_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_25_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_25_1 <= newCountRefill_1;
        end else begin
          regCount_25_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_25_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_25_2 <= newCountRefill_2;
        end else begin
          regCount_25_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_25_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_25_3 <= newCountRefill_3;
        end else begin
          regCount_25_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_26_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_26_0 <= newCountRefill_0;
        end else begin
          regCount_26_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_26_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_26_1 <= newCountRefill_1;
        end else begin
          regCount_26_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_26_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_26_2 <= newCountRefill_2;
        end else begin
          regCount_26_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_26_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_26_3 <= newCountRefill_3;
        end else begin
          regCount_26_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_27_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_27_0 <= newCountRefill_0;
        end else begin
          regCount_27_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_27_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_27_1 <= newCountRefill_1;
        end else begin
          regCount_27_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_27_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_27_2 <= newCountRefill_2;
        end else begin
          regCount_27_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_27_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_27_3 <= newCountRefill_3;
        end else begin
          regCount_27_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_28_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_28_0 <= newCountRefill_0;
        end else begin
          regCount_28_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_28_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_28_1 <= newCountRefill_1;
        end else begin
          regCount_28_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_28_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_28_2 <= newCountRefill_2;
        end else begin
          regCount_28_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_28_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_28_3 <= newCountRefill_3;
        end else begin
          regCount_28_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_29_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_29_0 <= newCountRefill_0;
        end else begin
          regCount_29_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_29_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_29_1 <= newCountRefill_1;
        end else begin
          regCount_29_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_29_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_29_2 <= newCountRefill_2;
        end else begin
          regCount_29_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_29_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_29_3 <= newCountRefill_3;
        end else begin
          regCount_29_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_30_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_30_0 <= newCountRefill_0;
        end else begin
          regCount_30_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_30_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_30_1 <= newCountRefill_1;
        end else begin
          regCount_30_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_30_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_30_2 <= newCountRefill_2;
        end else begin
          regCount_30_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_30_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_30_3 <= newCountRefill_3;
        end else begin
          regCount_30_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_31_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_31_0 <= newCountRefill_0;
        end else begin
          regCount_31_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_31_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_31_1 <= newCountRefill_1;
        end else begin
          regCount_31_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_31_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_31_2 <= newCountRefill_2;
        end else begin
          regCount_31_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_31_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_31_3 <= newCountRefill_3;
        end else begin
          regCount_31_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_32_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_32_0 <= newCountRefill_0;
        end else begin
          regCount_32_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_32_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_32_1 <= newCountRefill_1;
        end else begin
          regCount_32_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_32_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_32_2 <= newCountRefill_2;
        end else begin
          regCount_32_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_32_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_32_3 <= newCountRefill_3;
        end else begin
          regCount_32_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_33_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_33_0 <= newCountRefill_0;
        end else begin
          regCount_33_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_33_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_33_1 <= newCountRefill_1;
        end else begin
          regCount_33_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_33_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_33_2 <= newCountRefill_2;
        end else begin
          regCount_33_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_33_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_33_3 <= newCountRefill_3;
        end else begin
          regCount_33_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_34_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_34_0 <= newCountRefill_0;
        end else begin
          regCount_34_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_34_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_34_1 <= newCountRefill_1;
        end else begin
          regCount_34_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_34_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_34_2 <= newCountRefill_2;
        end else begin
          regCount_34_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_34_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_34_3 <= newCountRefill_3;
        end else begin
          regCount_34_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_35_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_35_0 <= newCountRefill_0;
        end else begin
          regCount_35_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_35_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_35_1 <= newCountRefill_1;
        end else begin
          regCount_35_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_35_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_35_2 <= newCountRefill_2;
        end else begin
          regCount_35_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_35_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_35_3 <= newCountRefill_3;
        end else begin
          regCount_35_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_36_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_36_0 <= newCountRefill_0;
        end else begin
          regCount_36_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_36_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_36_1 <= newCountRefill_1;
        end else begin
          regCount_36_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_36_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_36_2 <= newCountRefill_2;
        end else begin
          regCount_36_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_36_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_36_3 <= newCountRefill_3;
        end else begin
          regCount_36_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_37_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_37_0 <= newCountRefill_0;
        end else begin
          regCount_37_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_37_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_37_1 <= newCountRefill_1;
        end else begin
          regCount_37_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_37_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_37_2 <= newCountRefill_2;
        end else begin
          regCount_37_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_37_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_37_3 <= newCountRefill_3;
        end else begin
          regCount_37_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_38_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_38_0 <= newCountRefill_0;
        end else begin
          regCount_38_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_38_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_38_1 <= newCountRefill_1;
        end else begin
          regCount_38_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_38_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_38_2 <= newCountRefill_2;
        end else begin
          regCount_38_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_38_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_38_3 <= newCountRefill_3;
        end else begin
          regCount_38_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_39_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_39_0 <= newCountRefill_0;
        end else begin
          regCount_39_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_39_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_39_1 <= newCountRefill_1;
        end else begin
          regCount_39_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_39_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_39_2 <= newCountRefill_2;
        end else begin
          regCount_39_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_39_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_39_3 <= newCountRefill_3;
        end else begin
          regCount_39_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_40_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_40_0 <= newCountRefill_0;
        end else begin
          regCount_40_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_40_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_40_1 <= newCountRefill_1;
        end else begin
          regCount_40_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_40_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_40_2 <= newCountRefill_2;
        end else begin
          regCount_40_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_40_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_40_3 <= newCountRefill_3;
        end else begin
          regCount_40_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_41_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_41_0 <= newCountRefill_0;
        end else begin
          regCount_41_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_41_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_41_1 <= newCountRefill_1;
        end else begin
          regCount_41_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_41_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_41_2 <= newCountRefill_2;
        end else begin
          regCount_41_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_41_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_41_3 <= newCountRefill_3;
        end else begin
          regCount_41_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_42_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_42_0 <= newCountRefill_0;
        end else begin
          regCount_42_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_42_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_42_1 <= newCountRefill_1;
        end else begin
          regCount_42_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_42_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_42_2 <= newCountRefill_2;
        end else begin
          regCount_42_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_42_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_42_3 <= newCountRefill_3;
        end else begin
          regCount_42_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_43_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_43_0 <= newCountRefill_0;
        end else begin
          regCount_43_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_43_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_43_1 <= newCountRefill_1;
        end else begin
          regCount_43_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_43_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_43_2 <= newCountRefill_2;
        end else begin
          regCount_43_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_43_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_43_3 <= newCountRefill_3;
        end else begin
          regCount_43_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_44_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_44_0 <= newCountRefill_0;
        end else begin
          regCount_44_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_44_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_44_1 <= newCountRefill_1;
        end else begin
          regCount_44_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_44_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_44_2 <= newCountRefill_2;
        end else begin
          regCount_44_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_44_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_44_3 <= newCountRefill_3;
        end else begin
          regCount_44_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_45_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_45_0 <= newCountRefill_0;
        end else begin
          regCount_45_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_45_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_45_1 <= newCountRefill_1;
        end else begin
          regCount_45_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_45_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_45_2 <= newCountRefill_2;
        end else begin
          regCount_45_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_45_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_45_3 <= newCountRefill_3;
        end else begin
          regCount_45_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_46_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_46_0 <= newCountRefill_0;
        end else begin
          regCount_46_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_46_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_46_1 <= newCountRefill_1;
        end else begin
          regCount_46_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_46_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_46_2 <= newCountRefill_2;
        end else begin
          regCount_46_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_46_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_46_3 <= newCountRefill_3;
        end else begin
          regCount_46_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_47_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_47_0 <= newCountRefill_0;
        end else begin
          regCount_47_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_47_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_47_1 <= newCountRefill_1;
        end else begin
          regCount_47_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_47_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_47_2 <= newCountRefill_2;
        end else begin
          regCount_47_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_47_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_47_3 <= newCountRefill_3;
        end else begin
          regCount_47_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_48_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_48_0 <= newCountRefill_0;
        end else begin
          regCount_48_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_48_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_48_1 <= newCountRefill_1;
        end else begin
          regCount_48_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_48_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_48_2 <= newCountRefill_2;
        end else begin
          regCount_48_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_48_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_48_3 <= newCountRefill_3;
        end else begin
          regCount_48_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_49_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_49_0 <= newCountRefill_0;
        end else begin
          regCount_49_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_49_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_49_1 <= newCountRefill_1;
        end else begin
          regCount_49_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_49_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_49_2 <= newCountRefill_2;
        end else begin
          regCount_49_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_49_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_49_3 <= newCountRefill_3;
        end else begin
          regCount_49_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_50_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_50_0 <= newCountRefill_0;
        end else begin
          regCount_50_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_50_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_50_1 <= newCountRefill_1;
        end else begin
          regCount_50_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_50_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_50_2 <= newCountRefill_2;
        end else begin
          regCount_50_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_50_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_50_3 <= newCountRefill_3;
        end else begin
          regCount_50_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_51_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_51_0 <= newCountRefill_0;
        end else begin
          regCount_51_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_51_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_51_1 <= newCountRefill_1;
        end else begin
          regCount_51_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_51_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_51_2 <= newCountRefill_2;
        end else begin
          regCount_51_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_51_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_51_3 <= newCountRefill_3;
        end else begin
          regCount_51_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_52_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_52_0 <= newCountRefill_0;
        end else begin
          regCount_52_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_52_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_52_1 <= newCountRefill_1;
        end else begin
          regCount_52_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_52_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_52_2 <= newCountRefill_2;
        end else begin
          regCount_52_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_52_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_52_3 <= newCountRefill_3;
        end else begin
          regCount_52_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_53_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_53_0 <= newCountRefill_0;
        end else begin
          regCount_53_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_53_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_53_1 <= newCountRefill_1;
        end else begin
          regCount_53_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_53_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_53_2 <= newCountRefill_2;
        end else begin
          regCount_53_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_53_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_53_3 <= newCountRefill_3;
        end else begin
          regCount_53_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_54_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_54_0 <= newCountRefill_0;
        end else begin
          regCount_54_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_54_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_54_1 <= newCountRefill_1;
        end else begin
          regCount_54_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_54_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_54_2 <= newCountRefill_2;
        end else begin
          regCount_54_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_54_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_54_3 <= newCountRefill_3;
        end else begin
          regCount_54_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_55_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_55_0 <= newCountRefill_0;
        end else begin
          regCount_55_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_55_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_55_1 <= newCountRefill_1;
        end else begin
          regCount_55_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_55_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_55_2 <= newCountRefill_2;
        end else begin
          regCount_55_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_55_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_55_3 <= newCountRefill_3;
        end else begin
          regCount_55_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_56_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_56_0 <= newCountRefill_0;
        end else begin
          regCount_56_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_56_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_56_1 <= newCountRefill_1;
        end else begin
          regCount_56_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_56_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_56_2 <= newCountRefill_2;
        end else begin
          regCount_56_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_56_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_56_3 <= newCountRefill_3;
        end else begin
          regCount_56_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_57_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_57_0 <= newCountRefill_0;
        end else begin
          regCount_57_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_57_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_57_1 <= newCountRefill_1;
        end else begin
          regCount_57_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_57_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_57_2 <= newCountRefill_2;
        end else begin
          regCount_57_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_57_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_57_3 <= newCountRefill_3;
        end else begin
          regCount_57_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_58_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_58_0 <= newCountRefill_0;
        end else begin
          regCount_58_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_58_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_58_1 <= newCountRefill_1;
        end else begin
          regCount_58_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_58_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_58_2 <= newCountRefill_2;
        end else begin
          regCount_58_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_58_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_58_3 <= newCountRefill_3;
        end else begin
          regCount_58_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_59_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_59_0 <= newCountRefill_0;
        end else begin
          regCount_59_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_59_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_59_1 <= newCountRefill_1;
        end else begin
          regCount_59_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_59_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_59_2 <= newCountRefill_2;
        end else begin
          regCount_59_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_59_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_59_3 <= newCountRefill_3;
        end else begin
          regCount_59_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_60_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_60_0 <= newCountRefill_0;
        end else begin
          regCount_60_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_60_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_60_1 <= newCountRefill_1;
        end else begin
          regCount_60_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_60_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_60_2 <= newCountRefill_2;
        end else begin
          regCount_60_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_60_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_60_3 <= newCountRefill_3;
        end else begin
          regCount_60_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_61_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_61_0 <= newCountRefill_0;
        end else begin
          regCount_61_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_61_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_61_1 <= newCountRefill_1;
        end else begin
          regCount_61_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_61_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_61_2 <= newCountRefill_2;
        end else begin
          regCount_61_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_61_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_61_3 <= newCountRefill_3;
        end else begin
          regCount_61_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_62_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_62_0 <= newCountRefill_0;
        end else begin
          regCount_62_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_62_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_62_1 <= newCountRefill_1;
        end else begin
          regCount_62_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_62_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_62_2 <= newCountRefill_2;
        end else begin
          regCount_62_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_62_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_62_3 <= newCountRefill_3;
        end else begin
          regCount_62_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_63_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_63_0 <= newCountRefill_0;
        end else begin
          regCount_63_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_63_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_63_1 <= newCountRefill_1;
        end else begin
          regCount_63_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_63_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_63_2 <= newCountRefill_2;
        end else begin
          regCount_63_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_63_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == s2_pipeline_addr[9:4]) begin
        if (cacheUpdate) begin
          regCount_63_3 <= newCountRefill_3;
        end else begin
          regCount_63_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      s2_pipeline_valid <= 1'h0;
    end else begin
      s2_pipeline_valid <= _GEN_4;
    end
    if (reset) begin
      s2_pipeline_addr <= 32'h0;
    end else if (~s2_stall) begin
      s2_pipeline_addr <= io_in_req_bits_addr;
    end
    if (reset) begin
      s2_pipeline_size <= 2'h0;
    end else if (~s2_stall) begin
      s2_pipeline_size <= 2'h2;
    end
    if (reset) begin
      s2_pipeline_isMMIO <= 1'h0;
    end else if (~s2_stall) begin
      s2_pipeline_isMMIO <= s1_isMMIO_hit;
    end
    if (_T_33) begin
      mmioRespData <= io_mmio_resp_bits_rdata;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  icache_status = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  regCount_0_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  regCount_0_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  regCount_0_2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  regCount_0_3 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  regCount_1_0 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  regCount_1_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  regCount_1_2 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  regCount_1_3 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  regCount_2_0 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  regCount_2_1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  regCount_2_2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  regCount_2_3 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  regCount_3_0 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  regCount_3_1 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  regCount_3_2 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  regCount_3_3 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  regCount_4_0 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  regCount_4_1 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  regCount_4_2 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  regCount_4_3 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  regCount_5_0 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  regCount_5_1 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  regCount_5_2 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  regCount_5_3 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  regCount_6_0 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  regCount_6_1 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  regCount_6_2 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  regCount_6_3 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  regCount_7_0 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  regCount_7_1 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  regCount_7_2 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  regCount_7_3 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  regCount_8_0 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  regCount_8_1 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  regCount_8_2 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  regCount_8_3 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  regCount_9_0 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  regCount_9_1 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  regCount_9_2 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  regCount_9_3 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  regCount_10_0 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  regCount_10_1 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  regCount_10_2 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  regCount_10_3 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  regCount_11_0 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  regCount_11_1 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  regCount_11_2 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  regCount_11_3 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  regCount_12_0 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  regCount_12_1 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  regCount_12_2 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  regCount_12_3 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  regCount_13_0 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  regCount_13_1 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  regCount_13_2 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  regCount_13_3 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  regCount_14_0 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  regCount_14_1 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  regCount_14_2 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  regCount_14_3 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  regCount_15_0 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  regCount_15_1 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  regCount_15_2 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  regCount_15_3 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  regCount_16_0 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  regCount_16_1 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  regCount_16_2 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  regCount_16_3 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  regCount_17_0 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  regCount_17_1 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  regCount_17_2 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  regCount_17_3 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  regCount_18_0 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  regCount_18_1 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  regCount_18_2 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  regCount_18_3 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  regCount_19_0 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  regCount_19_1 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  regCount_19_2 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  regCount_19_3 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  regCount_20_0 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  regCount_20_1 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  regCount_20_2 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  regCount_20_3 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  regCount_21_0 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  regCount_21_1 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  regCount_21_2 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  regCount_21_3 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  regCount_22_0 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  regCount_22_1 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  regCount_22_2 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  regCount_22_3 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  regCount_23_0 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  regCount_23_1 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  regCount_23_2 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  regCount_23_3 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  regCount_24_0 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  regCount_24_1 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  regCount_24_2 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  regCount_24_3 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  regCount_25_0 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  regCount_25_1 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  regCount_25_2 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  regCount_25_3 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  regCount_26_0 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  regCount_26_1 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  regCount_26_2 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  regCount_26_3 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  regCount_27_0 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  regCount_27_1 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  regCount_27_2 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  regCount_27_3 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  regCount_28_0 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  regCount_28_1 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  regCount_28_2 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  regCount_28_3 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  regCount_29_0 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  regCount_29_1 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  regCount_29_2 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  regCount_29_3 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  regCount_30_0 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  regCount_30_1 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  regCount_30_2 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  regCount_30_3 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  regCount_31_0 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  regCount_31_1 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  regCount_31_2 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  regCount_31_3 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  regCount_32_0 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  regCount_32_1 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  regCount_32_2 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  regCount_32_3 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  regCount_33_0 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  regCount_33_1 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  regCount_33_2 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  regCount_33_3 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  regCount_34_0 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  regCount_34_1 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  regCount_34_2 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  regCount_34_3 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  regCount_35_0 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  regCount_35_1 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  regCount_35_2 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  regCount_35_3 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  regCount_36_0 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  regCount_36_1 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  regCount_36_2 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  regCount_36_3 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  regCount_37_0 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  regCount_37_1 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  regCount_37_2 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  regCount_37_3 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  regCount_38_0 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  regCount_38_1 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  regCount_38_2 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  regCount_38_3 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  regCount_39_0 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  regCount_39_1 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  regCount_39_2 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  regCount_39_3 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  regCount_40_0 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  regCount_40_1 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  regCount_40_2 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  regCount_40_3 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  regCount_41_0 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  regCount_41_1 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  regCount_41_2 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  regCount_41_3 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  regCount_42_0 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  regCount_42_1 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  regCount_42_2 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  regCount_42_3 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  regCount_43_0 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  regCount_43_1 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  regCount_43_2 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  regCount_43_3 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  regCount_44_0 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  regCount_44_1 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  regCount_44_2 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  regCount_44_3 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  regCount_45_0 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  regCount_45_1 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  regCount_45_2 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  regCount_45_3 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  regCount_46_0 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  regCount_46_1 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  regCount_46_2 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  regCount_46_3 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  regCount_47_0 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  regCount_47_1 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  regCount_47_2 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  regCount_47_3 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  regCount_48_0 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  regCount_48_1 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  regCount_48_2 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  regCount_48_3 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  regCount_49_0 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  regCount_49_1 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  regCount_49_2 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  regCount_49_3 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  regCount_50_0 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  regCount_50_1 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  regCount_50_2 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  regCount_50_3 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  regCount_51_0 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  regCount_51_1 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  regCount_51_2 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  regCount_51_3 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  regCount_52_0 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  regCount_52_1 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  regCount_52_2 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  regCount_52_3 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  regCount_53_0 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  regCount_53_1 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  regCount_53_2 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  regCount_53_3 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  regCount_54_0 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  regCount_54_1 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  regCount_54_2 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  regCount_54_3 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  regCount_55_0 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  regCount_55_1 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  regCount_55_2 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  regCount_55_3 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  regCount_56_0 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  regCount_56_1 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  regCount_56_2 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  regCount_56_3 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  regCount_57_0 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  regCount_57_1 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  regCount_57_2 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  regCount_57_3 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  regCount_58_0 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  regCount_58_1 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  regCount_58_2 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  regCount_58_3 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  regCount_59_0 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  regCount_59_1 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  regCount_59_2 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  regCount_59_3 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  regCount_60_0 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  regCount_60_1 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  regCount_60_2 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  regCount_60_3 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  regCount_61_0 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  regCount_61_1 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  regCount_61_2 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  regCount_61_3 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  regCount_62_0 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  regCount_62_1 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  regCount_62_2 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  regCount_62_3 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  regCount_63_0 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  regCount_63_1 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  regCount_63_2 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  regCount_63_3 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  s2_pipeline_valid = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  s2_pipeline_addr = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  s2_pipeline_size = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  s2_pipeline_isMMIO = _RAND_260[0:0];
  _RAND_261 = {2{`RANDOM}};
  mmioRespData = _RAND_261[63:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Arbiter(
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_addr,
  input  [127:0] io_in_0_bits_wdata,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [31:0]  io_in_1_bits_addr,
  input  [127:0] io_in_1_bits_wdata,
  input  [1:0]   io_in_1_bits_size,
  input  [2:0]   io_in_1_bits_cmd,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [127:0] io_out_bits_wdata,
  output [1:0]   io_out_bits_size,
  output [2:0]   io_out_bits_cmd
);
  wire  grant_1 = ~io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = grant_1 & io_out_ready;
  assign io_out_valid = ~grant_1 | io_in_1_valid;
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata;
  assign io_out_bits_size = io_in_0_valid ? 2'h3 : io_in_1_bits_size;
  assign io_out_bits_cmd = io_in_0_valid ? 3'h2 : io_in_1_bits_cmd;
endmodule
module ysyx_040656_DCache(
  input          clock,
  input          reset,
  output         io_in_req_ready,
  input          io_in_req_valid,
  input  [31:0]  io_in_req_bits_addr,
  input  [63:0]  io_in_req_bits_wdata,
  input  [1:0]   io_in_req_bits_size,
  input  [2:0]   io_in_req_bits_cmd,
  output         io_in_resp_valid,
  output [63:0]  io_in_resp_bits_rdata,
  input          io_out_req_ready,
  output         io_out_req_valid,
  output [31:0]  io_out_req_bits_addr,
  output [127:0] io_out_req_bits_wdata,
  output [2:0]   io_out_req_bits_cmd,
  output         io_out_resp_ready,
  input          io_out_resp_valid,
  input  [127:0] io_out_resp_bits_rdata,
  output         io_link_req_ready,
  input          io_link_req_valid,
  input  [31:0]  io_link_req_bits_addr,
  input  [127:0] io_link_req_bits_wdata,
  output         io_link_resp_valid,
  output [2:0]   io_link_resp_bits_cmd,
  output [127:0] io_link_resp_bits_rdata,
  input  [127:0] io_dataArray_0_rdata,
  output         io_dataArray_0_wen,
  output [5:0]   io_dataArray_0_addr,
  output [127:0] io_dataArray_0_wdata,
  input  [127:0] io_dataArray_1_rdata,
  output         io_dataArray_1_wen,
  output [5:0]   io_dataArray_1_addr,
  output [127:0] io_dataArray_1_wdata,
  input  [127:0] io_dataArray_2_rdata,
  output         io_dataArray_2_wen,
  output [5:0]   io_dataArray_2_addr,
  output [127:0] io_dataArray_2_wdata,
  input  [127:0] io_dataArray_3_rdata,
  output         io_dataArray_3_wen,
  output [5:0]   io_dataArray_3_addr,
  output [127:0] io_dataArray_3_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
`endif
  wire  metaArray_0_clock;
  wire  metaArray_0_reset;
  wire [5:0] metaArray_0_io_w_setIdx;
  wire [21:0] metaArray_0_io_w_data_tag;
  wire  metaArray_0_io_w_data_valid;
  wire  metaArray_0_io_w_data_needFlush;
  wire  metaArray_0_io_w_wen;
  wire [5:0] metaArray_0_io_r_setIdx;
  wire [21:0] metaArray_0_io_r_data_tag;
  wire  metaArray_0_io_r_data_valid;
  wire  metaArray_0_io_r_data_needFlush;
  wire  metaArray_0_io_r_ren;
  wire  metaArray_1_clock;
  wire  metaArray_1_reset;
  wire [5:0] metaArray_1_io_w_setIdx;
  wire [21:0] metaArray_1_io_w_data_tag;
  wire  metaArray_1_io_w_data_valid;
  wire  metaArray_1_io_w_data_needFlush;
  wire  metaArray_1_io_w_wen;
  wire [5:0] metaArray_1_io_r_setIdx;
  wire [21:0] metaArray_1_io_r_data_tag;
  wire  metaArray_1_io_r_data_valid;
  wire  metaArray_1_io_r_data_needFlush;
  wire  metaArray_1_io_r_ren;
  wire  metaArray_2_clock;
  wire  metaArray_2_reset;
  wire [5:0] metaArray_2_io_w_setIdx;
  wire [21:0] metaArray_2_io_w_data_tag;
  wire  metaArray_2_io_w_data_valid;
  wire  metaArray_2_io_w_data_needFlush;
  wire  metaArray_2_io_w_wen;
  wire [5:0] metaArray_2_io_r_setIdx;
  wire [21:0] metaArray_2_io_r_data_tag;
  wire  metaArray_2_io_r_data_valid;
  wire  metaArray_2_io_r_data_needFlush;
  wire  metaArray_2_io_r_ren;
  wire  metaArray_3_clock;
  wire  metaArray_3_reset;
  wire [5:0] metaArray_3_io_w_setIdx;
  wire [21:0] metaArray_3_io_w_data_tag;
  wire  metaArray_3_io_w_data_valid;
  wire  metaArray_3_io_w_data_needFlush;
  wire  metaArray_3_io_w_wen;
  wire [5:0] metaArray_3_io_r_setIdx;
  wire [21:0] metaArray_3_io_r_data_tag;
  wire  metaArray_3_io_r_data_valid;
  wire  metaArray_3_io_r_data_needFlush;
  wire  metaArray_3_io_r_ren;
  wire  arbiter_io_in_0_ready;
  wire  arbiter_io_in_0_valid;
  wire [31:0] arbiter_io_in_0_bits_addr;
  wire [127:0] arbiter_io_in_0_bits_wdata;
  wire  arbiter_io_in_1_ready;
  wire  arbiter_io_in_1_valid;
  wire [31:0] arbiter_io_in_1_bits_addr;
  wire [127:0] arbiter_io_in_1_bits_wdata;
  wire [1:0] arbiter_io_in_1_bits_size;
  wire [2:0] arbiter_io_in_1_bits_cmd;
  wire  arbiter_io_out_ready;
  wire  arbiter_io_out_valid;
  wire [31:0] arbiter_io_out_bits_addr;
  wire [127:0] arbiter_io_out_bits_wdata;
  wire [1:0] arbiter_io_out_bits_size;
  wire [2:0] arbiter_io_out_bits_cmd;
  wire  selTree_io_inWayValid_0;
  wire  selTree_io_inWayValid_1;
  wire  selTree_io_inWayValid_2;
  wire  selTree_io_inWayValid_3;
  wire [1:0] selTree_io_inValue_0;
  wire [1:0] selTree_io_inValue_1;
  wire [1:0] selTree_io_inValue_2;
  wire [1:0] selTree_io_inValue_3;
  wire [1:0] selTree_io_outIdx;
  reg [2:0] c_state;
  reg [1:0] regCount_0_0;
  reg [1:0] regCount_0_1;
  reg [1:0] regCount_0_2;
  reg [1:0] regCount_0_3;
  reg [1:0] regCount_1_0;
  reg [1:0] regCount_1_1;
  reg [1:0] regCount_1_2;
  reg [1:0] regCount_1_3;
  reg [1:0] regCount_2_0;
  reg [1:0] regCount_2_1;
  reg [1:0] regCount_2_2;
  reg [1:0] regCount_2_3;
  reg [1:0] regCount_3_0;
  reg [1:0] regCount_3_1;
  reg [1:0] regCount_3_2;
  reg [1:0] regCount_3_3;
  reg [1:0] regCount_4_0;
  reg [1:0] regCount_4_1;
  reg [1:0] regCount_4_2;
  reg [1:0] regCount_4_3;
  reg [1:0] regCount_5_0;
  reg [1:0] regCount_5_1;
  reg [1:0] regCount_5_2;
  reg [1:0] regCount_5_3;
  reg [1:0] regCount_6_0;
  reg [1:0] regCount_6_1;
  reg [1:0] regCount_6_2;
  reg [1:0] regCount_6_3;
  reg [1:0] regCount_7_0;
  reg [1:0] regCount_7_1;
  reg [1:0] regCount_7_2;
  reg [1:0] regCount_7_3;
  reg [1:0] regCount_8_0;
  reg [1:0] regCount_8_1;
  reg [1:0] regCount_8_2;
  reg [1:0] regCount_8_3;
  reg [1:0] regCount_9_0;
  reg [1:0] regCount_9_1;
  reg [1:0] regCount_9_2;
  reg [1:0] regCount_9_3;
  reg [1:0] regCount_10_0;
  reg [1:0] regCount_10_1;
  reg [1:0] regCount_10_2;
  reg [1:0] regCount_10_3;
  reg [1:0] regCount_11_0;
  reg [1:0] regCount_11_1;
  reg [1:0] regCount_11_2;
  reg [1:0] regCount_11_3;
  reg [1:0] regCount_12_0;
  reg [1:0] regCount_12_1;
  reg [1:0] regCount_12_2;
  reg [1:0] regCount_12_3;
  reg [1:0] regCount_13_0;
  reg [1:0] regCount_13_1;
  reg [1:0] regCount_13_2;
  reg [1:0] regCount_13_3;
  reg [1:0] regCount_14_0;
  reg [1:0] regCount_14_1;
  reg [1:0] regCount_14_2;
  reg [1:0] regCount_14_3;
  reg [1:0] regCount_15_0;
  reg [1:0] regCount_15_1;
  reg [1:0] regCount_15_2;
  reg [1:0] regCount_15_3;
  reg [1:0] regCount_16_0;
  reg [1:0] regCount_16_1;
  reg [1:0] regCount_16_2;
  reg [1:0] regCount_16_3;
  reg [1:0] regCount_17_0;
  reg [1:0] regCount_17_1;
  reg [1:0] regCount_17_2;
  reg [1:0] regCount_17_3;
  reg [1:0] regCount_18_0;
  reg [1:0] regCount_18_1;
  reg [1:0] regCount_18_2;
  reg [1:0] regCount_18_3;
  reg [1:0] regCount_19_0;
  reg [1:0] regCount_19_1;
  reg [1:0] regCount_19_2;
  reg [1:0] regCount_19_3;
  reg [1:0] regCount_20_0;
  reg [1:0] regCount_20_1;
  reg [1:0] regCount_20_2;
  reg [1:0] regCount_20_3;
  reg [1:0] regCount_21_0;
  reg [1:0] regCount_21_1;
  reg [1:0] regCount_21_2;
  reg [1:0] regCount_21_3;
  reg [1:0] regCount_22_0;
  reg [1:0] regCount_22_1;
  reg [1:0] regCount_22_2;
  reg [1:0] regCount_22_3;
  reg [1:0] regCount_23_0;
  reg [1:0] regCount_23_1;
  reg [1:0] regCount_23_2;
  reg [1:0] regCount_23_3;
  reg [1:0] regCount_24_0;
  reg [1:0] regCount_24_1;
  reg [1:0] regCount_24_2;
  reg [1:0] regCount_24_3;
  reg [1:0] regCount_25_0;
  reg [1:0] regCount_25_1;
  reg [1:0] regCount_25_2;
  reg [1:0] regCount_25_3;
  reg [1:0] regCount_26_0;
  reg [1:0] regCount_26_1;
  reg [1:0] regCount_26_2;
  reg [1:0] regCount_26_3;
  reg [1:0] regCount_27_0;
  reg [1:0] regCount_27_1;
  reg [1:0] regCount_27_2;
  reg [1:0] regCount_27_3;
  reg [1:0] regCount_28_0;
  reg [1:0] regCount_28_1;
  reg [1:0] regCount_28_2;
  reg [1:0] regCount_28_3;
  reg [1:0] regCount_29_0;
  reg [1:0] regCount_29_1;
  reg [1:0] regCount_29_2;
  reg [1:0] regCount_29_3;
  reg [1:0] regCount_30_0;
  reg [1:0] regCount_30_1;
  reg [1:0] regCount_30_2;
  reg [1:0] regCount_30_3;
  reg [1:0] regCount_31_0;
  reg [1:0] regCount_31_1;
  reg [1:0] regCount_31_2;
  reg [1:0] regCount_31_3;
  reg [1:0] regCount_32_0;
  reg [1:0] regCount_32_1;
  reg [1:0] regCount_32_2;
  reg [1:0] regCount_32_3;
  reg [1:0] regCount_33_0;
  reg [1:0] regCount_33_1;
  reg [1:0] regCount_33_2;
  reg [1:0] regCount_33_3;
  reg [1:0] regCount_34_0;
  reg [1:0] regCount_34_1;
  reg [1:0] regCount_34_2;
  reg [1:0] regCount_34_3;
  reg [1:0] regCount_35_0;
  reg [1:0] regCount_35_1;
  reg [1:0] regCount_35_2;
  reg [1:0] regCount_35_3;
  reg [1:0] regCount_36_0;
  reg [1:0] regCount_36_1;
  reg [1:0] regCount_36_2;
  reg [1:0] regCount_36_3;
  reg [1:0] regCount_37_0;
  reg [1:0] regCount_37_1;
  reg [1:0] regCount_37_2;
  reg [1:0] regCount_37_3;
  reg [1:0] regCount_38_0;
  reg [1:0] regCount_38_1;
  reg [1:0] regCount_38_2;
  reg [1:0] regCount_38_3;
  reg [1:0] regCount_39_0;
  reg [1:0] regCount_39_1;
  reg [1:0] regCount_39_2;
  reg [1:0] regCount_39_3;
  reg [1:0] regCount_40_0;
  reg [1:0] regCount_40_1;
  reg [1:0] regCount_40_2;
  reg [1:0] regCount_40_3;
  reg [1:0] regCount_41_0;
  reg [1:0] regCount_41_1;
  reg [1:0] regCount_41_2;
  reg [1:0] regCount_41_3;
  reg [1:0] regCount_42_0;
  reg [1:0] regCount_42_1;
  reg [1:0] regCount_42_2;
  reg [1:0] regCount_42_3;
  reg [1:0] regCount_43_0;
  reg [1:0] regCount_43_1;
  reg [1:0] regCount_43_2;
  reg [1:0] regCount_43_3;
  reg [1:0] regCount_44_0;
  reg [1:0] regCount_44_1;
  reg [1:0] regCount_44_2;
  reg [1:0] regCount_44_3;
  reg [1:0] regCount_45_0;
  reg [1:0] regCount_45_1;
  reg [1:0] regCount_45_2;
  reg [1:0] regCount_45_3;
  reg [1:0] regCount_46_0;
  reg [1:0] regCount_46_1;
  reg [1:0] regCount_46_2;
  reg [1:0] regCount_46_3;
  reg [1:0] regCount_47_0;
  reg [1:0] regCount_47_1;
  reg [1:0] regCount_47_2;
  reg [1:0] regCount_47_3;
  reg [1:0] regCount_48_0;
  reg [1:0] regCount_48_1;
  reg [1:0] regCount_48_2;
  reg [1:0] regCount_48_3;
  reg [1:0] regCount_49_0;
  reg [1:0] regCount_49_1;
  reg [1:0] regCount_49_2;
  reg [1:0] regCount_49_3;
  reg [1:0] regCount_50_0;
  reg [1:0] regCount_50_1;
  reg [1:0] regCount_50_2;
  reg [1:0] regCount_50_3;
  reg [1:0] regCount_51_0;
  reg [1:0] regCount_51_1;
  reg [1:0] regCount_51_2;
  reg [1:0] regCount_51_3;
  reg [1:0] regCount_52_0;
  reg [1:0] regCount_52_1;
  reg [1:0] regCount_52_2;
  reg [1:0] regCount_52_3;
  reg [1:0] regCount_53_0;
  reg [1:0] regCount_53_1;
  reg [1:0] regCount_53_2;
  reg [1:0] regCount_53_3;
  reg [1:0] regCount_54_0;
  reg [1:0] regCount_54_1;
  reg [1:0] regCount_54_2;
  reg [1:0] regCount_54_3;
  reg [1:0] regCount_55_0;
  reg [1:0] regCount_55_1;
  reg [1:0] regCount_55_2;
  reg [1:0] regCount_55_3;
  reg [1:0] regCount_56_0;
  reg [1:0] regCount_56_1;
  reg [1:0] regCount_56_2;
  reg [1:0] regCount_56_3;
  reg [1:0] regCount_57_0;
  reg [1:0] regCount_57_1;
  reg [1:0] regCount_57_2;
  reg [1:0] regCount_57_3;
  reg [1:0] regCount_58_0;
  reg [1:0] regCount_58_1;
  reg [1:0] regCount_58_2;
  reg [1:0] regCount_58_3;
  reg [1:0] regCount_59_0;
  reg [1:0] regCount_59_1;
  reg [1:0] regCount_59_2;
  reg [1:0] regCount_59_3;
  reg [1:0] regCount_60_0;
  reg [1:0] regCount_60_1;
  reg [1:0] regCount_60_2;
  reg [1:0] regCount_60_3;
  reg [1:0] regCount_61_0;
  reg [1:0] regCount_61_1;
  reg [1:0] regCount_61_2;
  reg [1:0] regCount_61_3;
  reg [1:0] regCount_62_0;
  reg [1:0] regCount_62_1;
  reg [1:0] regCount_62_2;
  reg [1:0] regCount_62_3;
  reg [1:0] regCount_63_0;
  reg [1:0] regCount_63_1;
  reg [1:0] regCount_63_2;
  reg [1:0] regCount_63_3;
  wire  s1_valid = arbiter_io_out_ready & arbiter_io_out_valid;
  reg [31:0] req_addr_r;
  wire [31:0] _GEN_0 = s1_valid ? arbiter_io_out_bits_addr : req_addr_r;
  wire [2:0] req_addr_byteOffset = _GEN_0[2:0];
  wire  req_addr_wordOffest = _GEN_0[3];
  wire [5:0] req_addr_index = _GEN_0[9:4];
  wire [21:0] req_addr_tag = _GEN_0[31:10];
  wire  s1_probe = arbiter_io_out_bits_cmd == 3'h2;
  wire [5:0] shift = {req_addr_byteOffset, 3'h0};
  wire [63:0] s1_wdata = arbiter_io_out_bits_wdata[63:0];
  wire  s1_wen = arbiter_io_out_bits_cmd == 3'h1 | arbiter_io_out_bits_cmd == 3'h4;
  wire [31:0] _s1_strb_T = {req_addr_tag,req_addr_index,req_addr_wordOffest,req_addr_byteOffset};
  wire [3:0] s1_strb_numValid = 4'h1 << arbiter_io_out_bits_size;
  wire [3:0] _GEN_1106 = {{1'd0}, _s1_strb_T[2:0]};
  wire [3:0] _s1_strb_wmask_0_T_4 = _GEN_1106 + s1_strb_numValid;
  wire  s1_strb_wmask_0 = _s1_strb_T[2:0] <= 3'h0 & _s1_strb_wmask_0_T_4 > 4'h0;
  wire  s1_strb_wmask_1 = _s1_strb_T[2:0] <= 3'h1 & _s1_strb_wmask_0_T_4 > 4'h1;
  wire  s1_strb_wmask_2 = _s1_strb_T[2:0] <= 3'h2 & _s1_strb_wmask_0_T_4 > 4'h2;
  wire  s1_strb_wmask_3 = _s1_strb_T[2:0] <= 3'h3 & _s1_strb_wmask_0_T_4 > 4'h3;
  wire  s1_strb_wmask_4 = _s1_strb_T[2:0] <= 3'h4 & _s1_strb_wmask_0_T_4 > 4'h4;
  wire  s1_strb_wmask_5 = _s1_strb_T[2:0] <= 3'h5 & _s1_strb_wmask_0_T_4 > 4'h5;
  wire  s1_strb_wmask_6 = _s1_strb_T[2:0] <= 3'h6 & _s1_strb_wmask_0_T_4 > 4'h6;
  wire  s1_strb_wmask_7 = _s1_strb_wmask_0_T_4 > 4'h7;
  wire [7:0] s1_strb = {s1_strb_wmask_7,s1_strb_wmask_6,s1_strb_wmask_5,s1_strb_wmask_4,s1_strb_wmask_3,s1_strb_wmask_2,
    s1_strb_wmask_1,s1_strb_wmask_0};
  wire [63:0] dataWays_0_0 = io_dataArray_0_rdata[63:0];
  wire [63:0] dataWays_0_1 = io_dataArray_0_rdata[127:64];
  wire [63:0] dataWays_1_0 = io_dataArray_1_rdata[63:0];
  wire [63:0] dataWays_1_1 = io_dataArray_1_rdata[127:64];
  wire [63:0] dataWays_2_0 = io_dataArray_2_rdata[63:0];
  wire [63:0] dataWays_2_1 = io_dataArray_2_rdata[127:64];
  wire [63:0] dataWays_3_0 = io_dataArray_3_rdata[63:0];
  wire [63:0] dataWays_3_1 = io_dataArray_3_rdata[127:64];
  reg  s2_reg_valid;
  reg [63:0] s2_reg_wdata;
  reg  s2_reg_wen;
  reg [7:0] s2_reg_strb;
  reg  s2_reg_probe;
  wire  _noprobeStall_T = ~s2_reg_probe;
  wire  metaWays_3_valid = metaArray_3_io_r_data_valid;
  wire [21:0] metaWays_3_tag = metaArray_3_io_r_data_tag;
  wire  hitVec_3 = metaWays_3_valid & metaWays_3_tag == _s1_strb_T[31:10];
  wire  metaWays_2_valid = metaArray_2_io_r_data_valid;
  wire [21:0] metaWays_2_tag = metaArray_2_io_r_data_tag;
  wire  hitVec_2 = metaWays_2_valid & metaWays_2_tag == _s1_strb_T[31:10];
  wire  metaWays_1_valid = metaArray_1_io_r_data_valid;
  wire [21:0] metaWays_1_tag = metaArray_1_io_r_data_tag;
  wire  hitVec_1 = metaWays_1_valid & metaWays_1_tag == _s1_strb_T[31:10];
  wire  metaWays_0_valid = metaArray_0_io_r_data_valid;
  wire [21:0] metaWays_0_tag = metaArray_0_io_r_data_tag;
  wire  hitVec_0 = metaWays_0_valid & metaWays_0_tag == _s1_strb_T[31:10];
  wire [3:0] _s2_hit_T = {hitVec_3,hitVec_2,hitVec_1,hitVec_0};
  wire  s2_hit = |_s2_hit_T & s2_reg_valid;
  wire  s2_miss = s2_reg_valid & ~s2_hit;
  wire  noprobeStall = ~s2_reg_probe & s2_miss;
  wire  probeStall = s2_reg_probe & ~io_link_resp_valid;
  wire  s2_stall = s2_reg_valid & (noprobeStall | probeStall);
  wire  _GEN_3 = s1_valid & s1_wen;
  wire  _GEN_5 = s1_valid & s1_probe;
  wire [1:0] _GEN_12 = 6'h1 == req_addr_index ? regCount_1_0 : regCount_0_0;
  wire [1:0] _GEN_13 = 6'h2 == req_addr_index ? regCount_2_0 : _GEN_12;
  wire [1:0] _GEN_14 = 6'h3 == req_addr_index ? regCount_3_0 : _GEN_13;
  wire [1:0] _GEN_15 = 6'h4 == req_addr_index ? regCount_4_0 : _GEN_14;
  wire [1:0] _GEN_16 = 6'h5 == req_addr_index ? regCount_5_0 : _GEN_15;
  wire [1:0] _GEN_17 = 6'h6 == req_addr_index ? regCount_6_0 : _GEN_16;
  wire [1:0] _GEN_18 = 6'h7 == req_addr_index ? regCount_7_0 : _GEN_17;
  wire [1:0] _GEN_19 = 6'h8 == req_addr_index ? regCount_8_0 : _GEN_18;
  wire [1:0] _GEN_20 = 6'h9 == req_addr_index ? regCount_9_0 : _GEN_19;
  wire [1:0] _GEN_21 = 6'ha == req_addr_index ? regCount_10_0 : _GEN_20;
  wire [1:0] _GEN_22 = 6'hb == req_addr_index ? regCount_11_0 : _GEN_21;
  wire [1:0] _GEN_23 = 6'hc == req_addr_index ? regCount_12_0 : _GEN_22;
  wire [1:0] _GEN_24 = 6'hd == req_addr_index ? regCount_13_0 : _GEN_23;
  wire [1:0] _GEN_25 = 6'he == req_addr_index ? regCount_14_0 : _GEN_24;
  wire [1:0] _GEN_26 = 6'hf == req_addr_index ? regCount_15_0 : _GEN_25;
  wire [1:0] _GEN_27 = 6'h10 == req_addr_index ? regCount_16_0 : _GEN_26;
  wire [1:0] _GEN_28 = 6'h11 == req_addr_index ? regCount_17_0 : _GEN_27;
  wire [1:0] _GEN_29 = 6'h12 == req_addr_index ? regCount_18_0 : _GEN_28;
  wire [1:0] _GEN_30 = 6'h13 == req_addr_index ? regCount_19_0 : _GEN_29;
  wire [1:0] _GEN_31 = 6'h14 == req_addr_index ? regCount_20_0 : _GEN_30;
  wire [1:0] _GEN_32 = 6'h15 == req_addr_index ? regCount_21_0 : _GEN_31;
  wire [1:0] _GEN_33 = 6'h16 == req_addr_index ? regCount_22_0 : _GEN_32;
  wire [1:0] _GEN_34 = 6'h17 == req_addr_index ? regCount_23_0 : _GEN_33;
  wire [1:0] _GEN_35 = 6'h18 == req_addr_index ? regCount_24_0 : _GEN_34;
  wire [1:0] _GEN_36 = 6'h19 == req_addr_index ? regCount_25_0 : _GEN_35;
  wire [1:0] _GEN_37 = 6'h1a == req_addr_index ? regCount_26_0 : _GEN_36;
  wire [1:0] _GEN_38 = 6'h1b == req_addr_index ? regCount_27_0 : _GEN_37;
  wire [1:0] _GEN_39 = 6'h1c == req_addr_index ? regCount_28_0 : _GEN_38;
  wire [1:0] _GEN_40 = 6'h1d == req_addr_index ? regCount_29_0 : _GEN_39;
  wire [1:0] _GEN_41 = 6'h1e == req_addr_index ? regCount_30_0 : _GEN_40;
  wire [1:0] _GEN_42 = 6'h1f == req_addr_index ? regCount_31_0 : _GEN_41;
  wire [1:0] _GEN_43 = 6'h20 == req_addr_index ? regCount_32_0 : _GEN_42;
  wire [1:0] _GEN_44 = 6'h21 == req_addr_index ? regCount_33_0 : _GEN_43;
  wire [1:0] _GEN_45 = 6'h22 == req_addr_index ? regCount_34_0 : _GEN_44;
  wire [1:0] _GEN_46 = 6'h23 == req_addr_index ? regCount_35_0 : _GEN_45;
  wire [1:0] _GEN_47 = 6'h24 == req_addr_index ? regCount_36_0 : _GEN_46;
  wire [1:0] _GEN_48 = 6'h25 == req_addr_index ? regCount_37_0 : _GEN_47;
  wire [1:0] _GEN_49 = 6'h26 == req_addr_index ? regCount_38_0 : _GEN_48;
  wire [1:0] _GEN_50 = 6'h27 == req_addr_index ? regCount_39_0 : _GEN_49;
  wire [1:0] _GEN_51 = 6'h28 == req_addr_index ? regCount_40_0 : _GEN_50;
  wire [1:0] _GEN_52 = 6'h29 == req_addr_index ? regCount_41_0 : _GEN_51;
  wire [1:0] _GEN_53 = 6'h2a == req_addr_index ? regCount_42_0 : _GEN_52;
  wire [1:0] _GEN_54 = 6'h2b == req_addr_index ? regCount_43_0 : _GEN_53;
  wire [1:0] _GEN_55 = 6'h2c == req_addr_index ? regCount_44_0 : _GEN_54;
  wire [1:0] _GEN_56 = 6'h2d == req_addr_index ? regCount_45_0 : _GEN_55;
  wire [1:0] _GEN_57 = 6'h2e == req_addr_index ? regCount_46_0 : _GEN_56;
  wire [1:0] _GEN_58 = 6'h2f == req_addr_index ? regCount_47_0 : _GEN_57;
  wire [1:0] _GEN_59 = 6'h30 == req_addr_index ? regCount_48_0 : _GEN_58;
  wire [1:0] _GEN_60 = 6'h31 == req_addr_index ? regCount_49_0 : _GEN_59;
  wire [1:0] _GEN_61 = 6'h32 == req_addr_index ? regCount_50_0 : _GEN_60;
  wire [1:0] _GEN_62 = 6'h33 == req_addr_index ? regCount_51_0 : _GEN_61;
  wire [1:0] _GEN_63 = 6'h34 == req_addr_index ? regCount_52_0 : _GEN_62;
  wire [1:0] _GEN_64 = 6'h35 == req_addr_index ? regCount_53_0 : _GEN_63;
  wire [1:0] _GEN_65 = 6'h36 == req_addr_index ? regCount_54_0 : _GEN_64;
  wire [1:0] _GEN_66 = 6'h37 == req_addr_index ? regCount_55_0 : _GEN_65;
  wire [1:0] _GEN_67 = 6'h38 == req_addr_index ? regCount_56_0 : _GEN_66;
  wire [1:0] _GEN_68 = 6'h39 == req_addr_index ? regCount_57_0 : _GEN_67;
  wire [1:0] _GEN_69 = 6'h3a == req_addr_index ? regCount_58_0 : _GEN_68;
  wire [1:0] _GEN_70 = 6'h3b == req_addr_index ? regCount_59_0 : _GEN_69;
  wire [1:0] _GEN_71 = 6'h3c == req_addr_index ? regCount_60_0 : _GEN_70;
  wire [1:0] _GEN_72 = 6'h3d == req_addr_index ? regCount_61_0 : _GEN_71;
  wire [1:0] _GEN_73 = 6'h3e == req_addr_index ? regCount_62_0 : _GEN_72;
  wire [1:0] _GEN_74 = 6'h3f == req_addr_index ? regCount_63_0 : _GEN_73;
  wire [1:0] _GEN_76 = 6'h1 == req_addr_index ? regCount_1_1 : regCount_0_1;
  wire [1:0] _GEN_77 = 6'h2 == req_addr_index ? regCount_2_1 : _GEN_76;
  wire [1:0] _GEN_78 = 6'h3 == req_addr_index ? regCount_3_1 : _GEN_77;
  wire [1:0] _GEN_79 = 6'h4 == req_addr_index ? regCount_4_1 : _GEN_78;
  wire [1:0] _GEN_80 = 6'h5 == req_addr_index ? regCount_5_1 : _GEN_79;
  wire [1:0] _GEN_81 = 6'h6 == req_addr_index ? regCount_6_1 : _GEN_80;
  wire [1:0] _GEN_82 = 6'h7 == req_addr_index ? regCount_7_1 : _GEN_81;
  wire [1:0] _GEN_83 = 6'h8 == req_addr_index ? regCount_8_1 : _GEN_82;
  wire [1:0] _GEN_84 = 6'h9 == req_addr_index ? regCount_9_1 : _GEN_83;
  wire [1:0] _GEN_85 = 6'ha == req_addr_index ? regCount_10_1 : _GEN_84;
  wire [1:0] _GEN_86 = 6'hb == req_addr_index ? regCount_11_1 : _GEN_85;
  wire [1:0] _GEN_87 = 6'hc == req_addr_index ? regCount_12_1 : _GEN_86;
  wire [1:0] _GEN_88 = 6'hd == req_addr_index ? regCount_13_1 : _GEN_87;
  wire [1:0] _GEN_89 = 6'he == req_addr_index ? regCount_14_1 : _GEN_88;
  wire [1:0] _GEN_90 = 6'hf == req_addr_index ? regCount_15_1 : _GEN_89;
  wire [1:0] _GEN_91 = 6'h10 == req_addr_index ? regCount_16_1 : _GEN_90;
  wire [1:0] _GEN_92 = 6'h11 == req_addr_index ? regCount_17_1 : _GEN_91;
  wire [1:0] _GEN_93 = 6'h12 == req_addr_index ? regCount_18_1 : _GEN_92;
  wire [1:0] _GEN_94 = 6'h13 == req_addr_index ? regCount_19_1 : _GEN_93;
  wire [1:0] _GEN_95 = 6'h14 == req_addr_index ? regCount_20_1 : _GEN_94;
  wire [1:0] _GEN_96 = 6'h15 == req_addr_index ? regCount_21_1 : _GEN_95;
  wire [1:0] _GEN_97 = 6'h16 == req_addr_index ? regCount_22_1 : _GEN_96;
  wire [1:0] _GEN_98 = 6'h17 == req_addr_index ? regCount_23_1 : _GEN_97;
  wire [1:0] _GEN_99 = 6'h18 == req_addr_index ? regCount_24_1 : _GEN_98;
  wire [1:0] _GEN_100 = 6'h19 == req_addr_index ? regCount_25_1 : _GEN_99;
  wire [1:0] _GEN_101 = 6'h1a == req_addr_index ? regCount_26_1 : _GEN_100;
  wire [1:0] _GEN_102 = 6'h1b == req_addr_index ? regCount_27_1 : _GEN_101;
  wire [1:0] _GEN_103 = 6'h1c == req_addr_index ? regCount_28_1 : _GEN_102;
  wire [1:0] _GEN_104 = 6'h1d == req_addr_index ? regCount_29_1 : _GEN_103;
  wire [1:0] _GEN_105 = 6'h1e == req_addr_index ? regCount_30_1 : _GEN_104;
  wire [1:0] _GEN_106 = 6'h1f == req_addr_index ? regCount_31_1 : _GEN_105;
  wire [1:0] _GEN_107 = 6'h20 == req_addr_index ? regCount_32_1 : _GEN_106;
  wire [1:0] _GEN_108 = 6'h21 == req_addr_index ? regCount_33_1 : _GEN_107;
  wire [1:0] _GEN_109 = 6'h22 == req_addr_index ? regCount_34_1 : _GEN_108;
  wire [1:0] _GEN_110 = 6'h23 == req_addr_index ? regCount_35_1 : _GEN_109;
  wire [1:0] _GEN_111 = 6'h24 == req_addr_index ? regCount_36_1 : _GEN_110;
  wire [1:0] _GEN_112 = 6'h25 == req_addr_index ? regCount_37_1 : _GEN_111;
  wire [1:0] _GEN_113 = 6'h26 == req_addr_index ? regCount_38_1 : _GEN_112;
  wire [1:0] _GEN_114 = 6'h27 == req_addr_index ? regCount_39_1 : _GEN_113;
  wire [1:0] _GEN_115 = 6'h28 == req_addr_index ? regCount_40_1 : _GEN_114;
  wire [1:0] _GEN_116 = 6'h29 == req_addr_index ? regCount_41_1 : _GEN_115;
  wire [1:0] _GEN_117 = 6'h2a == req_addr_index ? regCount_42_1 : _GEN_116;
  wire [1:0] _GEN_118 = 6'h2b == req_addr_index ? regCount_43_1 : _GEN_117;
  wire [1:0] _GEN_119 = 6'h2c == req_addr_index ? regCount_44_1 : _GEN_118;
  wire [1:0] _GEN_120 = 6'h2d == req_addr_index ? regCount_45_1 : _GEN_119;
  wire [1:0] _GEN_121 = 6'h2e == req_addr_index ? regCount_46_1 : _GEN_120;
  wire [1:0] _GEN_122 = 6'h2f == req_addr_index ? regCount_47_1 : _GEN_121;
  wire [1:0] _GEN_123 = 6'h30 == req_addr_index ? regCount_48_1 : _GEN_122;
  wire [1:0] _GEN_124 = 6'h31 == req_addr_index ? regCount_49_1 : _GEN_123;
  wire [1:0] _GEN_125 = 6'h32 == req_addr_index ? regCount_50_1 : _GEN_124;
  wire [1:0] _GEN_126 = 6'h33 == req_addr_index ? regCount_51_1 : _GEN_125;
  wire [1:0] _GEN_127 = 6'h34 == req_addr_index ? regCount_52_1 : _GEN_126;
  wire [1:0] _GEN_128 = 6'h35 == req_addr_index ? regCount_53_1 : _GEN_127;
  wire [1:0] _GEN_129 = 6'h36 == req_addr_index ? regCount_54_1 : _GEN_128;
  wire [1:0] _GEN_130 = 6'h37 == req_addr_index ? regCount_55_1 : _GEN_129;
  wire [1:0] _GEN_131 = 6'h38 == req_addr_index ? regCount_56_1 : _GEN_130;
  wire [1:0] _GEN_132 = 6'h39 == req_addr_index ? regCount_57_1 : _GEN_131;
  wire [1:0] _GEN_133 = 6'h3a == req_addr_index ? regCount_58_1 : _GEN_132;
  wire [1:0] _GEN_134 = 6'h3b == req_addr_index ? regCount_59_1 : _GEN_133;
  wire [1:0] _GEN_135 = 6'h3c == req_addr_index ? regCount_60_1 : _GEN_134;
  wire [1:0] _GEN_136 = 6'h3d == req_addr_index ? regCount_61_1 : _GEN_135;
  wire [1:0] _GEN_137 = 6'h3e == req_addr_index ? regCount_62_1 : _GEN_136;
  wire [1:0] _GEN_138 = 6'h3f == req_addr_index ? regCount_63_1 : _GEN_137;
  wire [1:0] _GEN_140 = 6'h1 == req_addr_index ? regCount_1_2 : regCount_0_2;
  wire [1:0] _GEN_141 = 6'h2 == req_addr_index ? regCount_2_2 : _GEN_140;
  wire [1:0] _GEN_142 = 6'h3 == req_addr_index ? regCount_3_2 : _GEN_141;
  wire [1:0] _GEN_143 = 6'h4 == req_addr_index ? regCount_4_2 : _GEN_142;
  wire [1:0] _GEN_144 = 6'h5 == req_addr_index ? regCount_5_2 : _GEN_143;
  wire [1:0] _GEN_145 = 6'h6 == req_addr_index ? regCount_6_2 : _GEN_144;
  wire [1:0] _GEN_146 = 6'h7 == req_addr_index ? regCount_7_2 : _GEN_145;
  wire [1:0] _GEN_147 = 6'h8 == req_addr_index ? regCount_8_2 : _GEN_146;
  wire [1:0] _GEN_148 = 6'h9 == req_addr_index ? regCount_9_2 : _GEN_147;
  wire [1:0] _GEN_149 = 6'ha == req_addr_index ? regCount_10_2 : _GEN_148;
  wire [1:0] _GEN_150 = 6'hb == req_addr_index ? regCount_11_2 : _GEN_149;
  wire [1:0] _GEN_151 = 6'hc == req_addr_index ? regCount_12_2 : _GEN_150;
  wire [1:0] _GEN_152 = 6'hd == req_addr_index ? regCount_13_2 : _GEN_151;
  wire [1:0] _GEN_153 = 6'he == req_addr_index ? regCount_14_2 : _GEN_152;
  wire [1:0] _GEN_154 = 6'hf == req_addr_index ? regCount_15_2 : _GEN_153;
  wire [1:0] _GEN_155 = 6'h10 == req_addr_index ? regCount_16_2 : _GEN_154;
  wire [1:0] _GEN_156 = 6'h11 == req_addr_index ? regCount_17_2 : _GEN_155;
  wire [1:0] _GEN_157 = 6'h12 == req_addr_index ? regCount_18_2 : _GEN_156;
  wire [1:0] _GEN_158 = 6'h13 == req_addr_index ? regCount_19_2 : _GEN_157;
  wire [1:0] _GEN_159 = 6'h14 == req_addr_index ? regCount_20_2 : _GEN_158;
  wire [1:0] _GEN_160 = 6'h15 == req_addr_index ? regCount_21_2 : _GEN_159;
  wire [1:0] _GEN_161 = 6'h16 == req_addr_index ? regCount_22_2 : _GEN_160;
  wire [1:0] _GEN_162 = 6'h17 == req_addr_index ? regCount_23_2 : _GEN_161;
  wire [1:0] _GEN_163 = 6'h18 == req_addr_index ? regCount_24_2 : _GEN_162;
  wire [1:0] _GEN_164 = 6'h19 == req_addr_index ? regCount_25_2 : _GEN_163;
  wire [1:0] _GEN_165 = 6'h1a == req_addr_index ? regCount_26_2 : _GEN_164;
  wire [1:0] _GEN_166 = 6'h1b == req_addr_index ? regCount_27_2 : _GEN_165;
  wire [1:0] _GEN_167 = 6'h1c == req_addr_index ? regCount_28_2 : _GEN_166;
  wire [1:0] _GEN_168 = 6'h1d == req_addr_index ? regCount_29_2 : _GEN_167;
  wire [1:0] _GEN_169 = 6'h1e == req_addr_index ? regCount_30_2 : _GEN_168;
  wire [1:0] _GEN_170 = 6'h1f == req_addr_index ? regCount_31_2 : _GEN_169;
  wire [1:0] _GEN_171 = 6'h20 == req_addr_index ? regCount_32_2 : _GEN_170;
  wire [1:0] _GEN_172 = 6'h21 == req_addr_index ? regCount_33_2 : _GEN_171;
  wire [1:0] _GEN_173 = 6'h22 == req_addr_index ? regCount_34_2 : _GEN_172;
  wire [1:0] _GEN_174 = 6'h23 == req_addr_index ? regCount_35_2 : _GEN_173;
  wire [1:0] _GEN_175 = 6'h24 == req_addr_index ? regCount_36_2 : _GEN_174;
  wire [1:0] _GEN_176 = 6'h25 == req_addr_index ? regCount_37_2 : _GEN_175;
  wire [1:0] _GEN_177 = 6'h26 == req_addr_index ? regCount_38_2 : _GEN_176;
  wire [1:0] _GEN_178 = 6'h27 == req_addr_index ? regCount_39_2 : _GEN_177;
  wire [1:0] _GEN_179 = 6'h28 == req_addr_index ? regCount_40_2 : _GEN_178;
  wire [1:0] _GEN_180 = 6'h29 == req_addr_index ? regCount_41_2 : _GEN_179;
  wire [1:0] _GEN_181 = 6'h2a == req_addr_index ? regCount_42_2 : _GEN_180;
  wire [1:0] _GEN_182 = 6'h2b == req_addr_index ? regCount_43_2 : _GEN_181;
  wire [1:0] _GEN_183 = 6'h2c == req_addr_index ? regCount_44_2 : _GEN_182;
  wire [1:0] _GEN_184 = 6'h2d == req_addr_index ? regCount_45_2 : _GEN_183;
  wire [1:0] _GEN_185 = 6'h2e == req_addr_index ? regCount_46_2 : _GEN_184;
  wire [1:0] _GEN_186 = 6'h2f == req_addr_index ? regCount_47_2 : _GEN_185;
  wire [1:0] _GEN_187 = 6'h30 == req_addr_index ? regCount_48_2 : _GEN_186;
  wire [1:0] _GEN_188 = 6'h31 == req_addr_index ? regCount_49_2 : _GEN_187;
  wire [1:0] _GEN_189 = 6'h32 == req_addr_index ? regCount_50_2 : _GEN_188;
  wire [1:0] _GEN_190 = 6'h33 == req_addr_index ? regCount_51_2 : _GEN_189;
  wire [1:0] _GEN_191 = 6'h34 == req_addr_index ? regCount_52_2 : _GEN_190;
  wire [1:0] _GEN_192 = 6'h35 == req_addr_index ? regCount_53_2 : _GEN_191;
  wire [1:0] _GEN_193 = 6'h36 == req_addr_index ? regCount_54_2 : _GEN_192;
  wire [1:0] _GEN_194 = 6'h37 == req_addr_index ? regCount_55_2 : _GEN_193;
  wire [1:0] _GEN_195 = 6'h38 == req_addr_index ? regCount_56_2 : _GEN_194;
  wire [1:0] _GEN_196 = 6'h39 == req_addr_index ? regCount_57_2 : _GEN_195;
  wire [1:0] _GEN_197 = 6'h3a == req_addr_index ? regCount_58_2 : _GEN_196;
  wire [1:0] _GEN_198 = 6'h3b == req_addr_index ? regCount_59_2 : _GEN_197;
  wire [1:0] _GEN_199 = 6'h3c == req_addr_index ? regCount_60_2 : _GEN_198;
  wire [1:0] _GEN_200 = 6'h3d == req_addr_index ? regCount_61_2 : _GEN_199;
  wire [1:0] _GEN_201 = 6'h3e == req_addr_index ? regCount_62_2 : _GEN_200;
  wire [1:0] _GEN_202 = 6'h3f == req_addr_index ? regCount_63_2 : _GEN_201;
  wire [1:0] _GEN_204 = 6'h1 == req_addr_index ? regCount_1_3 : regCount_0_3;
  wire [1:0] _GEN_205 = 6'h2 == req_addr_index ? regCount_2_3 : _GEN_204;
  wire [1:0] _GEN_206 = 6'h3 == req_addr_index ? regCount_3_3 : _GEN_205;
  wire [1:0] _GEN_207 = 6'h4 == req_addr_index ? regCount_4_3 : _GEN_206;
  wire [1:0] _GEN_208 = 6'h5 == req_addr_index ? regCount_5_3 : _GEN_207;
  wire [1:0] _GEN_209 = 6'h6 == req_addr_index ? regCount_6_3 : _GEN_208;
  wire [1:0] _GEN_210 = 6'h7 == req_addr_index ? regCount_7_3 : _GEN_209;
  wire [1:0] _GEN_211 = 6'h8 == req_addr_index ? regCount_8_3 : _GEN_210;
  wire [1:0] _GEN_212 = 6'h9 == req_addr_index ? regCount_9_3 : _GEN_211;
  wire [1:0] _GEN_213 = 6'ha == req_addr_index ? regCount_10_3 : _GEN_212;
  wire [1:0] _GEN_214 = 6'hb == req_addr_index ? regCount_11_3 : _GEN_213;
  wire [1:0] _GEN_215 = 6'hc == req_addr_index ? regCount_12_3 : _GEN_214;
  wire [1:0] _GEN_216 = 6'hd == req_addr_index ? regCount_13_3 : _GEN_215;
  wire [1:0] _GEN_217 = 6'he == req_addr_index ? regCount_14_3 : _GEN_216;
  wire [1:0] _GEN_218 = 6'hf == req_addr_index ? regCount_15_3 : _GEN_217;
  wire [1:0] _GEN_219 = 6'h10 == req_addr_index ? regCount_16_3 : _GEN_218;
  wire [1:0] _GEN_220 = 6'h11 == req_addr_index ? regCount_17_3 : _GEN_219;
  wire [1:0] _GEN_221 = 6'h12 == req_addr_index ? regCount_18_3 : _GEN_220;
  wire [1:0] _GEN_222 = 6'h13 == req_addr_index ? regCount_19_3 : _GEN_221;
  wire [1:0] _GEN_223 = 6'h14 == req_addr_index ? regCount_20_3 : _GEN_222;
  wire [1:0] _GEN_224 = 6'h15 == req_addr_index ? regCount_21_3 : _GEN_223;
  wire [1:0] _GEN_225 = 6'h16 == req_addr_index ? regCount_22_3 : _GEN_224;
  wire [1:0] _GEN_226 = 6'h17 == req_addr_index ? regCount_23_3 : _GEN_225;
  wire [1:0] _GEN_227 = 6'h18 == req_addr_index ? regCount_24_3 : _GEN_226;
  wire [1:0] _GEN_228 = 6'h19 == req_addr_index ? regCount_25_3 : _GEN_227;
  wire [1:0] _GEN_229 = 6'h1a == req_addr_index ? regCount_26_3 : _GEN_228;
  wire [1:0] _GEN_230 = 6'h1b == req_addr_index ? regCount_27_3 : _GEN_229;
  wire [1:0] _GEN_231 = 6'h1c == req_addr_index ? regCount_28_3 : _GEN_230;
  wire [1:0] _GEN_232 = 6'h1d == req_addr_index ? regCount_29_3 : _GEN_231;
  wire [1:0] _GEN_233 = 6'h1e == req_addr_index ? regCount_30_3 : _GEN_232;
  wire [1:0] _GEN_234 = 6'h1f == req_addr_index ? regCount_31_3 : _GEN_233;
  wire [1:0] _GEN_235 = 6'h20 == req_addr_index ? regCount_32_3 : _GEN_234;
  wire [1:0] _GEN_236 = 6'h21 == req_addr_index ? regCount_33_3 : _GEN_235;
  wire [1:0] _GEN_237 = 6'h22 == req_addr_index ? regCount_34_3 : _GEN_236;
  wire [1:0] _GEN_238 = 6'h23 == req_addr_index ? regCount_35_3 : _GEN_237;
  wire [1:0] _GEN_239 = 6'h24 == req_addr_index ? regCount_36_3 : _GEN_238;
  wire [1:0] _GEN_240 = 6'h25 == req_addr_index ? regCount_37_3 : _GEN_239;
  wire [1:0] _GEN_241 = 6'h26 == req_addr_index ? regCount_38_3 : _GEN_240;
  wire [1:0] _GEN_242 = 6'h27 == req_addr_index ? regCount_39_3 : _GEN_241;
  wire [1:0] _GEN_243 = 6'h28 == req_addr_index ? regCount_40_3 : _GEN_242;
  wire [1:0] _GEN_244 = 6'h29 == req_addr_index ? regCount_41_3 : _GEN_243;
  wire [1:0] _GEN_245 = 6'h2a == req_addr_index ? regCount_42_3 : _GEN_244;
  wire [1:0] _GEN_246 = 6'h2b == req_addr_index ? regCount_43_3 : _GEN_245;
  wire [1:0] _GEN_247 = 6'h2c == req_addr_index ? regCount_44_3 : _GEN_246;
  wire [1:0] _GEN_248 = 6'h2d == req_addr_index ? regCount_45_3 : _GEN_247;
  wire [1:0] _GEN_249 = 6'h2e == req_addr_index ? regCount_46_3 : _GEN_248;
  wire [1:0] _GEN_250 = 6'h2f == req_addr_index ? regCount_47_3 : _GEN_249;
  wire [1:0] _GEN_251 = 6'h30 == req_addr_index ? regCount_48_3 : _GEN_250;
  wire [1:0] _GEN_252 = 6'h31 == req_addr_index ? regCount_49_3 : _GEN_251;
  wire [1:0] _GEN_253 = 6'h32 == req_addr_index ? regCount_50_3 : _GEN_252;
  wire [1:0] _GEN_254 = 6'h33 == req_addr_index ? regCount_51_3 : _GEN_253;
  wire [1:0] _GEN_255 = 6'h34 == req_addr_index ? regCount_52_3 : _GEN_254;
  wire [1:0] _GEN_256 = 6'h35 == req_addr_index ? regCount_53_3 : _GEN_255;
  wire [1:0] _GEN_257 = 6'h36 == req_addr_index ? regCount_54_3 : _GEN_256;
  wire [1:0] _GEN_258 = 6'h37 == req_addr_index ? regCount_55_3 : _GEN_257;
  wire [1:0] _GEN_259 = 6'h38 == req_addr_index ? regCount_56_3 : _GEN_258;
  wire [1:0] _GEN_260 = 6'h39 == req_addr_index ? regCount_57_3 : _GEN_259;
  wire [1:0] _GEN_261 = 6'h3a == req_addr_index ? regCount_58_3 : _GEN_260;
  wire [1:0] _GEN_262 = 6'h3b == req_addr_index ? regCount_59_3 : _GEN_261;
  wire [1:0] _GEN_263 = 6'h3c == req_addr_index ? regCount_60_3 : _GEN_262;
  wire [1:0] _GEN_264 = 6'h3d == req_addr_index ? regCount_61_3 : _GEN_263;
  wire [1:0] _GEN_265 = 6'h3e == req_addr_index ? regCount_62_3 : _GEN_264;
  wire [1:0] _GEN_266 = 6'h3f == req_addr_index ? regCount_63_3 : _GEN_265;
  wire [1:0] s2_idxWayHit_hi_1 = _s2_hit_T[3:2];
  wire [1:0] s2_idxWayHit_lo_1 = _s2_hit_T[1:0];
  wire  _s2_idxWayHit_T_1 = |s2_idxWayHit_hi_1;
  wire [1:0] _s2_idxWayHit_T_2 = s2_idxWayHit_hi_1 | s2_idxWayHit_lo_1;
  wire [1:0] s2_idxWayHit = {_s2_idxWayHit_T_1,_s2_idxWayHit_T_2[1]};
  wire [1:0] s2_wordsMask = 2'h1 << req_addr_wordOffest;
  wire [63:0] _s2_dataBlockHit_T = hitVec_0 ? dataWays_0_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_1 = hitVec_1 ? dataWays_1_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_2 = hitVec_2 ? dataWays_2_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_3 = hitVec_3 ? dataWays_3_0 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_4 = _s2_dataBlockHit_T | _s2_dataBlockHit_T_1;
  wire [63:0] _s2_dataBlockHit_T_5 = _s2_dataBlockHit_T_4 | _s2_dataBlockHit_T_2;
  wire [63:0] s2_dataBlockHit_0 = _s2_dataBlockHit_T_5 | _s2_dataBlockHit_T_3;
  wire [63:0] _s2_dataBlockHit_T_7 = hitVec_0 ? dataWays_0_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_8 = hitVec_1 ? dataWays_1_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_9 = hitVec_2 ? dataWays_2_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_10 = hitVec_3 ? dataWays_3_1 : 64'h0;
  wire [63:0] _s2_dataBlockHit_T_11 = _s2_dataBlockHit_T_7 | _s2_dataBlockHit_T_8;
  wire [63:0] _s2_dataBlockHit_T_12 = _s2_dataBlockHit_T_11 | _s2_dataBlockHit_T_9;
  wire [63:0] s2_dataBlockHit_1 = _s2_dataBlockHit_T_12 | _s2_dataBlockHit_T_10;
  wire [63:0] _s2_hitWord_T_2 = s2_wordsMask[0] ? s2_dataBlockHit_0 : 64'h0;
  wire [63:0] _s2_hitWord_T_3 = s2_wordsMask[1] ? s2_dataBlockHit_1 : 64'h0;
  wire [63:0] rWord = _s2_hitWord_T_2 | _s2_hitWord_T_3;
  wire [7:0] _wmask_T_9 = s2_reg_strb[0] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_11 = s2_reg_strb[1] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_13 = s2_reg_strb[2] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_15 = s2_reg_strb[3] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_17 = s2_reg_strb[4] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_19 = s2_reg_strb[5] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_21 = s2_reg_strb[6] ? 8'hff : 8'h0;
  wire [7:0] _wmask_T_23 = s2_reg_strb[7] ? 8'hff : 8'h0;
  wire [63:0] wmask = {_wmask_T_23,_wmask_T_21,_wmask_T_19,_wmask_T_17,_wmask_T_15,_wmask_T_13,_wmask_T_11,_wmask_T_9};
  wire [63:0] _wordAfterWrite_T = s2_reg_wdata & wmask;
  wire [63:0] _wordAfterWrite_T_1 = ~wmask;
  wire [63:0] _wordAfterWrite_T_2 = rWord & _wordAfterWrite_T_1;
  wire [63:0] wordAfterWrite = _wordAfterWrite_T | _wordAfterWrite_T_2;
  wire [127:0] _s2_writeBlock_T = {s2_dataBlockHit_1,s2_dataBlockHit_0};
  wire [63:0] _GEN_267 = ~req_addr_wordOffest ? wordAfterWrite : _s2_writeBlock_T[63:0];
  wire [63:0] _GEN_268 = req_addr_wordOffest ? wordAfterWrite : _s2_writeBlock_T[127:64];
  wire [63:0] s2_writeBlock_0 = s2_reg_wen ? _GEN_267 : _s2_writeBlock_T[63:0];
  wire [63:0] s2_writeBlock_1 = s2_reg_wen ? _GEN_268 : _s2_writeBlock_T[127:64];
  wire [1:0] selectWay = selTree_io_outIdx;
  wire  metaWays_0_needFlush = metaArray_0_io_r_data_needFlush;
  wire  metaWays_1_needFlush = metaArray_1_io_r_data_needFlush;
  wire  _GEN_273 = 2'h1 == selectWay ? metaWays_1_needFlush : metaWays_0_needFlush;
  wire  metaWays_2_needFlush = metaArray_2_io_r_data_needFlush;
  wire  _GEN_274 = 2'h2 == selectWay ? metaWays_2_needFlush : _GEN_273;
  wire  metaWays_3_needFlush = metaArray_3_io_r_data_needFlush;
  wire  _GEN_275 = 2'h3 == selectWay ? metaWays_3_needFlush : _GEN_274;
  wire [2:0] _GEN_276 = _GEN_275 ? 3'h4 : 3'h2;
  wire [2:0] _GEN_277 = io_in_resp_valid ? 3'h0 : c_state;
  wire [2:0] _GEN_278 = s2_miss ? _GEN_276 : _GEN_277;
  wire [2:0] _GEN_279 = io_link_resp_valid ? 3'h0 : c_state;
  wire [2:0] _GEN_280 = io_link_resp_valid ? 3'h6 : c_state;
  wire [2:0] _GEN_281 = s2_miss ? _GEN_279 : _GEN_280;
  wire  _T_18 = io_out_req_ready & io_out_req_valid;
  wire [2:0] _GEN_283 = _T_18 ? 3'h3 : c_state;
  wire  _T_20 = io_out_resp_ready & io_out_resp_valid;
  wire [2:0] _GEN_284 = _T_20 ? 3'h7 : c_state;
  wire [2:0] _GEN_285 = _T_18 ? 3'h5 : c_state;
  wire [2:0] _GEN_286 = _T_20 ? 3'h2 : c_state;
  wire [2:0] _GEN_289 = 3'h7 == c_state ? _GEN_277 : c_state;
  wire [2:0] _GEN_290 = 3'h6 == c_state ? _GEN_279 : _GEN_289;
  wire [2:0] _GEN_291 = 3'h5 == c_state ? _GEN_286 : _GEN_290;
  wire [2:0] _GEN_292 = 3'h4 == c_state ? _GEN_285 : _GEN_291;
  wire [2:0] _GEN_293 = 3'h3 == c_state ? _GEN_284 : _GEN_292;
  wire  memRespUpdate = c_state == 3'h3 & _T_20;
  wire  _hitUpdate_T = c_state == 3'h1;
  wire  hitUpdate = c_state == 3'h1 & s2_hit;
  wire [21:0] _GEN_298 = 2'h1 == s2_idxWayHit ? metaWays_1_tag : metaWays_0_tag;
  wire [21:0] _GEN_299 = 2'h2 == s2_idxWayHit ? metaWays_2_tag : _GEN_298;
  wire [21:0] newMetaDirty_tag = 2'h3 == s2_idxWayHit ? metaWays_3_tag : _GEN_299;
  wire  _GEN_302 = 2'h1 == s2_idxWayHit ? metaWays_1_valid : metaWays_0_valid;
  wire  _GEN_303 = 2'h2 == s2_idxWayHit ? metaWays_2_valid : _GEN_302;
  wire  newMetaDirty_valid = 2'h3 == s2_idxWayHit ? metaWays_3_valid : _GEN_303;
  wire  _GEN_306 = 2'h1 == s2_idxWayHit ? metaWays_1_needFlush : metaWays_0_needFlush;
  wire  _GEN_307 = 2'h2 == s2_idxWayHit ? metaWays_2_needFlush : _GEN_306;
  wire  _GEN_308 = 2'h3 == s2_idxWayHit ? metaWays_3_needFlush : _GEN_307;
  wire  newMetaDirty_needFlush = s2_reg_wen | _GEN_308;
  wire  _cacheUpdate_T_2 = _hitUpdate_T | c_state == 3'h7;
  wire  cacheUpdate = memRespUpdate | (_hitUpdate_T | c_state == 3'h7) & s2_reg_wen & s2_hit;
  wire [1:0] wayWrite = memRespUpdate ? selectWay : s2_idxWayHit;
  wire  _metaArray_0_io_w_wen_T_1 = cacheUpdate & 2'h0 == wayWrite;
  wire  _metaArray_1_io_w_wen_T_1 = cacheUpdate & 2'h1 == wayWrite;
  wire  _metaArray_2_io_w_wen_T_1 = cacheUpdate & 2'h2 == wayWrite;
  wire  _metaArray_3_io_w_wen_T_1 = cacheUpdate & 2'h3 == wayWrite;
  wire [63:0] dataRefill_0 = io_out_resp_bits_rdata[63:0];
  wire [63:0] dataRefill_1 = io_out_resp_bits_rdata[127:64];
  wire [63:0] newBlock_0 = memRespUpdate ? dataRefill_0 : s2_writeBlock_0;
  wire [63:0] newBlock_1 = memRespUpdate ? dataRefill_1 : s2_writeBlock_1;
  wire [127:0] _io_dataArray_0_wdata_T_1 = {newBlock_1,newBlock_0};
  wire [1:0] _GEN_311 = 6'h0 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_0_1 : regCount_0_0;
  wire [1:0] _GEN_312 = 6'h0 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_0_2 : _GEN_311;
  wire [1:0] _GEN_313 = 6'h0 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_0_3 : _GEN_312;
  wire [1:0] _GEN_314 = 6'h1 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_1_0 : _GEN_313;
  wire [1:0] _GEN_315 = 6'h1 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_1_1 : _GEN_314;
  wire [1:0] _GEN_316 = 6'h1 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_1_2 : _GEN_315;
  wire [1:0] _GEN_317 = 6'h1 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_1_3 : _GEN_316;
  wire [1:0] _GEN_318 = 6'h2 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_2_0 : _GEN_317;
  wire [1:0] _GEN_319 = 6'h2 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_2_1 : _GEN_318;
  wire [1:0] _GEN_320 = 6'h2 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_2_2 : _GEN_319;
  wire [1:0] _GEN_321 = 6'h2 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_2_3 : _GEN_320;
  wire [1:0] _GEN_322 = 6'h3 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_3_0 : _GEN_321;
  wire [1:0] _GEN_323 = 6'h3 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_3_1 : _GEN_322;
  wire [1:0] _GEN_324 = 6'h3 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_3_2 : _GEN_323;
  wire [1:0] _GEN_325 = 6'h3 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_3_3 : _GEN_324;
  wire [1:0] _GEN_326 = 6'h4 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_4_0 : _GEN_325;
  wire [1:0] _GEN_327 = 6'h4 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_4_1 : _GEN_326;
  wire [1:0] _GEN_328 = 6'h4 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_4_2 : _GEN_327;
  wire [1:0] _GEN_329 = 6'h4 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_4_3 : _GEN_328;
  wire [1:0] _GEN_330 = 6'h5 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_5_0 : _GEN_329;
  wire [1:0] _GEN_331 = 6'h5 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_5_1 : _GEN_330;
  wire [1:0] _GEN_332 = 6'h5 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_5_2 : _GEN_331;
  wire [1:0] _GEN_333 = 6'h5 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_5_3 : _GEN_332;
  wire [1:0] _GEN_334 = 6'h6 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_6_0 : _GEN_333;
  wire [1:0] _GEN_335 = 6'h6 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_6_1 : _GEN_334;
  wire [1:0] _GEN_336 = 6'h6 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_6_2 : _GEN_335;
  wire [1:0] _GEN_337 = 6'h6 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_6_3 : _GEN_336;
  wire [1:0] _GEN_338 = 6'h7 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_7_0 : _GEN_337;
  wire [1:0] _GEN_339 = 6'h7 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_7_1 : _GEN_338;
  wire [1:0] _GEN_340 = 6'h7 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_7_2 : _GEN_339;
  wire [1:0] _GEN_341 = 6'h7 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_7_3 : _GEN_340;
  wire [1:0] _GEN_342 = 6'h8 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_8_0 : _GEN_341;
  wire [1:0] _GEN_343 = 6'h8 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_8_1 : _GEN_342;
  wire [1:0] _GEN_344 = 6'h8 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_8_2 : _GEN_343;
  wire [1:0] _GEN_345 = 6'h8 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_8_3 : _GEN_344;
  wire [1:0] _GEN_346 = 6'h9 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_9_0 : _GEN_345;
  wire [1:0] _GEN_347 = 6'h9 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_9_1 : _GEN_346;
  wire [1:0] _GEN_348 = 6'h9 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_9_2 : _GEN_347;
  wire [1:0] _GEN_349 = 6'h9 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_9_3 : _GEN_348;
  wire [1:0] _GEN_350 = 6'ha == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_10_0 : _GEN_349;
  wire [1:0] _GEN_351 = 6'ha == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_10_1 : _GEN_350;
  wire [1:0] _GEN_352 = 6'ha == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_10_2 : _GEN_351;
  wire [1:0] _GEN_353 = 6'ha == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_10_3 : _GEN_352;
  wire [1:0] _GEN_354 = 6'hb == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_11_0 : _GEN_353;
  wire [1:0] _GEN_355 = 6'hb == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_11_1 : _GEN_354;
  wire [1:0] _GEN_356 = 6'hb == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_11_2 : _GEN_355;
  wire [1:0] _GEN_357 = 6'hb == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_11_3 : _GEN_356;
  wire [1:0] _GEN_358 = 6'hc == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_12_0 : _GEN_357;
  wire [1:0] _GEN_359 = 6'hc == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_12_1 : _GEN_358;
  wire [1:0] _GEN_360 = 6'hc == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_12_2 : _GEN_359;
  wire [1:0] _GEN_361 = 6'hc == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_12_3 : _GEN_360;
  wire [1:0] _GEN_362 = 6'hd == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_13_0 : _GEN_361;
  wire [1:0] _GEN_363 = 6'hd == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_13_1 : _GEN_362;
  wire [1:0] _GEN_364 = 6'hd == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_13_2 : _GEN_363;
  wire [1:0] _GEN_365 = 6'hd == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_13_3 : _GEN_364;
  wire [1:0] _GEN_366 = 6'he == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_14_0 : _GEN_365;
  wire [1:0] _GEN_367 = 6'he == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_14_1 : _GEN_366;
  wire [1:0] _GEN_368 = 6'he == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_14_2 : _GEN_367;
  wire [1:0] _GEN_369 = 6'he == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_14_3 : _GEN_368;
  wire [1:0] _GEN_370 = 6'hf == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_15_0 : _GEN_369;
  wire [1:0] _GEN_371 = 6'hf == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_15_1 : _GEN_370;
  wire [1:0] _GEN_372 = 6'hf == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_15_2 : _GEN_371;
  wire [1:0] _GEN_373 = 6'hf == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_15_3 : _GEN_372;
  wire [1:0] _GEN_374 = 6'h10 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_16_0 : _GEN_373;
  wire [1:0] _GEN_375 = 6'h10 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_16_1 : _GEN_374;
  wire [1:0] _GEN_376 = 6'h10 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_16_2 : _GEN_375;
  wire [1:0] _GEN_377 = 6'h10 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_16_3 : _GEN_376;
  wire [1:0] _GEN_378 = 6'h11 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_17_0 : _GEN_377;
  wire [1:0] _GEN_379 = 6'h11 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_17_1 : _GEN_378;
  wire [1:0] _GEN_380 = 6'h11 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_17_2 : _GEN_379;
  wire [1:0] _GEN_381 = 6'h11 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_17_3 : _GEN_380;
  wire [1:0] _GEN_382 = 6'h12 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_18_0 : _GEN_381;
  wire [1:0] _GEN_383 = 6'h12 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_18_1 : _GEN_382;
  wire [1:0] _GEN_384 = 6'h12 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_18_2 : _GEN_383;
  wire [1:0] _GEN_385 = 6'h12 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_18_3 : _GEN_384;
  wire [1:0] _GEN_386 = 6'h13 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_19_0 : _GEN_385;
  wire [1:0] _GEN_387 = 6'h13 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_19_1 : _GEN_386;
  wire [1:0] _GEN_388 = 6'h13 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_19_2 : _GEN_387;
  wire [1:0] _GEN_389 = 6'h13 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_19_3 : _GEN_388;
  wire [1:0] _GEN_390 = 6'h14 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_20_0 : _GEN_389;
  wire [1:0] _GEN_391 = 6'h14 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_20_1 : _GEN_390;
  wire [1:0] _GEN_392 = 6'h14 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_20_2 : _GEN_391;
  wire [1:0] _GEN_393 = 6'h14 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_20_3 : _GEN_392;
  wire [1:0] _GEN_394 = 6'h15 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_21_0 : _GEN_393;
  wire [1:0] _GEN_395 = 6'h15 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_21_1 : _GEN_394;
  wire [1:0] _GEN_396 = 6'h15 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_21_2 : _GEN_395;
  wire [1:0] _GEN_397 = 6'h15 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_21_3 : _GEN_396;
  wire [1:0] _GEN_398 = 6'h16 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_22_0 : _GEN_397;
  wire [1:0] _GEN_399 = 6'h16 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_22_1 : _GEN_398;
  wire [1:0] _GEN_400 = 6'h16 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_22_2 : _GEN_399;
  wire [1:0] _GEN_401 = 6'h16 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_22_3 : _GEN_400;
  wire [1:0] _GEN_402 = 6'h17 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_23_0 : _GEN_401;
  wire [1:0] _GEN_403 = 6'h17 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_23_1 : _GEN_402;
  wire [1:0] _GEN_404 = 6'h17 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_23_2 : _GEN_403;
  wire [1:0] _GEN_405 = 6'h17 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_23_3 : _GEN_404;
  wire [1:0] _GEN_406 = 6'h18 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_24_0 : _GEN_405;
  wire [1:0] _GEN_407 = 6'h18 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_24_1 : _GEN_406;
  wire [1:0] _GEN_408 = 6'h18 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_24_2 : _GEN_407;
  wire [1:0] _GEN_409 = 6'h18 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_24_3 : _GEN_408;
  wire [1:0] _GEN_410 = 6'h19 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_25_0 : _GEN_409;
  wire [1:0] _GEN_411 = 6'h19 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_25_1 : _GEN_410;
  wire [1:0] _GEN_412 = 6'h19 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_25_2 : _GEN_411;
  wire [1:0] _GEN_413 = 6'h19 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_25_3 : _GEN_412;
  wire [1:0] _GEN_414 = 6'h1a == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_26_0 : _GEN_413;
  wire [1:0] _GEN_415 = 6'h1a == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_26_1 : _GEN_414;
  wire [1:0] _GEN_416 = 6'h1a == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_26_2 : _GEN_415;
  wire [1:0] _GEN_417 = 6'h1a == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_26_3 : _GEN_416;
  wire [1:0] _GEN_418 = 6'h1b == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_27_0 : _GEN_417;
  wire [1:0] _GEN_419 = 6'h1b == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_27_1 : _GEN_418;
  wire [1:0] _GEN_420 = 6'h1b == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_27_2 : _GEN_419;
  wire [1:0] _GEN_421 = 6'h1b == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_27_3 : _GEN_420;
  wire [1:0] _GEN_422 = 6'h1c == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_28_0 : _GEN_421;
  wire [1:0] _GEN_423 = 6'h1c == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_28_1 : _GEN_422;
  wire [1:0] _GEN_424 = 6'h1c == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_28_2 : _GEN_423;
  wire [1:0] _GEN_425 = 6'h1c == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_28_3 : _GEN_424;
  wire [1:0] _GEN_426 = 6'h1d == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_29_0 : _GEN_425;
  wire [1:0] _GEN_427 = 6'h1d == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_29_1 : _GEN_426;
  wire [1:0] _GEN_428 = 6'h1d == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_29_2 : _GEN_427;
  wire [1:0] _GEN_429 = 6'h1d == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_29_3 : _GEN_428;
  wire [1:0] _GEN_430 = 6'h1e == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_30_0 : _GEN_429;
  wire [1:0] _GEN_431 = 6'h1e == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_30_1 : _GEN_430;
  wire [1:0] _GEN_432 = 6'h1e == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_30_2 : _GEN_431;
  wire [1:0] _GEN_433 = 6'h1e == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_30_3 : _GEN_432;
  wire [1:0] _GEN_434 = 6'h1f == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_31_0 : _GEN_433;
  wire [1:0] _GEN_435 = 6'h1f == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_31_1 : _GEN_434;
  wire [1:0] _GEN_436 = 6'h1f == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_31_2 : _GEN_435;
  wire [1:0] _GEN_437 = 6'h1f == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_31_3 : _GEN_436;
  wire [1:0] _GEN_438 = 6'h20 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_32_0 : _GEN_437;
  wire [1:0] _GEN_439 = 6'h20 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_32_1 : _GEN_438;
  wire [1:0] _GEN_440 = 6'h20 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_32_2 : _GEN_439;
  wire [1:0] _GEN_441 = 6'h20 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_32_3 : _GEN_440;
  wire [1:0] _GEN_442 = 6'h21 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_33_0 : _GEN_441;
  wire [1:0] _GEN_443 = 6'h21 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_33_1 : _GEN_442;
  wire [1:0] _GEN_444 = 6'h21 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_33_2 : _GEN_443;
  wire [1:0] _GEN_445 = 6'h21 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_33_3 : _GEN_444;
  wire [1:0] _GEN_446 = 6'h22 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_34_0 : _GEN_445;
  wire [1:0] _GEN_447 = 6'h22 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_34_1 : _GEN_446;
  wire [1:0] _GEN_448 = 6'h22 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_34_2 : _GEN_447;
  wire [1:0] _GEN_449 = 6'h22 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_34_3 : _GEN_448;
  wire [1:0] _GEN_450 = 6'h23 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_35_0 : _GEN_449;
  wire [1:0] _GEN_451 = 6'h23 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_35_1 : _GEN_450;
  wire [1:0] _GEN_452 = 6'h23 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_35_2 : _GEN_451;
  wire [1:0] _GEN_453 = 6'h23 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_35_3 : _GEN_452;
  wire [1:0] _GEN_454 = 6'h24 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_36_0 : _GEN_453;
  wire [1:0] _GEN_455 = 6'h24 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_36_1 : _GEN_454;
  wire [1:0] _GEN_456 = 6'h24 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_36_2 : _GEN_455;
  wire [1:0] _GEN_457 = 6'h24 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_36_3 : _GEN_456;
  wire [1:0] _GEN_458 = 6'h25 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_37_0 : _GEN_457;
  wire [1:0] _GEN_459 = 6'h25 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_37_1 : _GEN_458;
  wire [1:0] _GEN_460 = 6'h25 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_37_2 : _GEN_459;
  wire [1:0] _GEN_461 = 6'h25 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_37_3 : _GEN_460;
  wire [1:0] _GEN_462 = 6'h26 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_38_0 : _GEN_461;
  wire [1:0] _GEN_463 = 6'h26 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_38_1 : _GEN_462;
  wire [1:0] _GEN_464 = 6'h26 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_38_2 : _GEN_463;
  wire [1:0] _GEN_465 = 6'h26 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_38_3 : _GEN_464;
  wire [1:0] _GEN_466 = 6'h27 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_39_0 : _GEN_465;
  wire [1:0] _GEN_467 = 6'h27 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_39_1 : _GEN_466;
  wire [1:0] _GEN_468 = 6'h27 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_39_2 : _GEN_467;
  wire [1:0] _GEN_469 = 6'h27 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_39_3 : _GEN_468;
  wire [1:0] _GEN_470 = 6'h28 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_40_0 : _GEN_469;
  wire [1:0] _GEN_471 = 6'h28 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_40_1 : _GEN_470;
  wire [1:0] _GEN_472 = 6'h28 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_40_2 : _GEN_471;
  wire [1:0] _GEN_473 = 6'h28 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_40_3 : _GEN_472;
  wire [1:0] _GEN_474 = 6'h29 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_41_0 : _GEN_473;
  wire [1:0] _GEN_475 = 6'h29 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_41_1 : _GEN_474;
  wire [1:0] _GEN_476 = 6'h29 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_41_2 : _GEN_475;
  wire [1:0] _GEN_477 = 6'h29 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_41_3 : _GEN_476;
  wire [1:0] _GEN_478 = 6'h2a == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_42_0 : _GEN_477;
  wire [1:0] _GEN_479 = 6'h2a == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_42_1 : _GEN_478;
  wire [1:0] _GEN_480 = 6'h2a == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_42_2 : _GEN_479;
  wire [1:0] _GEN_481 = 6'h2a == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_42_3 : _GEN_480;
  wire [1:0] _GEN_482 = 6'h2b == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_43_0 : _GEN_481;
  wire [1:0] _GEN_483 = 6'h2b == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_43_1 : _GEN_482;
  wire [1:0] _GEN_484 = 6'h2b == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_43_2 : _GEN_483;
  wire [1:0] _GEN_485 = 6'h2b == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_43_3 : _GEN_484;
  wire [1:0] _GEN_486 = 6'h2c == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_44_0 : _GEN_485;
  wire [1:0] _GEN_487 = 6'h2c == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_44_1 : _GEN_486;
  wire [1:0] _GEN_488 = 6'h2c == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_44_2 : _GEN_487;
  wire [1:0] _GEN_489 = 6'h2c == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_44_3 : _GEN_488;
  wire [1:0] _GEN_490 = 6'h2d == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_45_0 : _GEN_489;
  wire [1:0] _GEN_491 = 6'h2d == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_45_1 : _GEN_490;
  wire [1:0] _GEN_492 = 6'h2d == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_45_2 : _GEN_491;
  wire [1:0] _GEN_493 = 6'h2d == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_45_3 : _GEN_492;
  wire [1:0] _GEN_494 = 6'h2e == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_46_0 : _GEN_493;
  wire [1:0] _GEN_495 = 6'h2e == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_46_1 : _GEN_494;
  wire [1:0] _GEN_496 = 6'h2e == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_46_2 : _GEN_495;
  wire [1:0] _GEN_497 = 6'h2e == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_46_3 : _GEN_496;
  wire [1:0] _GEN_498 = 6'h2f == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_47_0 : _GEN_497;
  wire [1:0] _GEN_499 = 6'h2f == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_47_1 : _GEN_498;
  wire [1:0] _GEN_500 = 6'h2f == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_47_2 : _GEN_499;
  wire [1:0] _GEN_501 = 6'h2f == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_47_3 : _GEN_500;
  wire [1:0] _GEN_502 = 6'h30 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_48_0 : _GEN_501;
  wire [1:0] _GEN_503 = 6'h30 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_48_1 : _GEN_502;
  wire [1:0] _GEN_504 = 6'h30 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_48_2 : _GEN_503;
  wire [1:0] _GEN_505 = 6'h30 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_48_3 : _GEN_504;
  wire [1:0] _GEN_506 = 6'h31 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_49_0 : _GEN_505;
  wire [1:0] _GEN_507 = 6'h31 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_49_1 : _GEN_506;
  wire [1:0] _GEN_508 = 6'h31 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_49_2 : _GEN_507;
  wire [1:0] _GEN_509 = 6'h31 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_49_3 : _GEN_508;
  wire [1:0] _GEN_510 = 6'h32 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_50_0 : _GEN_509;
  wire [1:0] _GEN_511 = 6'h32 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_50_1 : _GEN_510;
  wire [1:0] _GEN_512 = 6'h32 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_50_2 : _GEN_511;
  wire [1:0] _GEN_513 = 6'h32 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_50_3 : _GEN_512;
  wire [1:0] _GEN_514 = 6'h33 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_51_0 : _GEN_513;
  wire [1:0] _GEN_515 = 6'h33 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_51_1 : _GEN_514;
  wire [1:0] _GEN_516 = 6'h33 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_51_2 : _GEN_515;
  wire [1:0] _GEN_517 = 6'h33 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_51_3 : _GEN_516;
  wire [1:0] _GEN_518 = 6'h34 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_52_0 : _GEN_517;
  wire [1:0] _GEN_519 = 6'h34 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_52_1 : _GEN_518;
  wire [1:0] _GEN_520 = 6'h34 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_52_2 : _GEN_519;
  wire [1:0] _GEN_521 = 6'h34 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_52_3 : _GEN_520;
  wire [1:0] _GEN_522 = 6'h35 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_53_0 : _GEN_521;
  wire [1:0] _GEN_523 = 6'h35 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_53_1 : _GEN_522;
  wire [1:0] _GEN_524 = 6'h35 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_53_2 : _GEN_523;
  wire [1:0] _GEN_525 = 6'h35 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_53_3 : _GEN_524;
  wire [1:0] _GEN_526 = 6'h36 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_54_0 : _GEN_525;
  wire [1:0] _GEN_527 = 6'h36 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_54_1 : _GEN_526;
  wire [1:0] _GEN_528 = 6'h36 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_54_2 : _GEN_527;
  wire [1:0] _GEN_529 = 6'h36 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_54_3 : _GEN_528;
  wire [1:0] _GEN_530 = 6'h37 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_55_0 : _GEN_529;
  wire [1:0] _GEN_531 = 6'h37 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_55_1 : _GEN_530;
  wire [1:0] _GEN_532 = 6'h37 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_55_2 : _GEN_531;
  wire [1:0] _GEN_533 = 6'h37 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_55_3 : _GEN_532;
  wire [1:0] _GEN_534 = 6'h38 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_56_0 : _GEN_533;
  wire [1:0] _GEN_535 = 6'h38 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_56_1 : _GEN_534;
  wire [1:0] _GEN_536 = 6'h38 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_56_2 : _GEN_535;
  wire [1:0] _GEN_537 = 6'h38 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_56_3 : _GEN_536;
  wire [1:0] _GEN_538 = 6'h39 == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_57_0 : _GEN_537;
  wire [1:0] _GEN_539 = 6'h39 == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_57_1 : _GEN_538;
  wire [1:0] _GEN_540 = 6'h39 == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_57_2 : _GEN_539;
  wire [1:0] _GEN_541 = 6'h39 == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_57_3 : _GEN_540;
  wire [1:0] _GEN_542 = 6'h3a == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_58_0 : _GEN_541;
  wire [1:0] _GEN_543 = 6'h3a == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_58_1 : _GEN_542;
  wire [1:0] _GEN_544 = 6'h3a == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_58_2 : _GEN_543;
  wire [1:0] _GEN_545 = 6'h3a == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_58_3 : _GEN_544;
  wire [1:0] _GEN_546 = 6'h3b == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_59_0 : _GEN_545;
  wire [1:0] _GEN_547 = 6'h3b == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_59_1 : _GEN_546;
  wire [1:0] _GEN_548 = 6'h3b == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_59_2 : _GEN_547;
  wire [1:0] _GEN_549 = 6'h3b == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_59_3 : _GEN_548;
  wire [1:0] _GEN_550 = 6'h3c == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_60_0 : _GEN_549;
  wire [1:0] _GEN_551 = 6'h3c == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_60_1 : _GEN_550;
  wire [1:0] _GEN_552 = 6'h3c == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_60_2 : _GEN_551;
  wire [1:0] _GEN_553 = 6'h3c == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_60_3 : _GEN_552;
  wire [1:0] _GEN_554 = 6'h3d == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_61_0 : _GEN_553;
  wire [1:0] _GEN_555 = 6'h3d == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_61_1 : _GEN_554;
  wire [1:0] _GEN_556 = 6'h3d == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_61_2 : _GEN_555;
  wire [1:0] _GEN_557 = 6'h3d == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_61_3 : _GEN_556;
  wire [1:0] _GEN_558 = 6'h3e == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_62_0 : _GEN_557;
  wire [1:0] _GEN_559 = 6'h3e == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_62_1 : _GEN_558;
  wire [1:0] _GEN_560 = 6'h3e == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_62_2 : _GEN_559;
  wire [1:0] _GEN_561 = 6'h3e == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_62_3 : _GEN_560;
  wire [1:0] _GEN_562 = 6'h3f == req_addr_index & 2'h0 == s2_idxWayHit ? regCount_63_0 : _GEN_561;
  wire [1:0] _GEN_563 = 6'h3f == req_addr_index & 2'h1 == s2_idxWayHit ? regCount_63_1 : _GEN_562;
  wire [1:0] _GEN_564 = 6'h3f == req_addr_index & 2'h2 == s2_idxWayHit ? regCount_63_2 : _GEN_563;
  wire [1:0] _GEN_565 = 6'h3f == req_addr_index & 2'h3 == s2_idxWayHit ? regCount_63_3 : _GEN_564;
  wire [1:0] _newCountHit_0_T_1 = _GEN_74 + 2'h1;
  wire [1:0] _GEN_566 = _GEN_74 < _GEN_565 ? _newCountHit_0_T_1 : _GEN_74;
  wire [1:0] newCountHit_0 = 2'h0 != s2_idxWayHit ? _GEN_566 : 2'h0;
  wire [1:0] _newCountHit_1_T_1 = _GEN_138 + 2'h1;
  wire [1:0] _GEN_568 = _GEN_138 < _GEN_565 ? _newCountHit_1_T_1 : _GEN_138;
  wire [1:0] newCountHit_1 = 2'h1 != s2_idxWayHit ? _GEN_568 : 2'h0;
  wire [1:0] _newCountHit_2_T_1 = _GEN_202 + 2'h1;
  wire [1:0] _GEN_570 = _GEN_202 < _GEN_565 ? _newCountHit_2_T_1 : _GEN_202;
  wire [1:0] newCountHit_2 = 2'h2 != s2_idxWayHit ? _GEN_570 : 2'h0;
  wire [1:0] _newCountHit_3_T_1 = _GEN_266 + 2'h1;
  wire [1:0] _GEN_572 = _GEN_266 < _GEN_565 ? _newCountHit_3_T_1 : _GEN_266;
  wire [1:0] newCountHit_3 = 2'h3 != s2_idxWayHit ? _GEN_572 : 2'h0;
  wire [1:0] _GEN_574 = metaWays_0_valid ? _newCountHit_0_T_1 : _GEN_74;
  wire [1:0] newCountRefill_0 = 2'h0 == selectWay ? 2'h0 : _GEN_574;
  wire [1:0] _GEN_576 = metaWays_1_valid ? _newCountHit_1_T_1 : _GEN_138;
  wire [1:0] newCountRefill_1 = 2'h1 == selectWay ? 2'h0 : _GEN_576;
  wire [1:0] _GEN_578 = metaWays_2_valid ? _newCountHit_2_T_1 : _GEN_202;
  wire [1:0] newCountRefill_2 = 2'h2 == selectWay ? 2'h0 : _GEN_578;
  wire [1:0] _GEN_580 = metaWays_3_valid ? _newCountHit_3_T_1 : _GEN_266;
  wire [1:0] newCountRefill_3 = 2'h3 == selectWay ? 2'h0 : _GEN_580;
  wire  countUpdate = hitUpdate | memRespUpdate;
  wire [31:0] _WIRE_9 = {{26'd0}, req_addr_index};
  wire  hitRespValid = _cacheUpdate_T_2 & s2_hit;
  wire [21:0] _GEN_1095 = 2'h1 == selectWay ? metaWays_1_tag : metaWays_0_tag;
  wire [21:0] _GEN_1096 = 2'h2 == selectWay ? metaWays_2_tag : _GEN_1095;
  wire [21:0] _GEN_1097 = 2'h3 == selectWay ? metaWays_3_tag : _GEN_1096;
  wire [31:0] writeBackAddr = {_GEN_1097,req_addr_index,4'h0};
  wire  _x1_T = c_state == 3'h4;
  wire [63:0] _GEN_1099 = 2'h1 == selectWay ? dataWays_1_1 : dataWays_0_1;
  wire [63:0] _GEN_1100 = 2'h2 == selectWay ? dataWays_2_1 : _GEN_1099;
  wire [63:0] _GEN_1101 = 2'h3 == selectWay ? dataWays_3_1 : _GEN_1100;
  wire [63:0] _GEN_1103 = 2'h1 == selectWay ? dataWays_1_0 : dataWays_0_0;
  wire [63:0] _GEN_1104 = 2'h2 == selectWay ? dataWays_2_0 : _GEN_1103;
  wire [63:0] _GEN_1105 = 2'h3 == selectWay ? dataWays_3_0 : _GEN_1104;
  wire [127:0] _x2_T_1 = {_GEN_1101,_GEN_1105};
  wire  probeCheck = _hitUpdate_T & s2_reg_probe;
  wire  probeResp = c_state == 3'h6;
  wire [2:0] _linkCmd_T = s2_hit ? 3'h5 : 3'h6;
  ysyx_040656_SRAM metaArray_0 (
    .clock(metaArray_0_clock),
    .reset(metaArray_0_reset),
    .io_w_setIdx(metaArray_0_io_w_setIdx),
    .io_w_data_tag(metaArray_0_io_w_data_tag),
    .io_w_data_valid(metaArray_0_io_w_data_valid),
    .io_w_data_needFlush(metaArray_0_io_w_data_needFlush),
    .io_w_wen(metaArray_0_io_w_wen),
    .io_r_setIdx(metaArray_0_io_r_setIdx),
    .io_r_data_tag(metaArray_0_io_r_data_tag),
    .io_r_data_valid(metaArray_0_io_r_data_valid),
    .io_r_data_needFlush(metaArray_0_io_r_data_needFlush),
    .io_r_ren(metaArray_0_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_1 (
    .clock(metaArray_1_clock),
    .reset(metaArray_1_reset),
    .io_w_setIdx(metaArray_1_io_w_setIdx),
    .io_w_data_tag(metaArray_1_io_w_data_tag),
    .io_w_data_valid(metaArray_1_io_w_data_valid),
    .io_w_data_needFlush(metaArray_1_io_w_data_needFlush),
    .io_w_wen(metaArray_1_io_w_wen),
    .io_r_setIdx(metaArray_1_io_r_setIdx),
    .io_r_data_tag(metaArray_1_io_r_data_tag),
    .io_r_data_valid(metaArray_1_io_r_data_valid),
    .io_r_data_needFlush(metaArray_1_io_r_data_needFlush),
    .io_r_ren(metaArray_1_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_2 (
    .clock(metaArray_2_clock),
    .reset(metaArray_2_reset),
    .io_w_setIdx(metaArray_2_io_w_setIdx),
    .io_w_data_tag(metaArray_2_io_w_data_tag),
    .io_w_data_valid(metaArray_2_io_w_data_valid),
    .io_w_data_needFlush(metaArray_2_io_w_data_needFlush),
    .io_w_wen(metaArray_2_io_w_wen),
    .io_r_setIdx(metaArray_2_io_r_setIdx),
    .io_r_data_tag(metaArray_2_io_r_data_tag),
    .io_r_data_valid(metaArray_2_io_r_data_valid),
    .io_r_data_needFlush(metaArray_2_io_r_data_needFlush),
    .io_r_ren(metaArray_2_io_r_ren)
  );
  ysyx_040656_SRAM metaArray_3 (
    .clock(metaArray_3_clock),
    .reset(metaArray_3_reset),
    .io_w_setIdx(metaArray_3_io_w_setIdx),
    .io_w_data_tag(metaArray_3_io_w_data_tag),
    .io_w_data_valid(metaArray_3_io_w_data_valid),
    .io_w_data_needFlush(metaArray_3_io_w_data_needFlush),
    .io_w_wen(metaArray_3_io_w_wen),
    .io_r_setIdx(metaArray_3_io_r_setIdx),
    .io_r_data_tag(metaArray_3_io_r_data_tag),
    .io_r_data_valid(metaArray_3_io_r_data_valid),
    .io_r_data_needFlush(metaArray_3_io_r_data_needFlush),
    .io_r_ren(metaArray_3_io_r_ren)
  );
  ysyx_040656_Arbiter arbiter (
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_wdata(arbiter_io_in_1_bits_wdata),
    .io_in_1_bits_size(arbiter_io_in_1_bits_size),
    .io_in_1_bits_cmd(arbiter_io_in_1_bits_cmd),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_size(arbiter_io_out_bits_size),
    .io_out_bits_cmd(arbiter_io_out_bits_cmd)
  );
  ysyx_040656_LRU selTree (
    .io_inWayValid_0(selTree_io_inWayValid_0),
    .io_inWayValid_1(selTree_io_inWayValid_1),
    .io_inWayValid_2(selTree_io_inWayValid_2),
    .io_inWayValid_3(selTree_io_inWayValid_3),
    .io_inValue_0(selTree_io_inValue_0),
    .io_inValue_1(selTree_io_inValue_1),
    .io_inValue_2(selTree_io_inValue_2),
    .io_inValue_3(selTree_io_inValue_3),
    .io_outIdx(selTree_io_outIdx)
  );
  assign io_in_req_ready = arbiter_io_in_1_ready;
  assign io_in_resp_valid = hitRespValid & _noprobeStall_T;
  assign io_in_resp_bits_rdata = rWord >> shift;
  assign io_out_req_valid = c_state == 3'h2 | _x1_T;
  assign io_out_req_bits_addr = c_state == 3'h4 ? writeBackAddr : _s1_strb_T;
  assign io_out_req_bits_wdata = c_state == 3'h4 ? _x2_T_1 : 128'h0;
  assign io_out_req_bits_cmd = {{2'd0}, _x1_T};
  assign io_out_resp_ready = 1'h1;
  assign io_link_req_ready = arbiter_io_in_0_ready;
  assign io_link_resp_valid = probeCheck | probeResp;
  assign io_link_resp_bits_cmd = probeResp ? 3'h3 : _linkCmd_T;
  assign io_link_resp_bits_rdata = {s2_dataBlockHit_1,s2_dataBlockHit_0};
  assign io_dataArray_0_wen = ~(reset | _metaArray_0_io_w_wen_T_1);
  assign io_dataArray_0_addr = _GEN_0[9:4];
  assign io_dataArray_0_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_1_wen = ~(reset | _metaArray_1_io_w_wen_T_1);
  assign io_dataArray_1_addr = _GEN_0[9:4];
  assign io_dataArray_1_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_2_wen = ~(reset | _metaArray_2_io_w_wen_T_1);
  assign io_dataArray_2_addr = _GEN_0[9:4];
  assign io_dataArray_2_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign io_dataArray_3_wen = ~(reset | _metaArray_3_io_w_wen_T_1);
  assign io_dataArray_3_addr = _GEN_0[9:4];
  assign io_dataArray_3_wdata = reset ? 128'h0 : _io_dataArray_0_wdata_T_1;
  assign metaArray_0_clock = clock;
  assign metaArray_0_reset = reset;
  assign metaArray_0_io_w_setIdx = _GEN_0[9:4];
  assign metaArray_0_io_w_data_tag = memRespUpdate ? req_addr_tag : newMetaDirty_tag;
  assign metaArray_0_io_w_data_valid = memRespUpdate | newMetaDirty_valid;
  assign metaArray_0_io_w_data_needFlush = memRespUpdate ? 1'h0 : newMetaDirty_needFlush;
  assign metaArray_0_io_w_wen = cacheUpdate & 2'h0 == wayWrite;
  assign metaArray_0_io_r_setIdx = _GEN_0[9:4];
  assign metaArray_0_io_r_ren = ~cacheUpdate;
  assign metaArray_1_clock = clock;
  assign metaArray_1_reset = reset;
  assign metaArray_1_io_w_setIdx = _GEN_0[9:4];
  assign metaArray_1_io_w_data_tag = memRespUpdate ? req_addr_tag : newMetaDirty_tag;
  assign metaArray_1_io_w_data_valid = memRespUpdate | newMetaDirty_valid;
  assign metaArray_1_io_w_data_needFlush = memRespUpdate ? 1'h0 : newMetaDirty_needFlush;
  assign metaArray_1_io_w_wen = cacheUpdate & 2'h1 == wayWrite;
  assign metaArray_1_io_r_setIdx = _GEN_0[9:4];
  assign metaArray_1_io_r_ren = ~cacheUpdate;
  assign metaArray_2_clock = clock;
  assign metaArray_2_reset = reset;
  assign metaArray_2_io_w_setIdx = _GEN_0[9:4];
  assign metaArray_2_io_w_data_tag = memRespUpdate ? req_addr_tag : newMetaDirty_tag;
  assign metaArray_2_io_w_data_valid = memRespUpdate | newMetaDirty_valid;
  assign metaArray_2_io_w_data_needFlush = memRespUpdate ? 1'h0 : newMetaDirty_needFlush;
  assign metaArray_2_io_w_wen = cacheUpdate & 2'h2 == wayWrite;
  assign metaArray_2_io_r_setIdx = _GEN_0[9:4];
  assign metaArray_2_io_r_ren = ~cacheUpdate;
  assign metaArray_3_clock = clock;
  assign metaArray_3_reset = reset;
  assign metaArray_3_io_w_setIdx = _GEN_0[9:4];
  assign metaArray_3_io_w_data_tag = memRespUpdate ? req_addr_tag : newMetaDirty_tag;
  assign metaArray_3_io_w_data_valid = memRespUpdate | newMetaDirty_valid;
  assign metaArray_3_io_w_data_needFlush = memRespUpdate ? 1'h0 : newMetaDirty_needFlush;
  assign metaArray_3_io_w_wen = cacheUpdate & 2'h3 == wayWrite;
  assign metaArray_3_io_r_setIdx = _GEN_0[9:4];
  assign metaArray_3_io_r_ren = ~cacheUpdate;
  assign arbiter_io_in_0_valid = io_link_req_valid;
  assign arbiter_io_in_0_bits_addr = io_link_req_bits_addr;
  assign arbiter_io_in_0_bits_wdata = io_link_req_bits_wdata;
  assign arbiter_io_in_1_valid = io_in_req_valid;
  assign arbiter_io_in_1_bits_addr = io_in_req_bits_addr;
  assign arbiter_io_in_1_bits_wdata = {{64'd0}, io_in_req_bits_wdata};
  assign arbiter_io_in_1_bits_size = io_in_req_bits_size;
  assign arbiter_io_in_1_bits_cmd = io_in_req_bits_cmd;
  assign arbiter_io_out_ready = c_state == 3'h0;
  assign selTree_io_inWayValid_0 = metaArray_0_io_r_data_valid;
  assign selTree_io_inWayValid_1 = metaArray_1_io_r_data_valid;
  assign selTree_io_inWayValid_2 = metaArray_2_io_r_data_valid;
  assign selTree_io_inWayValid_3 = metaArray_3_io_r_data_valid;
  assign selTree_io_inValue_0 = 6'h3f == req_addr_index ? regCount_63_0 : _GEN_73;
  assign selTree_io_inValue_1 = 6'h3f == req_addr_index ? regCount_63_1 : _GEN_137;
  assign selTree_io_inValue_2 = 6'h3f == req_addr_index ? regCount_63_2 : _GEN_201;
  assign selTree_io_inValue_3 = 6'h3f == req_addr_index ? regCount_63_3 : _GEN_265;
  always @(posedge clock) begin
    if (reset) begin
      c_state <= 3'h0;
    end else if (3'h0 == c_state) begin
      if (s1_valid) begin
        c_state <= 3'h1;
      end
    end else if (3'h1 == c_state) begin
      if (_noprobeStall_T) begin
        c_state <= _GEN_278;
      end else begin
        c_state <= _GEN_281;
      end
    end else if (3'h2 == c_state) begin
      c_state <= _GEN_283;
    end else begin
      c_state <= _GEN_293;
    end
    if (reset) begin
      regCount_0_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_0_0 <= newCountRefill_0;
        end else begin
          regCount_0_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_0_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_0_1 <= newCountRefill_1;
        end else begin
          regCount_0_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_0_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_0_2 <= newCountRefill_2;
        end else begin
          regCount_0_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_0_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h0 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_0_3 <= newCountRefill_3;
        end else begin
          regCount_0_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_1_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_1_0 <= newCountRefill_0;
        end else begin
          regCount_1_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_1_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_1_1 <= newCountRefill_1;
        end else begin
          regCount_1_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_1_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_1_2 <= newCountRefill_2;
        end else begin
          regCount_1_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_1_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_1_3 <= newCountRefill_3;
        end else begin
          regCount_1_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_2_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_2_0 <= newCountRefill_0;
        end else begin
          regCount_2_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_2_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_2_1 <= newCountRefill_1;
        end else begin
          regCount_2_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_2_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_2_2 <= newCountRefill_2;
        end else begin
          regCount_2_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_2_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_2_3 <= newCountRefill_3;
        end else begin
          regCount_2_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_3_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_3_0 <= newCountRefill_0;
        end else begin
          regCount_3_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_3_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_3_1 <= newCountRefill_1;
        end else begin
          regCount_3_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_3_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_3_2 <= newCountRefill_2;
        end else begin
          regCount_3_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_3_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_3_3 <= newCountRefill_3;
        end else begin
          regCount_3_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_4_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_4_0 <= newCountRefill_0;
        end else begin
          regCount_4_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_4_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_4_1 <= newCountRefill_1;
        end else begin
          regCount_4_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_4_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_4_2 <= newCountRefill_2;
        end else begin
          regCount_4_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_4_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h4 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_4_3 <= newCountRefill_3;
        end else begin
          regCount_4_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_5_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_5_0 <= newCountRefill_0;
        end else begin
          regCount_5_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_5_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_5_1 <= newCountRefill_1;
        end else begin
          regCount_5_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_5_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_5_2 <= newCountRefill_2;
        end else begin
          regCount_5_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_5_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h5 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_5_3 <= newCountRefill_3;
        end else begin
          regCount_5_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_6_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_6_0 <= newCountRefill_0;
        end else begin
          regCount_6_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_6_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_6_1 <= newCountRefill_1;
        end else begin
          regCount_6_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_6_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_6_2 <= newCountRefill_2;
        end else begin
          regCount_6_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_6_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h6 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_6_3 <= newCountRefill_3;
        end else begin
          regCount_6_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_7_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_7_0 <= newCountRefill_0;
        end else begin
          regCount_7_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_7_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_7_1 <= newCountRefill_1;
        end else begin
          regCount_7_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_7_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_7_2 <= newCountRefill_2;
        end else begin
          regCount_7_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_7_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h7 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_7_3 <= newCountRefill_3;
        end else begin
          regCount_7_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_8_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_8_0 <= newCountRefill_0;
        end else begin
          regCount_8_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_8_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_8_1 <= newCountRefill_1;
        end else begin
          regCount_8_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_8_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_8_2 <= newCountRefill_2;
        end else begin
          regCount_8_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_8_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h8 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_8_3 <= newCountRefill_3;
        end else begin
          regCount_8_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_9_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_9_0 <= newCountRefill_0;
        end else begin
          regCount_9_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_9_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_9_1 <= newCountRefill_1;
        end else begin
          regCount_9_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_9_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_9_2 <= newCountRefill_2;
        end else begin
          regCount_9_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_9_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h9 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_9_3 <= newCountRefill_3;
        end else begin
          regCount_9_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_10_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_10_0 <= newCountRefill_0;
        end else begin
          regCount_10_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_10_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_10_1 <= newCountRefill_1;
        end else begin
          regCount_10_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_10_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_10_2 <= newCountRefill_2;
        end else begin
          regCount_10_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_10_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'ha == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_10_3 <= newCountRefill_3;
        end else begin
          regCount_10_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_11_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_11_0 <= newCountRefill_0;
        end else begin
          regCount_11_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_11_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_11_1 <= newCountRefill_1;
        end else begin
          regCount_11_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_11_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_11_2 <= newCountRefill_2;
        end else begin
          regCount_11_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_11_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hb == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_11_3 <= newCountRefill_3;
        end else begin
          regCount_11_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_12_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_12_0 <= newCountRefill_0;
        end else begin
          regCount_12_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_12_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_12_1 <= newCountRefill_1;
        end else begin
          regCount_12_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_12_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_12_2 <= newCountRefill_2;
        end else begin
          regCount_12_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_12_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hc == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_12_3 <= newCountRefill_3;
        end else begin
          regCount_12_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_13_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_13_0 <= newCountRefill_0;
        end else begin
          regCount_13_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_13_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_13_1 <= newCountRefill_1;
        end else begin
          regCount_13_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_13_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_13_2 <= newCountRefill_2;
        end else begin
          regCount_13_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_13_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hd == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_13_3 <= newCountRefill_3;
        end else begin
          regCount_13_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_14_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_14_0 <= newCountRefill_0;
        end else begin
          regCount_14_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_14_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_14_1 <= newCountRefill_1;
        end else begin
          regCount_14_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_14_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_14_2 <= newCountRefill_2;
        end else begin
          regCount_14_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_14_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'he == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_14_3 <= newCountRefill_3;
        end else begin
          regCount_14_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_15_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_15_0 <= newCountRefill_0;
        end else begin
          regCount_15_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_15_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_15_1 <= newCountRefill_1;
        end else begin
          regCount_15_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_15_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_15_2 <= newCountRefill_2;
        end else begin
          regCount_15_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_15_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'hf == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_15_3 <= newCountRefill_3;
        end else begin
          regCount_15_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_16_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_16_0 <= newCountRefill_0;
        end else begin
          regCount_16_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_16_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_16_1 <= newCountRefill_1;
        end else begin
          regCount_16_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_16_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_16_2 <= newCountRefill_2;
        end else begin
          regCount_16_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_16_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h10 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_16_3 <= newCountRefill_3;
        end else begin
          regCount_16_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_17_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_17_0 <= newCountRefill_0;
        end else begin
          regCount_17_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_17_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_17_1 <= newCountRefill_1;
        end else begin
          regCount_17_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_17_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_17_2 <= newCountRefill_2;
        end else begin
          regCount_17_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_17_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h11 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_17_3 <= newCountRefill_3;
        end else begin
          regCount_17_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_18_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_18_0 <= newCountRefill_0;
        end else begin
          regCount_18_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_18_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_18_1 <= newCountRefill_1;
        end else begin
          regCount_18_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_18_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_18_2 <= newCountRefill_2;
        end else begin
          regCount_18_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_18_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h12 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_18_3 <= newCountRefill_3;
        end else begin
          regCount_18_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_19_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_19_0 <= newCountRefill_0;
        end else begin
          regCount_19_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_19_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_19_1 <= newCountRefill_1;
        end else begin
          regCount_19_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_19_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_19_2 <= newCountRefill_2;
        end else begin
          regCount_19_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_19_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h13 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_19_3 <= newCountRefill_3;
        end else begin
          regCount_19_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_20_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_20_0 <= newCountRefill_0;
        end else begin
          regCount_20_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_20_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_20_1 <= newCountRefill_1;
        end else begin
          regCount_20_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_20_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_20_2 <= newCountRefill_2;
        end else begin
          regCount_20_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_20_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h14 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_20_3 <= newCountRefill_3;
        end else begin
          regCount_20_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_21_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_21_0 <= newCountRefill_0;
        end else begin
          regCount_21_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_21_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_21_1 <= newCountRefill_1;
        end else begin
          regCount_21_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_21_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_21_2 <= newCountRefill_2;
        end else begin
          regCount_21_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_21_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h15 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_21_3 <= newCountRefill_3;
        end else begin
          regCount_21_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_22_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_22_0 <= newCountRefill_0;
        end else begin
          regCount_22_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_22_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_22_1 <= newCountRefill_1;
        end else begin
          regCount_22_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_22_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_22_2 <= newCountRefill_2;
        end else begin
          regCount_22_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_22_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h16 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_22_3 <= newCountRefill_3;
        end else begin
          regCount_22_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_23_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_23_0 <= newCountRefill_0;
        end else begin
          regCount_23_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_23_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_23_1 <= newCountRefill_1;
        end else begin
          regCount_23_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_23_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_23_2 <= newCountRefill_2;
        end else begin
          regCount_23_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_23_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h17 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_23_3 <= newCountRefill_3;
        end else begin
          regCount_23_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_24_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_24_0 <= newCountRefill_0;
        end else begin
          regCount_24_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_24_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_24_1 <= newCountRefill_1;
        end else begin
          regCount_24_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_24_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_24_2 <= newCountRefill_2;
        end else begin
          regCount_24_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_24_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h18 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_24_3 <= newCountRefill_3;
        end else begin
          regCount_24_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_25_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_25_0 <= newCountRefill_0;
        end else begin
          regCount_25_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_25_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_25_1 <= newCountRefill_1;
        end else begin
          regCount_25_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_25_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_25_2 <= newCountRefill_2;
        end else begin
          regCount_25_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_25_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h19 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_25_3 <= newCountRefill_3;
        end else begin
          regCount_25_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_26_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_26_0 <= newCountRefill_0;
        end else begin
          regCount_26_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_26_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_26_1 <= newCountRefill_1;
        end else begin
          regCount_26_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_26_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_26_2 <= newCountRefill_2;
        end else begin
          regCount_26_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_26_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_26_3 <= newCountRefill_3;
        end else begin
          regCount_26_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_27_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_27_0 <= newCountRefill_0;
        end else begin
          regCount_27_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_27_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_27_1 <= newCountRefill_1;
        end else begin
          regCount_27_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_27_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_27_2 <= newCountRefill_2;
        end else begin
          regCount_27_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_27_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_27_3 <= newCountRefill_3;
        end else begin
          regCount_27_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_28_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_28_0 <= newCountRefill_0;
        end else begin
          regCount_28_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_28_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_28_1 <= newCountRefill_1;
        end else begin
          regCount_28_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_28_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_28_2 <= newCountRefill_2;
        end else begin
          regCount_28_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_28_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_28_3 <= newCountRefill_3;
        end else begin
          regCount_28_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_29_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_29_0 <= newCountRefill_0;
        end else begin
          regCount_29_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_29_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_29_1 <= newCountRefill_1;
        end else begin
          regCount_29_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_29_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_29_2 <= newCountRefill_2;
        end else begin
          regCount_29_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_29_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_29_3 <= newCountRefill_3;
        end else begin
          regCount_29_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_30_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_30_0 <= newCountRefill_0;
        end else begin
          regCount_30_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_30_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_30_1 <= newCountRefill_1;
        end else begin
          regCount_30_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_30_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_30_2 <= newCountRefill_2;
        end else begin
          regCount_30_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_30_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_30_3 <= newCountRefill_3;
        end else begin
          regCount_30_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_31_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_31_0 <= newCountRefill_0;
        end else begin
          regCount_31_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_31_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_31_1 <= newCountRefill_1;
        end else begin
          regCount_31_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_31_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_31_2 <= newCountRefill_2;
        end else begin
          regCount_31_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_31_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h1f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_31_3 <= newCountRefill_3;
        end else begin
          regCount_31_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_32_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_32_0 <= newCountRefill_0;
        end else begin
          regCount_32_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_32_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_32_1 <= newCountRefill_1;
        end else begin
          regCount_32_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_32_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_32_2 <= newCountRefill_2;
        end else begin
          regCount_32_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_32_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h20 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_32_3 <= newCountRefill_3;
        end else begin
          regCount_32_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_33_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_33_0 <= newCountRefill_0;
        end else begin
          regCount_33_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_33_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_33_1 <= newCountRefill_1;
        end else begin
          regCount_33_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_33_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_33_2 <= newCountRefill_2;
        end else begin
          regCount_33_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_33_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h21 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_33_3 <= newCountRefill_3;
        end else begin
          regCount_33_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_34_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_34_0 <= newCountRefill_0;
        end else begin
          regCount_34_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_34_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_34_1 <= newCountRefill_1;
        end else begin
          regCount_34_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_34_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_34_2 <= newCountRefill_2;
        end else begin
          regCount_34_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_34_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h22 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_34_3 <= newCountRefill_3;
        end else begin
          regCount_34_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_35_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_35_0 <= newCountRefill_0;
        end else begin
          regCount_35_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_35_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_35_1 <= newCountRefill_1;
        end else begin
          regCount_35_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_35_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_35_2 <= newCountRefill_2;
        end else begin
          regCount_35_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_35_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h23 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_35_3 <= newCountRefill_3;
        end else begin
          regCount_35_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_36_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_36_0 <= newCountRefill_0;
        end else begin
          regCount_36_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_36_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_36_1 <= newCountRefill_1;
        end else begin
          regCount_36_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_36_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_36_2 <= newCountRefill_2;
        end else begin
          regCount_36_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_36_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h24 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_36_3 <= newCountRefill_3;
        end else begin
          regCount_36_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_37_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_37_0 <= newCountRefill_0;
        end else begin
          regCount_37_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_37_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_37_1 <= newCountRefill_1;
        end else begin
          regCount_37_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_37_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_37_2 <= newCountRefill_2;
        end else begin
          regCount_37_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_37_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h25 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_37_3 <= newCountRefill_3;
        end else begin
          regCount_37_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_38_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_38_0 <= newCountRefill_0;
        end else begin
          regCount_38_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_38_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_38_1 <= newCountRefill_1;
        end else begin
          regCount_38_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_38_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_38_2 <= newCountRefill_2;
        end else begin
          regCount_38_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_38_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h26 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_38_3 <= newCountRefill_3;
        end else begin
          regCount_38_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_39_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_39_0 <= newCountRefill_0;
        end else begin
          regCount_39_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_39_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_39_1 <= newCountRefill_1;
        end else begin
          regCount_39_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_39_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_39_2 <= newCountRefill_2;
        end else begin
          regCount_39_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_39_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h27 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_39_3 <= newCountRefill_3;
        end else begin
          regCount_39_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_40_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_40_0 <= newCountRefill_0;
        end else begin
          regCount_40_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_40_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_40_1 <= newCountRefill_1;
        end else begin
          regCount_40_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_40_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_40_2 <= newCountRefill_2;
        end else begin
          regCount_40_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_40_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h28 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_40_3 <= newCountRefill_3;
        end else begin
          regCount_40_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_41_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_41_0 <= newCountRefill_0;
        end else begin
          regCount_41_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_41_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_41_1 <= newCountRefill_1;
        end else begin
          regCount_41_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_41_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_41_2 <= newCountRefill_2;
        end else begin
          regCount_41_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_41_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h29 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_41_3 <= newCountRefill_3;
        end else begin
          regCount_41_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_42_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_42_0 <= newCountRefill_0;
        end else begin
          regCount_42_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_42_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_42_1 <= newCountRefill_1;
        end else begin
          regCount_42_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_42_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_42_2 <= newCountRefill_2;
        end else begin
          regCount_42_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_42_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_42_3 <= newCountRefill_3;
        end else begin
          regCount_42_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_43_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_43_0 <= newCountRefill_0;
        end else begin
          regCount_43_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_43_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_43_1 <= newCountRefill_1;
        end else begin
          regCount_43_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_43_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_43_2 <= newCountRefill_2;
        end else begin
          regCount_43_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_43_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_43_3 <= newCountRefill_3;
        end else begin
          regCount_43_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_44_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_44_0 <= newCountRefill_0;
        end else begin
          regCount_44_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_44_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_44_1 <= newCountRefill_1;
        end else begin
          regCount_44_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_44_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_44_2 <= newCountRefill_2;
        end else begin
          regCount_44_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_44_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_44_3 <= newCountRefill_3;
        end else begin
          regCount_44_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_45_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_45_0 <= newCountRefill_0;
        end else begin
          regCount_45_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_45_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_45_1 <= newCountRefill_1;
        end else begin
          regCount_45_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_45_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_45_2 <= newCountRefill_2;
        end else begin
          regCount_45_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_45_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_45_3 <= newCountRefill_3;
        end else begin
          regCount_45_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_46_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_46_0 <= newCountRefill_0;
        end else begin
          regCount_46_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_46_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_46_1 <= newCountRefill_1;
        end else begin
          regCount_46_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_46_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_46_2 <= newCountRefill_2;
        end else begin
          regCount_46_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_46_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_46_3 <= newCountRefill_3;
        end else begin
          regCount_46_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_47_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_47_0 <= newCountRefill_0;
        end else begin
          regCount_47_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_47_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_47_1 <= newCountRefill_1;
        end else begin
          regCount_47_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_47_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_47_2 <= newCountRefill_2;
        end else begin
          regCount_47_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_47_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h2f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_47_3 <= newCountRefill_3;
        end else begin
          regCount_47_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_48_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_48_0 <= newCountRefill_0;
        end else begin
          regCount_48_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_48_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_48_1 <= newCountRefill_1;
        end else begin
          regCount_48_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_48_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_48_2 <= newCountRefill_2;
        end else begin
          regCount_48_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_48_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h30 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_48_3 <= newCountRefill_3;
        end else begin
          regCount_48_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_49_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_49_0 <= newCountRefill_0;
        end else begin
          regCount_49_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_49_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_49_1 <= newCountRefill_1;
        end else begin
          regCount_49_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_49_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_49_2 <= newCountRefill_2;
        end else begin
          regCount_49_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_49_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h31 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_49_3 <= newCountRefill_3;
        end else begin
          regCount_49_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_50_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_50_0 <= newCountRefill_0;
        end else begin
          regCount_50_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_50_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_50_1 <= newCountRefill_1;
        end else begin
          regCount_50_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_50_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_50_2 <= newCountRefill_2;
        end else begin
          regCount_50_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_50_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h32 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_50_3 <= newCountRefill_3;
        end else begin
          regCount_50_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_51_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_51_0 <= newCountRefill_0;
        end else begin
          regCount_51_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_51_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_51_1 <= newCountRefill_1;
        end else begin
          regCount_51_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_51_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_51_2 <= newCountRefill_2;
        end else begin
          regCount_51_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_51_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h33 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_51_3 <= newCountRefill_3;
        end else begin
          regCount_51_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_52_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_52_0 <= newCountRefill_0;
        end else begin
          regCount_52_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_52_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_52_1 <= newCountRefill_1;
        end else begin
          regCount_52_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_52_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_52_2 <= newCountRefill_2;
        end else begin
          regCount_52_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_52_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h34 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_52_3 <= newCountRefill_3;
        end else begin
          regCount_52_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_53_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_53_0 <= newCountRefill_0;
        end else begin
          regCount_53_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_53_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_53_1 <= newCountRefill_1;
        end else begin
          regCount_53_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_53_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_53_2 <= newCountRefill_2;
        end else begin
          regCount_53_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_53_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h35 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_53_3 <= newCountRefill_3;
        end else begin
          regCount_53_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_54_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_54_0 <= newCountRefill_0;
        end else begin
          regCount_54_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_54_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_54_1 <= newCountRefill_1;
        end else begin
          regCount_54_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_54_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_54_2 <= newCountRefill_2;
        end else begin
          regCount_54_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_54_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h36 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_54_3 <= newCountRefill_3;
        end else begin
          regCount_54_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_55_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_55_0 <= newCountRefill_0;
        end else begin
          regCount_55_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_55_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_55_1 <= newCountRefill_1;
        end else begin
          regCount_55_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_55_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_55_2 <= newCountRefill_2;
        end else begin
          regCount_55_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_55_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h37 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_55_3 <= newCountRefill_3;
        end else begin
          regCount_55_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_56_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_56_0 <= newCountRefill_0;
        end else begin
          regCount_56_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_56_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_56_1 <= newCountRefill_1;
        end else begin
          regCount_56_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_56_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_56_2 <= newCountRefill_2;
        end else begin
          regCount_56_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_56_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h38 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_56_3 <= newCountRefill_3;
        end else begin
          regCount_56_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_57_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_57_0 <= newCountRefill_0;
        end else begin
          regCount_57_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_57_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_57_1 <= newCountRefill_1;
        end else begin
          regCount_57_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_57_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_57_2 <= newCountRefill_2;
        end else begin
          regCount_57_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_57_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h39 == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_57_3 <= newCountRefill_3;
        end else begin
          regCount_57_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_58_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_58_0 <= newCountRefill_0;
        end else begin
          regCount_58_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_58_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_58_1 <= newCountRefill_1;
        end else begin
          regCount_58_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_58_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_58_2 <= newCountRefill_2;
        end else begin
          regCount_58_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_58_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3a == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_58_3 <= newCountRefill_3;
        end else begin
          regCount_58_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_59_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_59_0 <= newCountRefill_0;
        end else begin
          regCount_59_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_59_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_59_1 <= newCountRefill_1;
        end else begin
          regCount_59_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_59_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_59_2 <= newCountRefill_2;
        end else begin
          regCount_59_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_59_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3b == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_59_3 <= newCountRefill_3;
        end else begin
          regCount_59_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_60_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_60_0 <= newCountRefill_0;
        end else begin
          regCount_60_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_60_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_60_1 <= newCountRefill_1;
        end else begin
          regCount_60_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_60_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_60_2 <= newCountRefill_2;
        end else begin
          regCount_60_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_60_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3c == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_60_3 <= newCountRefill_3;
        end else begin
          regCount_60_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_61_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_61_0 <= newCountRefill_0;
        end else begin
          regCount_61_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_61_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_61_1 <= newCountRefill_1;
        end else begin
          regCount_61_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_61_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_61_2 <= newCountRefill_2;
        end else begin
          regCount_61_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_61_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3d == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_61_3 <= newCountRefill_3;
        end else begin
          regCount_61_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_62_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_62_0 <= newCountRefill_0;
        end else begin
          regCount_62_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_62_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_62_1 <= newCountRefill_1;
        end else begin
          regCount_62_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_62_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_62_2 <= newCountRefill_2;
        end else begin
          regCount_62_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_62_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3e == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_62_3 <= newCountRefill_3;
        end else begin
          regCount_62_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      regCount_63_0 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_63_0 <= newCountRefill_0;
        end else begin
          regCount_63_0 <= newCountHit_0;
        end
      end
    end
    if (reset) begin
      regCount_63_1 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_63_1 <= newCountRefill_1;
        end else begin
          regCount_63_1 <= newCountHit_1;
        end
      end
    end
    if (reset) begin
      regCount_63_2 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_63_2 <= newCountRefill_2;
        end else begin
          regCount_63_2 <= newCountHit_2;
        end
      end
    end
    if (reset) begin
      regCount_63_3 <= 2'h0;
    end else if (countUpdate) begin
      if (6'h3f == _WIRE_9[9:4]) begin
        if (memRespUpdate) begin
          regCount_63_3 <= newCountRefill_3;
        end else begin
          regCount_63_3 <= newCountHit_3;
        end
      end
    end
    if (reset) begin
      req_addr_r <= 32'h0;
    end else if (s1_valid) begin
      req_addr_r <= arbiter_io_out_bits_addr;
    end
    if (reset) begin
      s2_reg_valid <= 1'h0;
    end else if (~s2_stall) begin
      s2_reg_valid <= s1_valid;
    end
    if (reset) begin
      s2_reg_wdata <= 64'h0;
    end else if (~s2_stall) begin
      if (s1_valid) begin
        s2_reg_wdata <= s1_wdata;
      end else begin
        s2_reg_wdata <= 64'h0;
      end
    end
    if (reset) begin
      s2_reg_wen <= 1'h0;
    end else if (~s2_stall) begin
      s2_reg_wen <= _GEN_3;
    end
    if (reset) begin
      s2_reg_strb <= 8'h0;
    end else if (~s2_stall) begin
      if (s1_valid) begin
        s2_reg_strb <= s1_strb;
      end else begin
        s2_reg_strb <= 8'h0;
      end
    end
    if (reset) begin
      s2_reg_probe <= 1'h0;
    end else if (~s2_stall) begin
      s2_reg_probe <= _GEN_5;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  regCount_0_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  regCount_0_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  regCount_0_2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  regCount_0_3 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  regCount_1_0 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  regCount_1_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  regCount_1_2 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  regCount_1_3 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  regCount_2_0 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  regCount_2_1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  regCount_2_2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  regCount_2_3 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  regCount_3_0 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  regCount_3_1 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  regCount_3_2 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  regCount_3_3 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  regCount_4_0 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  regCount_4_1 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  regCount_4_2 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  regCount_4_3 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  regCount_5_0 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  regCount_5_1 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  regCount_5_2 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  regCount_5_3 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  regCount_6_0 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  regCount_6_1 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  regCount_6_2 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  regCount_6_3 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  regCount_7_0 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  regCount_7_1 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  regCount_7_2 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  regCount_7_3 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  regCount_8_0 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  regCount_8_1 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  regCount_8_2 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  regCount_8_3 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  regCount_9_0 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  regCount_9_1 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  regCount_9_2 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  regCount_9_3 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  regCount_10_0 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  regCount_10_1 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  regCount_10_2 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  regCount_10_3 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  regCount_11_0 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  regCount_11_1 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  regCount_11_2 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  regCount_11_3 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  regCount_12_0 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  regCount_12_1 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  regCount_12_2 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  regCount_12_3 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  regCount_13_0 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  regCount_13_1 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  regCount_13_2 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  regCount_13_3 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  regCount_14_0 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  regCount_14_1 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  regCount_14_2 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  regCount_14_3 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  regCount_15_0 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  regCount_15_1 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  regCount_15_2 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  regCount_15_3 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  regCount_16_0 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  regCount_16_1 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  regCount_16_2 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  regCount_16_3 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  regCount_17_0 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  regCount_17_1 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  regCount_17_2 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  regCount_17_3 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  regCount_18_0 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  regCount_18_1 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  regCount_18_2 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  regCount_18_3 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  regCount_19_0 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  regCount_19_1 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  regCount_19_2 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  regCount_19_3 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  regCount_20_0 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  regCount_20_1 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  regCount_20_2 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  regCount_20_3 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  regCount_21_0 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  regCount_21_1 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  regCount_21_2 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  regCount_21_3 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  regCount_22_0 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  regCount_22_1 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  regCount_22_2 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  regCount_22_3 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  regCount_23_0 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  regCount_23_1 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  regCount_23_2 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  regCount_23_3 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  regCount_24_0 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  regCount_24_1 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  regCount_24_2 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  regCount_24_3 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  regCount_25_0 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  regCount_25_1 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  regCount_25_2 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  regCount_25_3 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  regCount_26_0 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  regCount_26_1 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  regCount_26_2 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  regCount_26_3 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  regCount_27_0 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  regCount_27_1 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  regCount_27_2 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  regCount_27_3 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  regCount_28_0 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  regCount_28_1 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  regCount_28_2 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  regCount_28_3 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  regCount_29_0 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  regCount_29_1 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  regCount_29_2 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  regCount_29_3 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  regCount_30_0 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  regCount_30_1 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  regCount_30_2 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  regCount_30_3 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  regCount_31_0 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  regCount_31_1 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  regCount_31_2 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  regCount_31_3 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  regCount_32_0 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  regCount_32_1 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  regCount_32_2 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  regCount_32_3 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  regCount_33_0 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  regCount_33_1 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  regCount_33_2 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  regCount_33_3 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  regCount_34_0 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  regCount_34_1 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  regCount_34_2 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  regCount_34_3 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  regCount_35_0 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  regCount_35_1 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  regCount_35_2 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  regCount_35_3 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  regCount_36_0 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  regCount_36_1 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  regCount_36_2 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  regCount_36_3 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  regCount_37_0 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  regCount_37_1 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  regCount_37_2 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  regCount_37_3 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  regCount_38_0 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  regCount_38_1 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  regCount_38_2 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  regCount_38_3 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  regCount_39_0 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  regCount_39_1 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  regCount_39_2 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  regCount_39_3 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  regCount_40_0 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  regCount_40_1 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  regCount_40_2 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  regCount_40_3 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  regCount_41_0 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  regCount_41_1 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  regCount_41_2 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  regCount_41_3 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  regCount_42_0 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  regCount_42_1 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  regCount_42_2 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  regCount_42_3 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  regCount_43_0 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  regCount_43_1 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  regCount_43_2 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  regCount_43_3 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  regCount_44_0 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  regCount_44_1 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  regCount_44_2 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  regCount_44_3 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  regCount_45_0 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  regCount_45_1 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  regCount_45_2 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  regCount_45_3 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  regCount_46_0 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  regCount_46_1 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  regCount_46_2 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  regCount_46_3 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  regCount_47_0 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  regCount_47_1 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  regCount_47_2 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  regCount_47_3 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  regCount_48_0 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  regCount_48_1 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  regCount_48_2 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  regCount_48_3 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  regCount_49_0 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  regCount_49_1 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  regCount_49_2 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  regCount_49_3 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  regCount_50_0 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  regCount_50_1 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  regCount_50_2 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  regCount_50_3 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  regCount_51_0 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  regCount_51_1 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  regCount_51_2 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  regCount_51_3 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  regCount_52_0 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  regCount_52_1 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  regCount_52_2 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  regCount_52_3 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  regCount_53_0 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  regCount_53_1 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  regCount_53_2 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  regCount_53_3 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  regCount_54_0 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  regCount_54_1 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  regCount_54_2 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  regCount_54_3 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  regCount_55_0 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  regCount_55_1 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  regCount_55_2 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  regCount_55_3 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  regCount_56_0 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  regCount_56_1 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  regCount_56_2 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  regCount_56_3 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  regCount_57_0 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  regCount_57_1 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  regCount_57_2 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  regCount_57_3 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  regCount_58_0 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  regCount_58_1 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  regCount_58_2 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  regCount_58_3 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  regCount_59_0 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  regCount_59_1 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  regCount_59_2 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  regCount_59_3 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  regCount_60_0 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  regCount_60_1 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  regCount_60_2 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  regCount_60_3 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  regCount_61_0 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  regCount_61_1 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  regCount_61_2 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  regCount_61_3 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  regCount_62_0 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  regCount_62_1 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  regCount_62_2 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  regCount_62_3 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  regCount_63_0 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  regCount_63_1 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  regCount_63_2 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  regCount_63_3 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  req_addr_r = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  s2_reg_valid = _RAND_258[0:0];
  _RAND_259 = {2{`RANDOM}};
  s2_reg_wdata = _RAND_259[63:0];
  _RAND_260 = {1{`RANDOM}};
  s2_reg_wen = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  s2_reg_strb = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  s2_reg_probe = _RAND_262[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_CoreOverlay(
  input          clock,
  input          reset,
  input          io_imem_req_ready,
  output         io_imem_req_valid,
  output [31:0]  io_imem_req_bits_addr,
  output [127:0] io_imem_req_bits_wdata,
  output [2:0]   io_imem_req_bits_cmd,
  input          io_imem_resp_valid,
  input  [127:0] io_imem_resp_bits_rdata,
  input          io_dmem_req_ready,
  output         io_dmem_req_valid,
  output [31:0]  io_dmem_req_bits_addr,
  output [127:0] io_dmem_req_bits_wdata,
  output [2:0]   io_dmem_req_bits_cmd,
  input          io_dmem_resp_valid,
  input  [127:0] io_dmem_resp_bits_rdata,
  output         io_link_req_ready,
  input          io_link_req_valid,
  input  [31:0]  io_link_req_bits_addr,
  input  [127:0] io_link_req_bits_wdata,
  output         io_link_resp_valid,
  output [2:0]   io_link_resp_bits_cmd,
  output [127:0] io_link_resp_bits_rdata,
  input          io_immio_req_ready,
  output         io_immio_req_valid,
  output [31:0]  io_immio_req_bits_addr,
  output [1:0]   io_immio_req_bits_size,
  input          io_immio_resp_valid,
  input  [63:0]  io_immio_resp_bits_rdata,
  input          io_dmmio_req_ready,
  output         io_dmmio_req_valid,
  output [31:0]  io_dmmio_req_bits_addr,
  output [63:0]  io_dmmio_req_bits_wdata,
  output [1:0]   io_dmmio_req_bits_size,
  output [2:0]   io_dmmio_req_bits_cmd,
  input          io_dmmio_resp_valid,
  input  [63:0]  io_dmmio_resp_bits_rdata,
  input  [127:0] io_sram0_rdata,
  output         io_sram0_wen,
  output [5:0]   io_sram0_addr,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram1_rdata,
  output         io_sram1_wen,
  output [5:0]   io_sram1_addr,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram2_rdata,
  output         io_sram2_wen,
  output [5:0]   io_sram2_addr,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram3_rdata,
  output         io_sram3_wen,
  output [5:0]   io_sram3_addr,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram4_rdata,
  output         io_sram4_wen,
  output [5:0]   io_sram4_addr,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram5_rdata,
  output         io_sram5_wen,
  output [5:0]   io_sram5_addr,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram6_rdata,
  output         io_sram6_wen,
  output [5:0]   io_sram6_addr,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram7_rdata,
  output         io_sram7_wen,
  output [5:0]   io_sram7_addr,
  output [127:0] io_sram7_wdata
);
  wire  myCore_clock;
  wire  myCore_reset;
  wire  myCore_io_dmem_req_ready;
  wire  myCore_io_dmem_req_valid;
  wire [31:0] myCore_io_dmem_req_bits_addr;
  wire [63:0] myCore_io_dmem_req_bits_wdata;
  wire [1:0] myCore_io_dmem_req_bits_size;
  wire [2:0] myCore_io_dmem_req_bits_cmd;
  wire  myCore_io_dmem_resp_valid;
  wire [63:0] myCore_io_dmem_resp_bits_rdata;
  wire  myCore_io_imem_req_ready;
  wire [31:0] myCore_io_imem_req_bits_addr;
  wire  myCore_io_imem_resp_ready;
  wire  myCore_io_imem_resp_valid;
  wire [63:0] myCore_io_imem_resp_bits_rdata;
  wire  myCore_io_dmmio_req_ready;
  wire  myCore_io_dmmio_req_valid;
  wire [31:0] myCore_io_dmmio_req_bits_addr;
  wire [63:0] myCore_io_dmmio_req_bits_wdata;
  wire [1:0] myCore_io_dmmio_req_bits_size;
  wire [2:0] myCore_io_dmmio_req_bits_cmd;
  wire  myCore_io_dmmio_resp_valid;
  wire [63:0] myCore_io_dmmio_resp_bits_rdata;
  wire  myCore_flushICache;
  wire  iCache_clock;
  wire  iCache_reset;
  wire  iCache_io_in_req_ready;
  wire [31:0] iCache_io_in_req_bits_addr;
  wire  iCache_io_in_resp_ready;
  wire  iCache_io_in_resp_valid;
  wire [31:0] iCache_io_in_resp_bits_rdata;
  wire  iCache_io_out_req_ready;
  wire  iCache_io_out_req_valid;
  wire [31:0] iCache_io_out_req_bits_addr;
  wire [127:0] iCache_io_out_req_bits_wdata;
  wire [2:0] iCache_io_out_req_bits_cmd;
  wire  iCache_io_out_resp_ready;
  wire  iCache_io_out_resp_valid;
  wire [127:0] iCache_io_out_resp_bits_rdata;
  wire  iCache_io_mmio_req_ready;
  wire  iCache_io_mmio_req_valid;
  wire [31:0] iCache_io_mmio_req_bits_addr;
  wire [1:0] iCache_io_mmio_req_bits_size;
  wire  iCache_io_mmio_resp_ready;
  wire  iCache_io_mmio_resp_valid;
  wire [63:0] iCache_io_mmio_resp_bits_rdata;
  wire [127:0] iCache_io_dataArray_0_rdata;
  wire  iCache_io_dataArray_0_wen;
  wire [5:0] iCache_io_dataArray_0_addr;
  wire [127:0] iCache_io_dataArray_0_wdata;
  wire [127:0] iCache_io_dataArray_1_rdata;
  wire  iCache_io_dataArray_1_wen;
  wire [5:0] iCache_io_dataArray_1_addr;
  wire [127:0] iCache_io_dataArray_1_wdata;
  wire [127:0] iCache_io_dataArray_2_rdata;
  wire  iCache_io_dataArray_2_wen;
  wire [5:0] iCache_io_dataArray_2_addr;
  wire [127:0] iCache_io_dataArray_2_wdata;
  wire [127:0] iCache_io_dataArray_3_rdata;
  wire  iCache_io_dataArray_3_wen;
  wire [5:0] iCache_io_dataArray_3_addr;
  wire [127:0] iCache_io_dataArray_3_wdata;
  wire  iCache_difftestFENCEI;
  wire  dCache_clock;
  wire  dCache_reset;
  wire  dCache_io_in_req_ready;
  wire  dCache_io_in_req_valid;
  wire [31:0] dCache_io_in_req_bits_addr;
  wire [63:0] dCache_io_in_req_bits_wdata;
  wire [1:0] dCache_io_in_req_bits_size;
  wire [2:0] dCache_io_in_req_bits_cmd;
  wire  dCache_io_in_resp_valid;
  wire [63:0] dCache_io_in_resp_bits_rdata;
  wire  dCache_io_out_req_ready;
  wire  dCache_io_out_req_valid;
  wire [31:0] dCache_io_out_req_bits_addr;
  wire [127:0] dCache_io_out_req_bits_wdata;
  wire [2:0] dCache_io_out_req_bits_cmd;
  wire  dCache_io_out_resp_ready;
  wire  dCache_io_out_resp_valid;
  wire [127:0] dCache_io_out_resp_bits_rdata;
  wire  dCache_io_link_req_ready;
  wire  dCache_io_link_req_valid;
  wire [31:0] dCache_io_link_req_bits_addr;
  wire [127:0] dCache_io_link_req_bits_wdata;
  wire  dCache_io_link_resp_valid;
  wire [2:0] dCache_io_link_resp_bits_cmd;
  wire [127:0] dCache_io_link_resp_bits_rdata;
  wire [127:0] dCache_io_dataArray_0_rdata;
  wire  dCache_io_dataArray_0_wen;
  wire [5:0] dCache_io_dataArray_0_addr;
  wire [127:0] dCache_io_dataArray_0_wdata;
  wire [127:0] dCache_io_dataArray_1_rdata;
  wire  dCache_io_dataArray_1_wen;
  wire [5:0] dCache_io_dataArray_1_addr;
  wire [127:0] dCache_io_dataArray_1_wdata;
  wire [127:0] dCache_io_dataArray_2_rdata;
  wire  dCache_io_dataArray_2_wen;
  wire [5:0] dCache_io_dataArray_2_addr;
  wire [127:0] dCache_io_dataArray_2_wdata;
  wire [127:0] dCache_io_dataArray_3_rdata;
  wire  dCache_io_dataArray_3_wen;
  wire [5:0] dCache_io_dataArray_3_addr;
  wire [127:0] dCache_io_dataArray_3_wdata;
  ysyx_040656_MyCore myCore (
    .clock(myCore_clock),
    .reset(myCore_reset),
    .io_dmem_req_ready(myCore_io_dmem_req_ready),
    .io_dmem_req_valid(myCore_io_dmem_req_valid),
    .io_dmem_req_bits_addr(myCore_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(myCore_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_size(myCore_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(myCore_io_dmem_req_bits_cmd),
    .io_dmem_resp_valid(myCore_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(myCore_io_dmem_resp_bits_rdata),
    .io_imem_req_ready(myCore_io_imem_req_ready),
    .io_imem_req_bits_addr(myCore_io_imem_req_bits_addr),
    .io_imem_resp_ready(myCore_io_imem_resp_ready),
    .io_imem_resp_valid(myCore_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(myCore_io_imem_resp_bits_rdata),
    .io_dmmio_req_ready(myCore_io_dmmio_req_ready),
    .io_dmmio_req_valid(myCore_io_dmmio_req_valid),
    .io_dmmio_req_bits_addr(myCore_io_dmmio_req_bits_addr),
    .io_dmmio_req_bits_wdata(myCore_io_dmmio_req_bits_wdata),
    .io_dmmio_req_bits_size(myCore_io_dmmio_req_bits_size),
    .io_dmmio_req_bits_cmd(myCore_io_dmmio_req_bits_cmd),
    .io_dmmio_resp_valid(myCore_io_dmmio_resp_valid),
    .io_dmmio_resp_bits_rdata(myCore_io_dmmio_resp_bits_rdata),
    .flushICache(myCore_flushICache)
  );
  ysyx_040656_ICache iCache (
    .clock(iCache_clock),
    .reset(iCache_reset),
    .io_in_req_ready(iCache_io_in_req_ready),
    .io_in_req_bits_addr(iCache_io_in_req_bits_addr),
    .io_in_resp_ready(iCache_io_in_resp_ready),
    .io_in_resp_valid(iCache_io_in_resp_valid),
    .io_in_resp_bits_rdata(iCache_io_in_resp_bits_rdata),
    .io_out_req_ready(iCache_io_out_req_ready),
    .io_out_req_valid(iCache_io_out_req_valid),
    .io_out_req_bits_addr(iCache_io_out_req_bits_addr),
    .io_out_req_bits_wdata(iCache_io_out_req_bits_wdata),
    .io_out_req_bits_cmd(iCache_io_out_req_bits_cmd),
    .io_out_resp_ready(iCache_io_out_resp_ready),
    .io_out_resp_valid(iCache_io_out_resp_valid),
    .io_out_resp_bits_rdata(iCache_io_out_resp_bits_rdata),
    .io_mmio_req_ready(iCache_io_mmio_req_ready),
    .io_mmio_req_valid(iCache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(iCache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(iCache_io_mmio_req_bits_size),
    .io_mmio_resp_ready(iCache_io_mmio_resp_ready),
    .io_mmio_resp_valid(iCache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(iCache_io_mmio_resp_bits_rdata),
    .io_dataArray_0_rdata(iCache_io_dataArray_0_rdata),
    .io_dataArray_0_wen(iCache_io_dataArray_0_wen),
    .io_dataArray_0_addr(iCache_io_dataArray_0_addr),
    .io_dataArray_0_wdata(iCache_io_dataArray_0_wdata),
    .io_dataArray_1_rdata(iCache_io_dataArray_1_rdata),
    .io_dataArray_1_wen(iCache_io_dataArray_1_wen),
    .io_dataArray_1_addr(iCache_io_dataArray_1_addr),
    .io_dataArray_1_wdata(iCache_io_dataArray_1_wdata),
    .io_dataArray_2_rdata(iCache_io_dataArray_2_rdata),
    .io_dataArray_2_wen(iCache_io_dataArray_2_wen),
    .io_dataArray_2_addr(iCache_io_dataArray_2_addr),
    .io_dataArray_2_wdata(iCache_io_dataArray_2_wdata),
    .io_dataArray_3_rdata(iCache_io_dataArray_3_rdata),
    .io_dataArray_3_wen(iCache_io_dataArray_3_wen),
    .io_dataArray_3_addr(iCache_io_dataArray_3_addr),
    .io_dataArray_3_wdata(iCache_io_dataArray_3_wdata),
    .difftestFENCEI(iCache_difftestFENCEI)
  );
  ysyx_040656_DCache dCache (
    .clock(dCache_clock),
    .reset(dCache_reset),
    .io_in_req_ready(dCache_io_in_req_ready),
    .io_in_req_valid(dCache_io_in_req_valid),
    .io_in_req_bits_addr(dCache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(dCache_io_in_req_bits_wdata),
    .io_in_req_bits_size(dCache_io_in_req_bits_size),
    .io_in_req_bits_cmd(dCache_io_in_req_bits_cmd),
    .io_in_resp_valid(dCache_io_in_resp_valid),
    .io_in_resp_bits_rdata(dCache_io_in_resp_bits_rdata),
    .io_out_req_ready(dCache_io_out_req_ready),
    .io_out_req_valid(dCache_io_out_req_valid),
    .io_out_req_bits_addr(dCache_io_out_req_bits_addr),
    .io_out_req_bits_wdata(dCache_io_out_req_bits_wdata),
    .io_out_req_bits_cmd(dCache_io_out_req_bits_cmd),
    .io_out_resp_ready(dCache_io_out_resp_ready),
    .io_out_resp_valid(dCache_io_out_resp_valid),
    .io_out_resp_bits_rdata(dCache_io_out_resp_bits_rdata),
    .io_link_req_ready(dCache_io_link_req_ready),
    .io_link_req_valid(dCache_io_link_req_valid),
    .io_link_req_bits_addr(dCache_io_link_req_bits_addr),
    .io_link_req_bits_wdata(dCache_io_link_req_bits_wdata),
    .io_link_resp_valid(dCache_io_link_resp_valid),
    .io_link_resp_bits_cmd(dCache_io_link_resp_bits_cmd),
    .io_link_resp_bits_rdata(dCache_io_link_resp_bits_rdata),
    .io_dataArray_0_rdata(dCache_io_dataArray_0_rdata),
    .io_dataArray_0_wen(dCache_io_dataArray_0_wen),
    .io_dataArray_0_addr(dCache_io_dataArray_0_addr),
    .io_dataArray_0_wdata(dCache_io_dataArray_0_wdata),
    .io_dataArray_1_rdata(dCache_io_dataArray_1_rdata),
    .io_dataArray_1_wen(dCache_io_dataArray_1_wen),
    .io_dataArray_1_addr(dCache_io_dataArray_1_addr),
    .io_dataArray_1_wdata(dCache_io_dataArray_1_wdata),
    .io_dataArray_2_rdata(dCache_io_dataArray_2_rdata),
    .io_dataArray_2_wen(dCache_io_dataArray_2_wen),
    .io_dataArray_2_addr(dCache_io_dataArray_2_addr),
    .io_dataArray_2_wdata(dCache_io_dataArray_2_wdata),
    .io_dataArray_3_rdata(dCache_io_dataArray_3_rdata),
    .io_dataArray_3_wen(dCache_io_dataArray_3_wen),
    .io_dataArray_3_addr(dCache_io_dataArray_3_addr),
    .io_dataArray_3_wdata(dCache_io_dataArray_3_wdata)
  );
  assign io_imem_req_valid = iCache_io_out_req_valid;
  assign io_imem_req_bits_addr = iCache_io_out_req_bits_addr;
  assign io_imem_req_bits_wdata = iCache_io_out_req_bits_wdata;
  assign io_imem_req_bits_cmd = iCache_io_out_req_bits_cmd;
  assign io_dmem_req_valid = dCache_io_out_req_valid;
  assign io_dmem_req_bits_addr = dCache_io_out_req_bits_addr;
  assign io_dmem_req_bits_wdata = dCache_io_out_req_bits_wdata;
  assign io_dmem_req_bits_cmd = dCache_io_out_req_bits_cmd;
  assign io_link_req_ready = dCache_io_link_req_ready;
  assign io_link_resp_valid = dCache_io_link_resp_valid;
  assign io_link_resp_bits_cmd = dCache_io_link_resp_bits_cmd;
  assign io_link_resp_bits_rdata = dCache_io_link_resp_bits_rdata;
  assign io_immio_req_valid = iCache_io_mmio_req_valid;
  assign io_immio_req_bits_addr = iCache_io_mmio_req_bits_addr;
  assign io_immio_req_bits_size = iCache_io_mmio_req_bits_size;
  assign io_dmmio_req_valid = myCore_io_dmmio_req_valid;
  assign io_dmmio_req_bits_addr = myCore_io_dmmio_req_bits_addr;
  assign io_dmmio_req_bits_wdata = myCore_io_dmmio_req_bits_wdata;
  assign io_dmmio_req_bits_size = myCore_io_dmmio_req_bits_size;
  assign io_dmmio_req_bits_cmd = myCore_io_dmmio_req_bits_cmd;
  assign io_sram0_wen = dCache_io_dataArray_0_wen;
  assign io_sram0_addr = dCache_io_dataArray_0_addr;
  assign io_sram0_wdata = dCache_io_dataArray_0_wdata;
  assign io_sram1_wen = dCache_io_dataArray_1_wen;
  assign io_sram1_addr = dCache_io_dataArray_1_addr;
  assign io_sram1_wdata = dCache_io_dataArray_1_wdata;
  assign io_sram2_wen = dCache_io_dataArray_2_wen;
  assign io_sram2_addr = dCache_io_dataArray_2_addr;
  assign io_sram2_wdata = dCache_io_dataArray_2_wdata;
  assign io_sram3_wen = dCache_io_dataArray_3_wen;
  assign io_sram3_addr = dCache_io_dataArray_3_addr;
  assign io_sram3_wdata = dCache_io_dataArray_3_wdata;
  assign io_sram4_wen = iCache_io_dataArray_0_wen;
  assign io_sram4_addr = iCache_io_dataArray_0_addr;
  assign io_sram4_wdata = iCache_io_dataArray_0_wdata;
  assign io_sram5_wen = iCache_io_dataArray_1_wen;
  assign io_sram5_addr = iCache_io_dataArray_1_addr;
  assign io_sram5_wdata = iCache_io_dataArray_1_wdata;
  assign io_sram6_wen = iCache_io_dataArray_2_wen;
  assign io_sram6_addr = iCache_io_dataArray_2_addr;
  assign io_sram6_wdata = iCache_io_dataArray_2_wdata;
  assign io_sram7_wen = iCache_io_dataArray_3_wen;
  assign io_sram7_addr = iCache_io_dataArray_3_addr;
  assign io_sram7_wdata = iCache_io_dataArray_3_wdata;
  assign myCore_clock = clock;
  assign myCore_reset = reset;
  assign myCore_io_dmem_req_ready = dCache_io_in_req_ready;
  assign myCore_io_dmem_resp_valid = dCache_io_in_resp_valid;
  assign myCore_io_dmem_resp_bits_rdata = dCache_io_in_resp_bits_rdata;
  assign myCore_io_imem_req_ready = iCache_io_in_req_ready;
  assign myCore_io_imem_resp_valid = iCache_io_in_resp_valid;
  assign myCore_io_imem_resp_bits_rdata = {{32'd0}, iCache_io_in_resp_bits_rdata};
  assign myCore_io_dmmio_req_ready = io_dmmio_req_ready;
  assign myCore_io_dmmio_resp_valid = io_dmmio_resp_valid;
  assign myCore_io_dmmio_resp_bits_rdata = io_dmmio_resp_bits_rdata;
  assign iCache_clock = clock;
  assign iCache_reset = reset;
  assign iCache_io_in_req_bits_addr = myCore_io_imem_req_bits_addr;
  assign iCache_io_in_resp_ready = myCore_io_imem_resp_ready;
  assign iCache_io_out_req_ready = io_imem_req_ready;
  assign iCache_io_out_resp_valid = io_imem_resp_valid;
  assign iCache_io_out_resp_bits_rdata = io_imem_resp_bits_rdata;
  assign iCache_io_mmio_req_ready = io_immio_req_ready;
  assign iCache_io_mmio_resp_valid = io_immio_resp_valid;
  assign iCache_io_mmio_resp_bits_rdata = io_immio_resp_bits_rdata;
  assign iCache_io_dataArray_0_rdata = io_sram4_rdata;
  assign iCache_io_dataArray_1_rdata = io_sram5_rdata;
  assign iCache_io_dataArray_2_rdata = io_sram6_rdata;
  assign iCache_io_dataArray_3_rdata = io_sram7_rdata;
  assign iCache_difftestFENCEI = myCore_flushICache;
  assign dCache_clock = clock;
  assign dCache_reset = reset;
  assign dCache_io_in_req_valid = myCore_io_dmem_req_valid;
  assign dCache_io_in_req_bits_addr = myCore_io_dmem_req_bits_addr;
  assign dCache_io_in_req_bits_wdata = myCore_io_dmem_req_bits_wdata;
  assign dCache_io_in_req_bits_size = myCore_io_dmem_req_bits_size;
  assign dCache_io_in_req_bits_cmd = myCore_io_dmem_req_bits_cmd;
  assign dCache_io_out_req_ready = io_dmem_req_ready;
  assign dCache_io_out_resp_valid = io_dmem_resp_valid;
  assign dCache_io_out_resp_bits_rdata = io_dmem_resp_bits_rdata;
  assign dCache_io_link_req_valid = io_link_req_valid;
  assign dCache_io_link_req_bits_addr = io_link_req_bits_addr;
  assign dCache_io_link_req_bits_wdata = io_link_req_bits_wdata;
  assign dCache_io_dataArray_0_rdata = io_sram0_rdata;
  assign dCache_io_dataArray_1_rdata = io_sram1_rdata;
  assign dCache_io_dataArray_2_rdata = io_sram2_rdata;
  assign dCache_io_dataArray_3_rdata = io_sram3_rdata;
endmodule
module ysyx_040656_XConnect(
  input          clock,
  input          reset,
  output         io_in_req_ready,
  input          io_in_req_valid,
  input  [31:0]  io_in_req_bits_addr,
  input  [127:0] io_in_req_bits_wdata,
  input  [2:0]   io_in_req_bits_cmd,
  output         io_in_resp_valid,
  output [127:0] io_in_resp_bits_rdata,
  input          io_out_mem_req_ready,
  output         io_out_mem_req_valid,
  output [31:0]  io_out_mem_req_bits_addr,
  output [127:0] io_out_mem_req_bits_wdata,
  output [2:0]   io_out_mem_req_bits_cmd,
  output         io_out_mem_resp_ready,
  input          io_out_mem_resp_valid,
  input  [2:0]   io_out_mem_resp_bits_cmd,
  input  [127:0] io_out_mem_resp_bits_rdata,
  input          io_out_link_req_ready,
  output         io_out_link_req_valid,
  output [31:0]  io_out_link_req_bits_addr,
  output [127:0] io_out_link_req_bits_wdata,
  output         io_out_link_resp_ready,
  input          io_out_link_resp_valid,
  input  [2:0]   io_out_link_resp_bits_cmd,
  input  [127:0] io_out_link_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif
  reg [2:0] state;
  wire  running = state != 3'h0;
  wire  _requestBuffer_T = ~running;
  wire  _requestBuffer_T_3 = io_in_req_bits_cmd == 3'h0 | io_in_req_bits_cmd == 3'h3;
  wire  _requestBuffer_T_4 = ~running & _requestBuffer_T_3;
  reg [31:0] requestBuffer_addr;
  reg [127:0] requestBuffer_wdata;
  reg [2:0] requestBuffer_cmd;
  wire  _T_2 = io_in_req_bits_cmd == 3'h1 | io_in_req_bits_cmd == 3'h4;
  wire  _io_out_mem_req_valid_T_1 = io_in_req_valid & _requestBuffer_T;
  wire  _GEN_4 = _requestBuffer_T_3 & _io_out_mem_req_valid_T_1;
  wire  _GEN_5 = _requestBuffer_T_3 & (io_out_link_req_ready & _requestBuffer_T);
  wire  _GEN_6 = _T_2 & (io_in_req_valid & _requestBuffer_T);
  reg [127:0] respBuffer_rdata;
  reg  respBufferValid;
  wire  _T_7 = io_in_req_ready & io_in_req_valid;
  wire [2:0] _GEN_9 = _T_2 ? 3'h5 : state;
  wire  _T_15 = io_out_link_resp_ready & io_out_link_resp_valid;
  wire  _state_T = io_out_link_resp_bits_cmd == 3'h5;
  wire [2:0] _state_T_1 = _state_T ? 3'h2 : 3'h3;
  wire  _T_18 = io_out_link_resp_bits_cmd == 3'h3;
  wire [127:0] _GEN_14 = _T_15 & _T_18 ? io_out_link_resp_bits_rdata : respBuffer_rdata;
  wire  _GEN_15 = _T_15 & _T_18 | respBufferValid;
  wire [2:0] _GEN_16 = _T_15 & _T_18 ? 3'h0 : state;
  wire  _T_21 = io_out_mem_req_ready & io_out_mem_req_valid;
  wire [2:0] _GEN_17 = _T_21 ? 3'h4 : state;
  wire  _T_23 = io_out_mem_resp_ready & io_out_mem_resp_valid;
  wire  _T_24 = io_out_mem_resp_bits_cmd == 3'h3;
  wire [127:0] _GEN_19 = _T_23 & _T_24 ? io_out_mem_resp_bits_rdata : respBuffer_rdata;
  wire  _GEN_20 = _T_23 & _T_24 | respBufferValid;
  wire [2:0] _GEN_21 = _T_23 & _T_24 ? 3'h0 : state;
  wire [2:0] _GEN_22 = _T_23 ? 3'h0 : state;
  wire [2:0] _GEN_23 = 3'h5 == state ? _GEN_22 : state;
  wire [127:0] _GEN_25 = 3'h4 == state ? _GEN_19 : respBuffer_rdata;
  wire  _GEN_26 = 3'h4 == state ? _GEN_20 : respBufferValid;
  wire [2:0] _GEN_27 = 3'h4 == state ? _GEN_21 : _GEN_23;
  wire [31:0] _GEN_28 = 3'h3 == state ? requestBuffer_addr : io_in_req_bits_addr;
  wire [127:0] _GEN_29 = 3'h3 == state ? requestBuffer_wdata : io_in_req_bits_wdata;
  wire [2:0] _GEN_31 = 3'h3 == state ? requestBuffer_cmd : io_in_req_bits_cmd;
  wire  _GEN_32 = 3'h3 == state | _GEN_6;
  wire [2:0] _GEN_33 = 3'h3 == state ? _GEN_17 : _GEN_27;
  wire [127:0] _GEN_35 = 3'h3 == state ? respBuffer_rdata : _GEN_25;
  wire  _GEN_36 = 3'h3 == state ? respBufferValid : _GEN_26;
  wire [31:0] _GEN_41 = 3'h2 == state ? io_in_req_bits_addr : _GEN_28;
  wire [127:0] _GEN_42 = 3'h2 == state ? io_in_req_bits_wdata : _GEN_29;
  wire [2:0] _GEN_44 = 3'h2 == state ? io_in_req_bits_cmd : _GEN_31;
  wire  _GEN_45 = 3'h2 == state ? _GEN_6 : _GEN_32;
  wire [31:0] _GEN_50 = 3'h1 == state ? io_in_req_bits_addr : _GEN_41;
  wire [127:0] _GEN_51 = 3'h1 == state ? io_in_req_bits_wdata : _GEN_42;
  wire [2:0] _GEN_53 = 3'h1 == state ? io_in_req_bits_cmd : _GEN_44;
  wire  _GEN_54 = 3'h1 == state ? _GEN_6 : _GEN_45;
  assign io_in_req_ready = _T_2 ? io_out_mem_req_ready & _requestBuffer_T : _GEN_5;
  assign io_in_resp_valid = respBufferValid;
  assign io_in_resp_bits_rdata = respBuffer_rdata;
  assign io_out_mem_req_valid = 3'h0 == state ? _GEN_6 : _GEN_54;
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_50;
  assign io_out_mem_req_bits_wdata = 3'h0 == state ? io_in_req_bits_wdata : _GEN_51;
  assign io_out_mem_req_bits_cmd = 3'h0 == state ? io_in_req_bits_cmd : _GEN_53;
  assign io_out_mem_resp_ready = 1'h1;
  assign io_out_link_req_valid = _T_2 ? 1'h0 : _GEN_4;
  assign io_out_link_req_bits_addr = io_in_req_bits_addr;
  assign io_out_link_req_bits_wdata = io_in_req_bits_wdata;
  assign io_out_link_resp_ready = 1'h1;
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (3'h0 == state) begin
      if (_T_7) begin
        if (_requestBuffer_T_3) begin
          state <= 3'h1;
        end else begin
          state <= _GEN_9;
        end
      end
    end else if (3'h1 == state) begin
      if (_T_15) begin
        state <= _state_T_1;
      end
    end else if (3'h2 == state) begin
      state <= _GEN_16;
    end else begin
      state <= _GEN_33;
    end
    if (_requestBuffer_T_4) begin
      requestBuffer_addr <= io_in_req_bits_addr;
    end
    if (_requestBuffer_T_4) begin
      requestBuffer_wdata <= io_in_req_bits_wdata;
    end
    if (_requestBuffer_T_4) begin
      requestBuffer_cmd <= io_in_req_bits_cmd;
    end
    if (reset) begin
      respBuffer_rdata <= 128'h0;
    end else if (!(3'h0 == state)) begin
      if (!(3'h1 == state)) begin
        if (3'h2 == state) begin
          respBuffer_rdata <= _GEN_14;
        end else begin
          respBuffer_rdata <= _GEN_35;
        end
      end
    end
    if (reset) begin
      respBufferValid <= 1'h0;
    end else if (3'h0 == state) begin
      respBufferValid <= 1'h0;
    end else if (!(3'h1 == state)) begin
      if (3'h2 == state) begin
        respBufferValid <= _GEN_15;
      end else begin
        respBufferValid <= _GEN_36;
      end
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  requestBuffer_addr = _RAND_1[31:0];
  _RAND_2 = {4{`RANDOM}};
  requestBuffer_wdata = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  requestBuffer_cmd = _RAND_3[2:0];
  _RAND_4 = {4{`RANDOM}};
  respBuffer_rdata = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  respBufferValid = _RAND_5[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_AXI4CLINT(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [7:0]  io_in_w_bits_strb,
  input  [63:0] io_in_w_bits_data,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif
  wire [7:0] _fullMask_T_9 = io_in_w_bits_strb[0] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_11 = io_in_w_bits_strb[1] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_13 = io_in_w_bits_strb[2] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_15 = io_in_w_bits_strb[3] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_17 = io_in_w_bits_strb[4] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_19 = io_in_w_bits_strb[5] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_21 = io_in_w_bits_strb[6] ? 8'hff : 8'h0;
  wire [7:0] _fullMask_T_23 = io_in_w_bits_strb[7] ? 8'hff : 8'h0;
  wire [63:0] fullMask = {_fullMask_T_23,_fullMask_T_21,_fullMask_T_19,_fullMask_T_17,_fullMask_T_15,_fullMask_T_13,
    _fullMask_T_11,_fullMask_T_9};
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid;
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid;
  reg  r_busy;
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy;
  wire  _GEN_1 = _r_busy_T | _GEN_0;
  reg  ren_REG;
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy);
  reg  io_in_r_valid_r;
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r;
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2;
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid;
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid;
  reg  w_busy;
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy;
  wire  _GEN_5 = _w_busy_T | _GEN_4;
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid;
  reg  io_in_b_valid_r;
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r;
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6;
  reg [63:0] msip;
  reg [63:0] mtime;
  reg [63:0] mtimecmp;
  reg [15:0] freq;
  reg [15:0] inc;
  reg [15:0] cnt;
  wire [15:0] nextCnt = cnt + 16'h1;
  wire  tick = nextCnt == freq;
  wire [63:0] _GEN_29 = {{48'd0}, inc};
  wire [63:0] _mtime_T_1 = mtime + _GEN_29;
  wire [63:0] _GEN_8 = tick ? _mtime_T_1 : mtime;
  wire [15:0] reg_raddr = io_in_ar_bits_addr[15:0];
  wire [15:0] reg_wadrr = io_in_aw_bits_addr[15:0];
  wire  _io_in_r_bits_data_T = reg_raddr == 16'h0;
  wire  _io_in_r_bits_data_T_1 = reg_raddr == 16'h4000;
  wire  _io_in_r_bits_data_T_2 = reg_raddr == 16'h8000;
  wire  _io_in_r_bits_data_T_3 = reg_raddr == 16'h8008;
  wire  _io_in_r_bits_data_T_4 = reg_raddr == 16'hbff8;
  wire [63:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_4 ? mtime : 64'h0;
  wire [63:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_3 ? {{48'd0}, inc} : _io_in_r_bits_data_T_5;
  wire [63:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_2 ? {{48'd0}, freq} : _io_in_r_bits_data_T_6;
  wire [63:0] _io_in_r_bits_data_T_8 = _io_in_r_bits_data_T_1 ? mtimecmp : _io_in_r_bits_data_T_7;
  wire [63:0] _msip_T_25 = io_in_w_bits_data & fullMask;
  wire [63:0] _msip_T_26 = ~fullMask;
  wire [63:0] _msip_T_27 = msip & _msip_T_26;
  wire [63:0] _msip_T_28 = _msip_T_25 | _msip_T_27;
  wire [63:0] _mtimecmp_T_27 = mtimecmp & _msip_T_26;
  wire [63:0] _mtimecmp_T_28 = _msip_T_25 | _mtimecmp_T_27;
  wire [63:0] _GEN_30 = {{48'd0}, freq};
  wire [63:0] _freq_T_27 = _GEN_30 & _msip_T_26;
  wire [63:0] _freq_T_28 = _msip_T_25 | _freq_T_27;
  wire [63:0] _inc_T_27 = _GEN_29 & _msip_T_26;
  wire [63:0] _inc_T_28 = _msip_T_25 | _inc_T_27;
  wire [63:0] _mtime_T_29 = mtime & _msip_T_26;
  wire [63:0] _mtime_T_30 = _msip_T_25 | _mtime_T_29;
  wire [63:0] _GEN_9 = reg_wadrr == 16'hbff8 ? _mtime_T_30 : _GEN_8;
  wire [63:0] _GEN_10 = reg_wadrr == 16'h8008 ? _inc_T_28 : {{48'd0}, inc};
  wire [63:0] _GEN_11 = reg_wadrr == 16'h8008 ? _GEN_8 : _GEN_9;
  wire [63:0] _GEN_12 = reg_wadrr == 16'h8000 ? _freq_T_28 : {{48'd0}, freq};
  wire [63:0] _GEN_13 = reg_wadrr == 16'h8000 ? {{48'd0}, inc} : _GEN_10;
  wire [63:0] _GEN_14 = reg_wadrr == 16'h8000 ? _GEN_8 : _GEN_11;
  wire [63:0] _GEN_16 = reg_wadrr == 16'h4000 ? {{48'd0}, freq} : _GEN_12;
  wire [63:0] _GEN_17 = reg_wadrr == 16'h4000 ? {{48'd0}, inc} : _GEN_13;
  wire [63:0] _GEN_21 = reg_wadrr == 16'h0 ? {{48'd0}, freq} : _GEN_16;
  wire [63:0] _GEN_22 = reg_wadrr == 16'h0 ? {{48'd0}, inc} : _GEN_17;
  wire [63:0] _GEN_26 = _io_in_b_valid_T ? _GEN_21 : {{48'd0}, freq};
  wire [63:0] _GEN_27 = _io_in_b_valid_T ? _GEN_22 : {{48'd0}, inc};
  wire [63:0] _GEN_32 = reset ? 64'ha : _GEN_26;
  wire [63:0] _GEN_33 = reset ? 64'h1 : _GEN_27;
  assign io_in_aw_ready = ~w_busy;
  assign io_in_w_ready = io_in_aw_valid | w_busy;
  assign io_in_b_valid = io_in_b_valid_r;
  assign io_in_ar_ready = io_in_r_ready | ~r_busy;
  assign io_in_r_valid = io_in_r_valid_r;
  assign io_in_r_bits_data = _io_in_r_bits_data_T ? msip : _io_in_r_bits_data_T_8;
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren_REG <= 1'h0;
    end else begin
      ren_REG <= _r_busy_T;
    end
    if (reset) begin
      io_in_r_valid_r <= 1'h0;
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      io_in_b_valid_r <= 1'h0;
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin
      msip <= 64'h0;
    end else if (_io_in_b_valid_T) begin
      if (reg_wadrr == 16'h0) begin
        msip <= _msip_T_28;
      end
    end
    if (reset) begin
      mtime <= 64'h0;
    end else if (_io_in_b_valid_T) begin
      if (reg_wadrr == 16'h0) begin
        mtime <= _GEN_8;
      end else if (reg_wadrr == 16'h4000) begin
        mtime <= _GEN_8;
      end else begin
        mtime <= _GEN_14;
      end
    end else begin
      mtime <= _GEN_8;
    end
    if (reset) begin
      mtimecmp <= 64'h0;
    end else if (_io_in_b_valid_T) begin
      if (!(reg_wadrr == 16'h0)) begin
        if (reg_wadrr == 16'h4000) begin
          mtimecmp <= _mtimecmp_T_28;
        end
      end
    end
    freq <= _GEN_32[15:0];
    inc <= _GEN_33[15:0];
    if (reset) begin
      cnt <= 16'h0;
    end else if (nextCnt < freq) begin
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  msip = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtime = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mtimecmp = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_Arbiter_1(
  output       io_in_0_ready,
  input        io_in_0_valid,
  output       io_in_1_ready,
  input        io_in_1_valid,
  output       io_in_2_ready,
  input        io_in_2_valid,
  output       io_in_3_ready,
  input        io_in_3_valid,
  output       io_in_4_ready,
  input        io_in_4_valid,
  output       io_in_5_ready,
  input        io_out_ready,
  output [2:0] io_chosen
);
  wire [2:0] _GEN_0 = io_in_4_valid ? 3'h4 : 3'h5;
  wire [2:0] _GEN_6 = io_in_3_valid ? 3'h3 : _GEN_0;
  wire [2:0] _GEN_12 = io_in_2_valid ? 3'h2 : _GEN_6;
  wire [2:0] _GEN_18 = io_in_1_valid ? 3'h1 : _GEN_12;
  wire  grant_1 = ~io_in_0_valid;
  wire  grant_2 = ~(io_in_0_valid | io_in_1_valid);
  wire  grant_3 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid);
  wire  grant_4 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid);
  wire  grant_5 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid);
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = grant_1 & io_out_ready;
  assign io_in_2_ready = grant_2 & io_out_ready;
  assign io_in_3_ready = grant_3 & io_out_ready;
  assign io_in_4_ready = grant_4 & io_out_ready;
  assign io_in_5_ready = grant_5 & io_out_ready;
  assign io_chosen = io_in_0_valid ? 3'h0 : _GEN_18;
endmodule
module ysyx_040656_AXI4XBar_Nto1(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [31:0] io_in_0_aw_bits_addr,
  input  [2:0]  io_in_0_aw_bits_size,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [31:0] io_in_0_ar_bits_addr,
  input  [2:0]  io_in_0_ar_bits_size,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [63:0] io_in_0_r_bits_data,
  output        io_in_0_r_bits_last,
  output        io_in_1_aw_ready,
  input         io_in_1_aw_valid,
  input  [31:0] io_in_1_aw_bits_addr,
  input  [2:0]  io_in_1_aw_bits_size,
  output        io_in_1_w_ready,
  input         io_in_1_w_valid,
  input  [63:0] io_in_1_w_bits_data,
  input         io_in_1_w_bits_last,
  input         io_in_1_b_ready,
  output        io_in_1_b_valid,
  output        io_in_1_ar_ready,
  input         io_in_1_ar_valid,
  input  [31:0] io_in_1_ar_bits_addr,
  input  [2:0]  io_in_1_ar_bits_size,
  input         io_in_1_r_ready,
  output        io_in_1_r_valid,
  output [63:0] io_in_1_r_bits_data,
  output        io_in_1_r_bits_last,
  output        io_in_2_aw_ready,
  input         io_in_2_aw_valid,
  input  [31:0] io_in_2_aw_bits_addr,
  input  [3:0]  io_in_2_aw_bits_id,
  input  [7:0]  io_in_2_aw_bits_len,
  input  [2:0]  io_in_2_aw_bits_size,
  input  [1:0]  io_in_2_aw_bits_burst,
  output        io_in_2_w_ready,
  input         io_in_2_w_valid,
  input  [7:0]  io_in_2_w_bits_strb,
  input  [63:0] io_in_2_w_bits_data,
  input         io_in_2_b_ready,
  output        io_in_2_b_valid,
  output        io_in_2_ar_ready,
  input         io_in_2_ar_valid,
  input  [31:0] io_in_2_ar_bits_addr,
  input  [2:0]  io_in_2_ar_bits_size,
  input         io_in_2_r_ready,
  output        io_in_2_r_valid,
  output [63:0] io_in_2_r_bits_data,
  output        io_in_2_r_bits_last,
  output        io_in_3_aw_ready,
  input         io_in_3_aw_valid,
  input  [31:0] io_in_3_aw_bits_addr,
  input  [3:0]  io_in_3_aw_bits_id,
  input  [7:0]  io_in_3_aw_bits_len,
  input  [2:0]  io_in_3_aw_bits_size,
  input  [1:0]  io_in_3_aw_bits_burst,
  output        io_in_3_w_ready,
  input         io_in_3_w_valid,
  input  [7:0]  io_in_3_w_bits_strb,
  input  [63:0] io_in_3_w_bits_data,
  input         io_in_3_b_ready,
  output        io_in_3_b_valid,
  output        io_in_3_ar_ready,
  input         io_in_3_ar_valid,
  input  [31:0] io_in_3_ar_bits_addr,
  input  [2:0]  io_in_3_ar_bits_size,
  input         io_in_3_r_ready,
  output        io_in_3_r_valid,
  output [63:0] io_in_3_r_bits_data,
  output        io_in_3_r_bits_last,
  output        io_in_4_aw_ready,
  input         io_in_4_aw_valid,
  input  [31:0] io_in_4_aw_bits_addr,
  input  [3:0]  io_in_4_aw_bits_id,
  input  [7:0]  io_in_4_aw_bits_len,
  input  [2:0]  io_in_4_aw_bits_size,
  input  [1:0]  io_in_4_aw_bits_burst,
  output        io_in_4_w_ready,
  input         io_in_4_w_valid,
  input  [7:0]  io_in_4_w_bits_strb,
  input  [63:0] io_in_4_w_bits_data,
  input         io_in_4_b_ready,
  output        io_in_4_b_valid,
  output        io_in_4_ar_ready,
  input         io_in_4_ar_valid,
  input  [31:0] io_in_4_ar_bits_addr,
  input  [2:0]  io_in_4_ar_bits_size,
  input         io_in_4_r_ready,
  output        io_in_4_r_valid,
  output [63:0] io_in_4_r_bits_data,
  output        io_in_4_r_bits_last,
  output        io_in_5_aw_ready,
  input         io_in_5_aw_valid,
  input  [31:0] io_in_5_aw_bits_addr,
  input  [3:0]  io_in_5_aw_bits_id,
  input  [7:0]  io_in_5_aw_bits_len,
  input  [2:0]  io_in_5_aw_bits_size,
  input  [1:0]  io_in_5_aw_bits_burst,
  output        io_in_5_w_ready,
  input         io_in_5_w_valid,
  input  [7:0]  io_in_5_w_bits_strb,
  input  [63:0] io_in_5_w_bits_data,
  input         io_in_5_b_ready,
  output        io_in_5_b_valid,
  output        io_in_5_ar_ready,
  input         io_in_5_ar_valid,
  input  [31:0] io_in_5_ar_bits_addr,
  input  [2:0]  io_in_5_ar_bits_size,
  input         io_in_5_r_ready,
  output        io_in_5_r_valid,
  output [63:0] io_in_5_r_bits_data,
  output        io_in_5_r_bits_last,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  output [3:0]  io_out_aw_bits_id,
  output [7:0]  io_out_aw_bits_len,
  output [2:0]  io_out_aw_bits_size,
  output [1:0]  io_out_aw_bits_burst,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [7:0]  io_out_w_bits_strb,
  output [63:0] io_out_w_bits_data,
  output        io_out_w_bits_last,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output [1:0]  io_out_ar_bits_burst,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data,
  input         io_out_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif
  wire  r_arb_io_in_0_ready;
  wire  r_arb_io_in_0_valid;
  wire  r_arb_io_in_1_ready;
  wire  r_arb_io_in_1_valid;
  wire  r_arb_io_in_2_ready;
  wire  r_arb_io_in_2_valid;
  wire  r_arb_io_in_3_ready;
  wire  r_arb_io_in_3_valid;
  wire  r_arb_io_in_4_ready;
  wire  r_arb_io_in_4_valid;
  wire  r_arb_io_in_5_ready;
  wire  r_arb_io_out_ready;
  wire [2:0] r_arb_io_chosen;
  wire  w_arb_io_in_0_ready;
  wire  w_arb_io_in_0_valid;
  wire  w_arb_io_in_1_ready;
  wire  w_arb_io_in_1_valid;
  wire  w_arb_io_in_2_ready;
  wire  w_arb_io_in_2_valid;
  wire  w_arb_io_in_3_ready;
  wire  w_arb_io_in_3_valid;
  wire  w_arb_io_in_4_ready;
  wire  w_arb_io_in_4_valid;
  wire  w_arb_io_in_5_ready;
  wire  w_arb_io_out_ready;
  wire [2:0] w_arb_io_chosen;
  reg [2:0] r_port;
  reg [2:0] w_port;
  reg  r_state;
  wire  _r_chosen_mux_T = ~r_state;
  wire [5:0] r_chosen = {{3'd0}, r_arb_io_chosen};
  wire [5:0] r_chosen_mux = ~r_state ? r_chosen : {{3'd0}, r_port};
  wire  _GEN_1 = 3'h1 == r_chosen_mux[2:0] ? io_in_1_ar_valid : io_in_0_ar_valid;
  wire  _GEN_2 = 3'h2 == r_chosen_mux[2:0] ? io_in_2_ar_valid : _GEN_1;
  wire  _GEN_3 = 3'h3 == r_chosen_mux[2:0] ? io_in_3_ar_valid : _GEN_2;
  wire  _GEN_4 = 3'h4 == r_chosen_mux[2:0] ? io_in_4_ar_valid : _GEN_3;
  wire  _GEN_5 = 3'h5 == r_chosen_mux[2:0] ? io_in_5_ar_valid : _GEN_4;
  wire [31:0] _GEN_7 = 3'h1 == r_chosen_mux[2:0] ? io_in_1_ar_bits_addr : io_in_0_ar_bits_addr;
  wire [31:0] _GEN_8 = 3'h2 == r_chosen_mux[2:0] ? io_in_2_ar_bits_addr : _GEN_7;
  wire [31:0] _GEN_9 = 3'h3 == r_chosen_mux[2:0] ? io_in_3_ar_bits_addr : _GEN_8;
  wire [31:0] _GEN_10 = 3'h4 == r_chosen_mux[2:0] ? io_in_4_ar_bits_addr : _GEN_9;
  wire [7:0] _GEN_20 = 3'h2 == r_chosen_mux[2:0] ? 8'h0 : 8'h1;
  wire [7:0] _GEN_21 = 3'h3 == r_chosen_mux[2:0] ? 8'h0 : _GEN_20;
  wire [7:0] _GEN_22 = 3'h4 == r_chosen_mux[2:0] ? 8'h0 : _GEN_21;
  wire [2:0] _GEN_25 = 3'h1 == r_chosen_mux[2:0] ? io_in_1_ar_bits_size : io_in_0_ar_bits_size;
  wire [2:0] _GEN_26 = 3'h2 == r_chosen_mux[2:0] ? io_in_2_ar_bits_size : _GEN_25;
  wire [2:0] _GEN_27 = 3'h3 == r_chosen_mux[2:0] ? io_in_3_ar_bits_size : _GEN_26;
  wire [2:0] _GEN_28 = 3'h4 == r_chosen_mux[2:0] ? io_in_4_ar_bits_size : _GEN_27;
  wire [1:0] _GEN_32 = 3'h2 == r_chosen_mux[2:0] ? 2'h1 : 2'h2;
  wire [1:0] _GEN_33 = 3'h3 == r_chosen_mux[2:0] ? 2'h1 : _GEN_32;
  wire [1:0] _GEN_34 = 3'h4 == r_chosen_mux[2:0] ? 2'h1 : _GEN_33;
  wire  _GEN_49 = 3'h1 == r_port ? io_in_1_r_ready : io_in_0_r_ready;
  wire  _GEN_50 = 3'h2 == r_port ? io_in_2_r_ready : _GEN_49;
  wire  _GEN_51 = 3'h3 == r_port ? io_in_3_r_ready : _GEN_50;
  wire  _GEN_52 = 3'h4 == r_port ? io_in_4_r_ready : _GEN_51;
  wire  _GEN_53 = 3'h5 == r_port ? io_in_5_r_ready : _GEN_52;
  wire  _GEN_55 = 3'h1 == r_chosen[2:0] ? io_in_1_ar_ready : io_in_0_ar_ready;
  wire  _GEN_56 = 3'h2 == r_chosen[2:0] ? io_in_2_ar_ready : _GEN_55;
  wire  _GEN_57 = 3'h3 == r_chosen[2:0] ? io_in_3_ar_ready : _GEN_56;
  wire  _GEN_58 = 3'h4 == r_chosen[2:0] ? io_in_4_ar_ready : _GEN_57;
  wire  _GEN_59 = 3'h5 == r_chosen[2:0] ? io_in_5_ar_ready : _GEN_58;
  wire  _GEN_61 = 3'h1 == r_chosen[2:0] ? io_in_1_ar_valid : io_in_0_ar_valid;
  wire  _GEN_62 = 3'h2 == r_chosen[2:0] ? io_in_2_ar_valid : _GEN_61;
  wire  _GEN_63 = 3'h3 == r_chosen[2:0] ? io_in_3_ar_valid : _GEN_62;
  wire  _GEN_64 = 3'h4 == r_chosen[2:0] ? io_in_4_ar_valid : _GEN_63;
  wire  _GEN_65 = 3'h5 == r_chosen[2:0] ? io_in_5_ar_valid : _GEN_64;
  wire  _T_2 = _GEN_59 & _GEN_65;
  wire [5:0] _GEN_66 = _T_2 ? r_chosen : {{3'd0}, r_port};
  wire  _GEN_67 = _T_2 | r_state;
  wire  _GEN_69 = 3'h1 == r_port ? io_in_1_r_valid : io_in_0_r_valid;
  wire  _GEN_70 = 3'h2 == r_port ? io_in_2_r_valid : _GEN_69;
  wire  _GEN_71 = 3'h3 == r_port ? io_in_3_r_valid : _GEN_70;
  wire  _GEN_72 = 3'h4 == r_port ? io_in_4_r_valid : _GEN_71;
  wire  _GEN_73 = 3'h5 == r_port ? io_in_5_r_valid : _GEN_72;
  wire  _T_4 = _GEN_53 & _GEN_73;
  wire  _GEN_75 = 3'h1 == r_port ? io_in_1_r_bits_last : io_in_0_r_bits_last;
  wire  _GEN_76 = 3'h2 == r_port ? io_in_2_r_bits_last : _GEN_75;
  wire  _GEN_77 = 3'h3 == r_port ? io_in_3_r_bits_last : _GEN_76;
  wire  _GEN_78 = 3'h4 == r_port ? io_in_4_r_bits_last : _GEN_77;
  wire  _GEN_79 = 3'h5 == r_port ? io_in_5_r_bits_last : _GEN_78;
  wire [5:0] _GEN_82 = _r_chosen_mux_T ? _GEN_66 : {{3'd0}, r_port};
  reg [1:0] w_state;
  wire  _w_chosen_mux_T = w_state == 2'h0;
  wire [5:0] w_chosen = {{3'd0}, w_arb_io_chosen};
  wire [5:0] w_chosen_mux = w_state == 2'h0 ? w_chosen : {{3'd0}, w_port};
  wire  _GEN_85 = 3'h1 == w_chosen_mux[2:0] ? io_in_1_aw_valid : io_in_0_aw_valid;
  wire  _GEN_86 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_valid : _GEN_85;
  wire  _GEN_87 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_valid : _GEN_86;
  wire  _GEN_88 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_valid : _GEN_87;
  wire  _GEN_89 = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_valid : _GEN_88;
  wire [31:0] _GEN_91 = 3'h1 == w_chosen_mux[2:0] ? io_in_1_aw_bits_addr : io_in_0_aw_bits_addr;
  wire [31:0] _GEN_92 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_bits_addr : _GEN_91;
  wire [31:0] _GEN_93 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_bits_addr : _GEN_92;
  wire [31:0] _GEN_94 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_bits_addr : _GEN_93;
  wire [3:0] _GEN_98 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_bits_id : 4'h0;
  wire [3:0] _GEN_99 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_bits_id : _GEN_98;
  wire [3:0] _GEN_100 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_bits_id : _GEN_99;
  wire [7:0] _GEN_104 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_bits_len : 8'h1;
  wire [7:0] _GEN_105 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_bits_len : _GEN_104;
  wire [7:0] _GEN_106 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_bits_len : _GEN_105;
  wire [2:0] _GEN_109 = 3'h1 == w_chosen_mux[2:0] ? io_in_1_aw_bits_size : io_in_0_aw_bits_size;
  wire [2:0] _GEN_110 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_bits_size : _GEN_109;
  wire [2:0] _GEN_111 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_bits_size : _GEN_110;
  wire [2:0] _GEN_112 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_bits_size : _GEN_111;
  wire [1:0] _GEN_116 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_bits_burst : 2'h2;
  wire [1:0] _GEN_117 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_bits_burst : _GEN_116;
  wire [1:0] _GEN_118 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_bits_burst : _GEN_117;
  wire  _GEN_127 = 3'h1 == w_chosen_mux[2:0] ? io_in_1_aw_ready : io_in_0_aw_ready;
  wire  _GEN_128 = 3'h2 == w_chosen_mux[2:0] ? io_in_2_aw_ready : _GEN_127;
  wire  _GEN_129 = 3'h3 == w_chosen_mux[2:0] ? io_in_3_aw_ready : _GEN_128;
  wire  _GEN_130 = 3'h4 == w_chosen_mux[2:0] ? io_in_4_aw_ready : _GEN_129;
  wire  _GEN_131 = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_ready : _GEN_130;
  wire  _w_port_T = _GEN_131 & _GEN_89;
  reg [5:0] w_port_r;
  wire [5:0] _GEN_132 = _w_port_T ? w_chosen : w_port_r;
  wire  _GEN_134 = 3'h1 == w_port ? io_in_1_w_valid : io_in_0_w_valid;
  wire  _GEN_135 = 3'h2 == w_port ? io_in_2_w_valid : _GEN_134;
  wire  _GEN_136 = 3'h3 == w_port ? io_in_3_w_valid : _GEN_135;
  wire  _GEN_137 = 3'h4 == w_port ? io_in_4_w_valid : _GEN_136;
  wire [7:0] _GEN_141 = 3'h2 == w_port ? io_in_2_w_bits_strb : 8'hff;
  wire [7:0] _GEN_142 = 3'h3 == w_port ? io_in_3_w_bits_strb : _GEN_141;
  wire [7:0] _GEN_143 = 3'h4 == w_port ? io_in_4_w_bits_strb : _GEN_142;
  wire [63:0] _GEN_146 = 3'h1 == w_port ? io_in_1_w_bits_data : io_in_0_w_bits_data;
  wire [63:0] _GEN_147 = 3'h2 == w_port ? io_in_2_w_bits_data : _GEN_146;
  wire [63:0] _GEN_148 = 3'h3 == w_port ? io_in_3_w_bits_data : _GEN_147;
  wire [63:0] _GEN_149 = 3'h4 == w_port ? io_in_4_w_bits_data : _GEN_148;
  wire  _GEN_152 = 3'h1 == w_port ? io_in_1_w_bits_last : io_in_0_w_bits_last;
  wire  _GEN_206 = 3'h2 == w_port;
  wire  _GEN_207 = 3'h3 == w_port;
  wire  _GEN_208 = 3'h4 == w_port;
  wire  _GEN_209 = 3'h5 == w_port;
  wire  _GEN_210 = 3'h0 == w_port;
  wire  _GEN_211 = 3'h1 == w_port;
  wire  _GEN_170 = 3'h1 == w_port ? io_in_1_b_ready : io_in_0_b_ready;
  wire  _GEN_171 = 3'h2 == w_port ? io_in_2_b_ready : _GEN_170;
  wire  _GEN_172 = 3'h3 == w_port ? io_in_3_b_ready : _GEN_171;
  wire  _GEN_173 = 3'h4 == w_port ? io_in_4_b_ready : _GEN_172;
  wire  _GEN_174 = 3'h5 == w_port ? io_in_5_b_ready : _GEN_173;
  wire  _GEN_176 = 3'h1 == w_chosen[2:0] ? io_in_1_aw_ready : io_in_0_aw_ready;
  wire  _GEN_177 = 3'h2 == w_chosen[2:0] ? io_in_2_aw_ready : _GEN_176;
  wire  _GEN_178 = 3'h3 == w_chosen[2:0] ? io_in_3_aw_ready : _GEN_177;
  wire  _GEN_179 = 3'h4 == w_chosen[2:0] ? io_in_4_aw_ready : _GEN_178;
  wire  _GEN_180 = 3'h5 == w_chosen[2:0] ? io_in_5_aw_ready : _GEN_179;
  wire  _GEN_182 = 3'h1 == w_chosen[2:0] ? io_in_1_aw_valid : io_in_0_aw_valid;
  wire  _GEN_183 = 3'h2 == w_chosen[2:0] ? io_in_2_aw_valid : _GEN_182;
  wire  _GEN_184 = 3'h3 == w_chosen[2:0] ? io_in_3_aw_valid : _GEN_183;
  wire  _GEN_185 = 3'h4 == w_chosen[2:0] ? io_in_4_aw_valid : _GEN_184;
  wire  _GEN_186 = 3'h5 == w_chosen[2:0] ? io_in_5_aw_valid : _GEN_185;
  wire  _T_8 = _GEN_180 & _GEN_186;
  wire  _T_9 = io_out_w_ready & io_out_w_valid;
  wire  _T_10 = _T_9 & io_out_w_bits_last;
  wire  _GEN_191 = 3'h1 == w_port ? io_in_1_b_valid : io_in_0_b_valid;
  wire  _GEN_192 = 3'h2 == w_port ? io_in_2_b_valid : _GEN_191;
  wire  _GEN_193 = 3'h3 == w_port ? io_in_3_b_valid : _GEN_192;
  wire  _GEN_194 = 3'h4 == w_port ? io_in_4_b_valid : _GEN_193;
  wire  _GEN_195 = 3'h5 == w_port ? io_in_5_b_valid : _GEN_194;
  wire  _T_15 = _GEN_174 & _GEN_195;
  wire [1:0] _GEN_196 = _T_15 ? 2'h0 : w_state;
  wire [5:0] _GEN_241 = reset ? 6'h0 : _GEN_82;
  wire [5:0] _GEN_242 = reset ? 6'h0 : _GEN_132;
  ysyx_040656_Arbiter_1 r_arb (
    .io_in_0_ready(r_arb_io_in_0_ready),
    .io_in_0_valid(r_arb_io_in_0_valid),
    .io_in_1_ready(r_arb_io_in_1_ready),
    .io_in_1_valid(r_arb_io_in_1_valid),
    .io_in_2_ready(r_arb_io_in_2_ready),
    .io_in_2_valid(r_arb_io_in_2_valid),
    .io_in_3_ready(r_arb_io_in_3_ready),
    .io_in_3_valid(r_arb_io_in_3_valid),
    .io_in_4_ready(r_arb_io_in_4_ready),
    .io_in_4_valid(r_arb_io_in_4_valid),
    .io_in_5_ready(r_arb_io_in_5_ready),
    .io_out_ready(r_arb_io_out_ready),
    .io_chosen(r_arb_io_chosen)
  );
  ysyx_040656_Arbiter_1 w_arb (
    .io_in_0_ready(w_arb_io_in_0_ready),
    .io_in_0_valid(w_arb_io_in_0_valid),
    .io_in_1_ready(w_arb_io_in_1_ready),
    .io_in_1_valid(w_arb_io_in_1_valid),
    .io_in_2_ready(w_arb_io_in_2_ready),
    .io_in_2_valid(w_arb_io_in_2_valid),
    .io_in_3_ready(w_arb_io_in_3_ready),
    .io_in_3_valid(w_arb_io_in_3_valid),
    .io_in_4_ready(w_arb_io_in_4_ready),
    .io_in_4_valid(w_arb_io_in_4_valid),
    .io_in_5_ready(w_arb_io_in_5_ready),
    .io_out_ready(w_arb_io_out_ready),
    .io_chosen(w_arb_io_chosen)
  );
  assign io_in_0_aw_ready = 3'h0 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_0_ready;
  assign io_in_0_w_ready = 3'h0 == w_port & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_0_b_valid = _GEN_210 & io_out_b_valid;
  assign io_in_0_ar_ready = 3'h0 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_0_ready;
  assign io_in_0_r_valid = 3'h0 == r_port & io_out_r_valid;
  assign io_in_0_r_bits_data = io_out_r_bits_data;
  assign io_in_0_r_bits_last = io_out_r_bits_last;
  assign io_in_1_aw_ready = 3'h1 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_1_ready;
  assign io_in_1_w_ready = 3'h1 == w_port & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_1_b_valid = _GEN_211 & io_out_b_valid;
  assign io_in_1_ar_ready = 3'h1 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_1_ready;
  assign io_in_1_r_valid = 3'h1 == r_port & io_out_r_valid;
  assign io_in_1_r_bits_data = io_out_r_bits_data;
  assign io_in_1_r_bits_last = io_out_r_bits_last;
  assign io_in_2_aw_ready = 3'h2 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_2_ready;
  assign io_in_2_w_ready = _GEN_206 & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_2_b_valid = _GEN_206 & io_out_b_valid;
  assign io_in_2_ar_ready = 3'h2 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_2_ready;
  assign io_in_2_r_valid = 3'h2 == r_port & io_out_r_valid;
  assign io_in_2_r_bits_data = io_out_r_bits_data;
  assign io_in_2_r_bits_last = io_out_r_bits_last;
  assign io_in_3_aw_ready = 3'h3 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_3_ready;
  assign io_in_3_w_ready = _GEN_207 & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_3_b_valid = _GEN_207 & io_out_b_valid;
  assign io_in_3_ar_ready = 3'h3 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_3_ready;
  assign io_in_3_r_valid = 3'h3 == r_port & io_out_r_valid;
  assign io_in_3_r_bits_data = io_out_r_bits_data;
  assign io_in_3_r_bits_last = io_out_r_bits_last;
  assign io_in_4_aw_ready = 3'h4 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_4_ready;
  assign io_in_4_w_ready = _GEN_208 & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_4_b_valid = _GEN_208 & io_out_b_valid;
  assign io_in_4_ar_ready = 3'h4 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_4_ready;
  assign io_in_4_r_valid = 3'h4 == r_port & io_out_r_valid;
  assign io_in_4_r_bits_data = io_out_r_bits_data;
  assign io_in_4_r_bits_last = io_out_r_bits_last;
  assign io_in_5_aw_ready = 3'h5 == w_chosen_mux[2:0] ? io_out_aw_ready & _w_chosen_mux_T : w_arb_io_in_5_ready;
  assign io_in_5_w_ready = _GEN_209 & (io_out_w_ready & (w_state == 2'h1 | _w_chosen_mux_T));
  assign io_in_5_b_valid = _GEN_209 & io_out_b_valid;
  assign io_in_5_ar_ready = 3'h5 == r_chosen_mux[2:0] ? io_out_ar_ready & _r_chosen_mux_T : r_arb_io_in_5_ready;
  assign io_in_5_r_valid = 3'h5 == r_port & io_out_r_valid;
  assign io_in_5_r_bits_data = io_out_r_bits_data;
  assign io_in_5_r_bits_last = io_out_r_bits_last;
  assign io_out_aw_valid = _GEN_89 & _w_chosen_mux_T;
  assign io_out_aw_bits_addr = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_bits_addr : _GEN_94;
  assign io_out_aw_bits_id = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_bits_id : _GEN_100;
  assign io_out_aw_bits_len = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_bits_len : _GEN_106;
  assign io_out_aw_bits_size = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_bits_size : _GEN_112;
  assign io_out_aw_bits_burst = 3'h5 == w_chosen_mux[2:0] ? io_in_5_aw_bits_burst : _GEN_118;
  assign io_out_w_valid = 3'h5 == w_port ? io_in_5_w_valid : _GEN_137;
  assign io_out_w_bits_strb = 3'h5 == w_port ? io_in_5_w_bits_strb : _GEN_143;
  assign io_out_w_bits_data = 3'h5 == w_port ? io_in_5_w_bits_data : _GEN_149;
  assign io_out_w_bits_last = 3'h5 == w_port | (3'h4 == w_port | (3'h3 == w_port | (3'h2 == w_port | _GEN_152)));
  assign io_out_b_ready = 3'h5 == w_port ? io_in_5_b_ready : _GEN_173;
  assign io_out_ar_valid = _GEN_5 & _r_chosen_mux_T;
  assign io_out_ar_bits_addr = 3'h5 == r_chosen_mux[2:0] ? io_in_5_ar_bits_addr : _GEN_10;
  assign io_out_ar_bits_len = 3'h5 == r_chosen_mux[2:0] ? 8'h0 : _GEN_22;
  assign io_out_ar_bits_size = 3'h5 == r_chosen_mux[2:0] ? io_in_5_ar_bits_size : _GEN_28;
  assign io_out_ar_bits_burst = 3'h5 == r_chosen_mux[2:0] ? 2'h1 : _GEN_34;
  assign io_out_r_ready = 3'h5 == r_port ? io_in_5_r_ready : _GEN_52;
  assign r_arb_io_in_0_valid = io_in_0_ar_valid;
  assign r_arb_io_in_1_valid = io_in_1_ar_valid;
  assign r_arb_io_in_2_valid = io_in_2_ar_valid;
  assign r_arb_io_in_3_valid = io_in_3_ar_valid;
  assign r_arb_io_in_4_valid = io_in_4_ar_valid;
  assign r_arb_io_out_ready = io_out_ar_ready & _r_chosen_mux_T;
  assign w_arb_io_in_0_valid = io_in_0_aw_valid;
  assign w_arb_io_in_1_valid = io_in_1_aw_valid;
  assign w_arb_io_in_2_valid = io_in_2_aw_valid;
  assign w_arb_io_in_3_valid = io_in_3_aw_valid;
  assign w_arb_io_in_4_valid = io_in_4_aw_valid;
  assign w_arb_io_out_ready = io_out_aw_ready & _w_chosen_mux_T;
  always @(posedge clock) begin
    r_port <= _GEN_241[2:0];
    w_port <= _GEN_242[2:0];
    if (reset) begin
      r_state <= 1'h0;
    end else if (_r_chosen_mux_T) begin
      r_state <= _GEN_67;
    end else if (r_state) begin
      if (_T_4 & _GEN_79) begin
        r_state <= 1'h0;
      end
    end
    if (reset) begin
      w_state <= 2'h0;
    end else if (2'h0 == w_state) begin
      if (_T_8) begin
        if (_T_9 & io_out_w_bits_last) begin
          w_state <= 2'h2;
        end else begin
          w_state <= 2'h1;
        end
      end
    end else if (2'h1 == w_state) begin
      if (_T_10) begin
        w_state <= 2'h2;
      end
    end else if (2'h2 == w_state) begin
      w_state <= _GEN_196;
    end
    if (reset) begin
      w_port_r <= 6'h0;
    end else if (_w_port_T) begin
      w_port_r <= w_chosen;
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_port = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  w_port = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  r_state = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  w_port_r = _RAND_4[5:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_CoreLinkXBar(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [1:0]  io_in_req_bits_size,
  input  [2:0]  io_in_req_bits_cmd,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [63:0] io_out_0_req_bits_wdata,
  output [1:0]  io_out_0_req_bits_size,
  output [2:0]  io_out_0_req_bits_cmd,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [63:0] io_out_1_req_bits_wdata,
  output [1:0]  io_out_1_req_bits_size,
  output [2:0]  io_out_1_req_bits_cmd,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [63:0] io_out_2_req_bits_wdata,
  output [1:0]  io_out_2_req_bits_size,
  output [2:0]  io_out_2_req_bits_cmd,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata,
  input         io_out_3_req_ready,
  output        io_out_3_req_valid,
  output [31:0] io_out_3_req_bits_addr,
  output [63:0] io_out_3_req_bits_wdata,
  output [1:0]  io_out_3_req_bits_size,
  output [2:0]  io_out_3_req_bits_cmd,
  output        io_out_3_resp_ready,
  input         io_out_3_resp_valid,
  input  [63:0] io_out_3_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif
  reg [1:0] state;
  wire  outSelVec_0 = io_in_req_bits_addr <= 32'h1ffffff;
  wire  outSelVec_1 = io_in_req_bits_addr >= 32'h2000000 & io_in_req_bits_addr <= 32'h200ffff;
  wire  outSelVec_2 = io_in_req_bits_addr >= 32'h2010000 & io_in_req_bits_addr <= 32'h7fffffff;
  wire  outSelVec_3 = io_in_req_bits_addr >= 32'hfc000000;
  wire [1:0] _outSelIdx_T = outSelVec_2 ? 2'h2 : 2'h3;
  wire [1:0] _outSelIdx_T_1 = outSelVec_1 ? 2'h1 : _outSelIdx_T;
  wire [1:0] outSelIdx = outSelVec_0 ? 2'h0 : _outSelIdx_T_1;
  wire  _GEN_1 = 2'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready;
  wire  _GEN_2 = 2'h2 == outSelIdx ? io_out_2_req_ready : _GEN_1;
  wire  _GEN_3 = 2'h3 == outSelIdx ? io_out_3_req_ready : _GEN_2;
  wire  _GEN_5 = 2'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid;
  wire  _GEN_6 = 2'h2 == outSelIdx ? io_out_2_req_valid : _GEN_5;
  wire  _GEN_7 = 2'h3 == outSelIdx ? io_out_3_req_valid : _GEN_6;
  wire  _outSelIdxResp_T = _GEN_3 & _GEN_7;
  wire  _outSelIdxResp_T_1 = state == 2'h0;
  wire  _outSelIdxResp_T_2 = _outSelIdxResp_T & state == 2'h0;
  reg [1:0] outSelIdxResp;
  wire [3:0] _reqInvalidAddr_hit_T = {outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0};
  wire  reqInvalidAddr_hit = |_reqInvalidAddr_hit_T;
  wire  reqInvalidAddr = io_in_req_valid & reqInvalidAddr_hit & ~reqInvalidAddr_hit;
  wire  _GEN_12 = 2'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready;
  wire  _GEN_13 = 2'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_12;
  wire  _GEN_14 = 2'h3 == outSelIdxResp ? io_out_3_resp_ready : _GEN_13;
  wire  _GEN_16 = 2'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid;
  wire  _GEN_17 = 2'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_16;
  wire  _GEN_18 = 2'h3 == outSelIdxResp ? io_out_3_resp_valid : _GEN_17;
  wire  _T_3 = _GEN_14 & _GEN_18;
  wire [1:0] _GEN_20 = io_in_resp_valid ? 2'h0 : state;
  wire [63:0] _GEN_29 = 2'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata;
  wire [63:0] _GEN_30 = 2'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_29;
  assign io_in_req_ready = _GEN_3 | reqInvalidAddr;
  assign io_in_resp_valid = _T_3 | state == 2'h2;
  assign io_in_resp_bits_rdata = 2'h3 == outSelIdxResp ? io_out_3_resp_bits_rdata : _GEN_30;
  assign io_out_0_req_valid = outSelVec_0 & (io_in_req_valid & _outSelIdxResp_T_1);
  assign io_out_0_req_bits_addr = io_in_req_bits_addr;
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata;
  assign io_out_0_req_bits_size = io_in_req_bits_size;
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd;
  assign io_out_0_resp_ready = 2'h0 == outSelIdxResp | outSelVec_0;
  assign io_out_1_req_valid = outSelVec_1 & (io_in_req_valid & _outSelIdxResp_T_1);
  assign io_out_1_req_bits_addr = io_in_req_bits_addr;
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata;
  assign io_out_1_req_bits_size = io_in_req_bits_size;
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd;
  assign io_out_1_resp_ready = 2'h1 == outSelIdxResp | outSelVec_1;
  assign io_out_2_req_valid = outSelVec_2 & (io_in_req_valid & _outSelIdxResp_T_1);
  assign io_out_2_req_bits_addr = io_in_req_bits_addr;
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata;
  assign io_out_2_req_bits_size = io_in_req_bits_size;
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd;
  assign io_out_2_resp_ready = 2'h2 == outSelIdxResp | outSelVec_2;
  assign io_out_3_req_valid = outSelVec_3 & (io_in_req_valid & _outSelIdxResp_T_1);
  assign io_out_3_req_bits_addr = io_in_req_bits_addr;
  assign io_out_3_req_bits_wdata = io_in_req_bits_wdata;
  assign io_out_3_req_bits_size = io_in_req_bits_size;
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd;
  assign io_out_3_resp_ready = 2'h3 == outSelIdxResp | outSelVec_3;
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (2'h0 == state) begin
      if (reqInvalidAddr) begin
        state <= 2'h2;
      end else if (_outSelIdxResp_T) begin
        state <= 2'h1;
      end
    end else if (2'h1 == state) begin
      if (_T_3) begin
        state <= 2'h0;
      end
    end else if (2'h2 == state) begin
      state <= _GEN_20;
    end
    if (_outSelIdxResp_T_2) begin
      if (outSelVec_0) begin
        outSelIdxResp <= 2'h0;
      end else if (outSelVec_1) begin
        outSelIdxResp <= 2'h1;
      end else if (outSelVec_2) begin
        outSelIdxResp <= 2'h2;
      end else begin
        outSelIdxResp <= 2'h3;
      end
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[1:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_AXI4Bridge(
  input          clock,
  input          reset,
  output         io_in_req_ready,
  input          io_in_req_valid,
  input  [31:0]  io_in_req_bits_addr,
  input  [127:0] io_in_req_bits_wdata,
  input  [2:0]   io_in_req_bits_cmd,
  output         io_in_resp_valid,
  output [2:0]   io_in_resp_bits_cmd,
  output [127:0] io_in_resp_bits_rdata,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  output [2:0]   io_out_aw_bits_size,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output         io_out_w_bits_last,
  output         io_out_b_ready,
  input          io_out_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output [2:0]   io_out_ar_bits_size,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif
  reg [2:0] reg_state;
  reg [127:0] dataReadBuffer;
  reg [127:0] dataWriterBuffer;
  reg  readBeatCnt_value;
  reg  writeBeatCnt_value;
  reg [31:0] startAddr;
  reg [1:0] size;
  reg  axi_wen;
  wire  _io_in_resp_valid_T = reg_state == 3'h5;
  wire [31:0] addr = {io_in_req_bits_addr[31:3],3'h0};
  wire [63:0] wblock_0 = dataWriterBuffer[63:0];
  wire [63:0] wblock_1 = dataWriterBuffer[127:64];
  wire  _T_1 = io_in_req_ready & io_in_req_valid;
  wire  _T_3 = io_out_ar_ready & io_out_ar_valid;
  wire [31:0] _value_T = startAddr >> size;
  wire [31:0] _value_T_1 = _value_T & 32'h1;
  wire  _T_4 = io_out_aw_ready & io_out_aw_valid;
  wire [2:0] _GEN_5 = _T_4 ? 3'h2 : reg_state;
  wire [31:0] _GEN_7 = _T_3 ? _value_T_1 : {{31'd0}, readBeatCnt_value};
  wire  _T_6 = io_out_w_ready & io_out_w_valid;
  wire  _GEN_8 = writeBeatCnt_value ? 1'h0 : writeBeatCnt_value + 1'h1;
  wire [2:0] _GEN_9 = writeBeatCnt_value ? 3'h4 : reg_state;
  wire  _GEN_10 = _T_6 ? _GEN_8 : writeBeatCnt_value;
  wire [2:0] _GEN_11 = _T_6 ? _GEN_9 : reg_state;
  wire  _T_8 = io_out_r_ready & io_out_r_valid;
  wire [63:0] nextBlock_0 = ~readBeatCnt_value ? io_out_r_bits_data : dataReadBuffer[63:0];
  wire [63:0] nextBlock_1 = readBeatCnt_value ? io_out_r_bits_data : dataReadBuffer[127:64];
  wire [127:0] _dataReadBuffer_T = {nextBlock_1,nextBlock_0};
  wire  _GEN_14 = io_out_r_bits_last ? 1'h0 : readBeatCnt_value + 1'h1;
  wire [2:0] _GEN_15 = io_out_r_bits_last ? 3'h5 : reg_state;
  wire  _GEN_16 = readBeatCnt_value ? 1'h0 : _GEN_14;
  wire [127:0] _GEN_17 = _T_8 ? _dataReadBuffer_T : dataReadBuffer;
  wire  _GEN_18 = _T_8 ? _GEN_16 : readBeatCnt_value;
  wire [2:0] _GEN_19 = _T_8 ? _GEN_15 : reg_state;
  wire  _T_11 = io_out_b_ready & io_out_b_valid;
  wire [2:0] _GEN_20 = _T_11 ? 3'h5 : reg_state;
  wire [2:0] _GEN_21 = io_in_resp_valid ? 3'h0 : reg_state;
  wire [2:0] _GEN_22 = 3'h5 == reg_state ? _GEN_21 : reg_state;
  wire [2:0] _GEN_23 = 3'h4 == reg_state ? _GEN_20 : _GEN_22;
  wire [127:0] _GEN_24 = 3'h3 == reg_state ? _GEN_17 : dataReadBuffer;
  wire  _GEN_25 = 3'h3 == reg_state ? _GEN_18 : readBeatCnt_value;
  wire [2:0] _GEN_26 = 3'h3 == reg_state ? _GEN_19 : _GEN_23;
  wire  _GEN_30 = 3'h2 == reg_state ? readBeatCnt_value : _GEN_25;
  wire [31:0] _GEN_32 = 3'h1 == reg_state ? _GEN_7 : {{31'd0}, _GEN_30};
  wire [31:0] _GEN_40 = 3'h0 == reg_state ? {{31'd0}, readBeatCnt_value} : _GEN_32;
  wire  _io_out_ar_valid_T = reg_state == 3'h1;
  wire [31:0] _GEN_45 = reset ? 32'h0 : _GEN_40;
  assign io_in_req_ready = reg_state == 3'h0;
  assign io_in_resp_valid = reg_state == 3'h5;
  assign io_in_resp_bits_cmd = axi_wen ? 3'h4 : 3'h3;
  assign io_in_resp_bits_rdata = _io_in_resp_valid_T ? dataReadBuffer : 128'h0;
  assign io_out_aw_valid = _io_out_ar_valid_T & axi_wen;
  assign io_out_aw_bits_addr = startAddr;
  assign io_out_aw_bits_size = {{1'd0}, size};
  assign io_out_w_valid = reg_state == 3'h2 & axi_wen;
  assign io_out_w_bits_data = writeBeatCnt_value ? wblock_1 : wblock_0;
  assign io_out_w_bits_last = writeBeatCnt_value;
  assign io_out_b_ready = reg_state == 3'h4;
  assign io_out_ar_valid = reg_state == 3'h1 & ~axi_wen;
  assign io_out_ar_bits_addr = startAddr;
  assign io_out_ar_bits_size = {{1'd0}, size};
  assign io_out_r_ready = reg_state == 3'h3;
  always @(posedge clock) begin
    if (reset) begin
      reg_state <= 3'h0;
    end else if (3'h0 == reg_state) begin
      if (_T_1) begin
        reg_state <= 3'h1;
      end
    end else if (3'h1 == reg_state) begin
      if (_T_3) begin
        reg_state <= 3'h3;
      end else begin
        reg_state <= _GEN_5;
      end
    end else if (3'h2 == reg_state) begin
      reg_state <= _GEN_11;
    end else begin
      reg_state <= _GEN_26;
    end
    if (reset) begin
      dataReadBuffer <= 128'h0;
    end else if (!(3'h0 == reg_state)) begin
      if (!(3'h1 == reg_state)) begin
        if (!(3'h2 == reg_state)) begin
          dataReadBuffer <= _GEN_24;
        end
      end
    end
    if (reset) begin
      dataWriterBuffer <= 128'h0;
    end else if (3'h0 == reg_state) begin
      if (_T_1) begin
        dataWriterBuffer <= io_in_req_bits_wdata;
      end
    end
    readBeatCnt_value <= _GEN_45[0];
    if (reset) begin
      writeBeatCnt_value <= 1'h0;
    end else if (!(3'h0 == reg_state)) begin
      if (!(3'h1 == reg_state)) begin
        if (3'h2 == reg_state) begin
          writeBeatCnt_value <= _GEN_10;
        end
      end
    end
    if (reset) begin
      startAddr <= 32'h0;
    end else if (3'h0 == reg_state) begin
      if (_T_1) begin
        startAddr <= addr;
      end
    end
    if (reset) begin
      size <= 2'h0;
    end else if (3'h0 == reg_state) begin
      if (_T_1) begin
        size <= 2'h3;
      end
    end
    if (reset) begin
      axi_wen <= 1'h0;
    end else if (3'h0 == reg_state) begin
      if (_T_1) begin
        axi_wen <= io_in_req_bits_cmd == 3'h1;
      end
    end
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_state = _RAND_0[2:0];
  _RAND_1 = {4{`RANDOM}};
  dataReadBuffer = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  dataWriterBuffer = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  readBeatCnt_value = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  writeBeatCnt_value = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  startAddr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  size = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  axi_wen = _RAND_7[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_CoreLink2AXI4(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [1:0]  io_in_req_bits_size,
  input  [2:0]  io_in_req_bits_cmd,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [7:0]  io_out_w_bits_strb,
  output [63:0] io_out_w_bits_data,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif
  wire [3:0] io_out_w_bits_strb_numValid = 4'h1 << io_in_req_bits_size;
  wire [3:0] _GEN_5 = {{1'd0}, io_in_req_bits_addr[2:0]};
  wire [3:0] _io_out_w_bits_strb_wmask_0_T_4 = _GEN_5 + io_out_w_bits_strb_numValid;
  wire  io_out_w_bits_strb_wmask_0 = io_in_req_bits_addr[2:0] <= 3'h0 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h0;
  wire  io_out_w_bits_strb_wmask_1 = io_in_req_bits_addr[2:0] <= 3'h1 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h1;
  wire  io_out_w_bits_strb_wmask_2 = io_in_req_bits_addr[2:0] <= 3'h2 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h2;
  wire  io_out_w_bits_strb_wmask_3 = io_in_req_bits_addr[2:0] <= 3'h3 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h3;
  wire  io_out_w_bits_strb_wmask_4 = io_in_req_bits_addr[2:0] <= 3'h4 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h4;
  wire  io_out_w_bits_strb_wmask_5 = io_in_req_bits_addr[2:0] <= 3'h5 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h5;
  wire  io_out_w_bits_strb_wmask_6 = io_in_req_bits_addr[2:0] <= 3'h6 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h6;
  wire  io_out_w_bits_strb_wmask_7 = _io_out_w_bits_strb_wmask_0_T_4 > 4'h7;
  wire [3:0] io_out_w_bits_strb_lo = {io_out_w_bits_strb_wmask_3,io_out_w_bits_strb_wmask_2,io_out_w_bits_strb_wmask_1,
    io_out_w_bits_strb_wmask_0};
  wire [3:0] io_out_w_bits_strb_hi = {io_out_w_bits_strb_wmask_7,io_out_w_bits_strb_wmask_6,io_out_w_bits_strb_wmask_5,
    io_out_w_bits_strb_wmask_4};
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid;
  reg  awAck;
  wire  _GEN_0 = _awAck_T | awAck;
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid;
  reg  wAck;
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck;
  wire  _GEN_2 = _wSend_T_1 | wAck;
  wire  _wen_T_2 = io_in_req_bits_cmd == 3'h1 | io_in_req_bits_cmd == 3'h4;
  wire  _wen_T_3 = io_in_req_ready & io_in_req_valid;
  reg  wen;
  wire  _io_out_ar_valid_T_2 = io_in_req_bits_cmd == 3'h0 | io_in_req_bits_cmd == 3'h3;
  wire  _io_out_aw_valid_T_3 = io_in_req_valid & _wen_T_2;
  wire  _io_out_w_valid_T_4 = ~wAck;
  assign io_in_req_ready = _wen_T_2 ? _io_out_w_valid_T_4 & io_out_w_ready : io_out_ar_ready;
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid;
  assign io_in_resp_bits_rdata = io_out_r_bits_data;
  assign io_out_aw_valid = _io_out_aw_valid_T_3 & ~awAck;
  assign io_out_aw_bits_addr = io_out_ar_bits_addr;
  assign io_out_w_valid = _io_out_aw_valid_T_3 & ~wAck;
  assign io_out_w_bits_strb = {io_out_w_bits_strb_hi,io_out_w_bits_strb_lo};
  assign io_out_w_bits_data = io_in_req_bits_wdata;
  assign io_out_b_ready = io_in_resp_ready;
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_2;
  assign io_out_ar_bits_addr = io_in_req_bits_addr;
  assign io_out_r_ready = io_in_resp_ready;
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_3) begin
      wen <= _wen_T_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656_CoreLink2AXI4_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [1:0]  io_in_req_bits_size,
  input  [2:0]  io_in_req_bits_cmd,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  output [3:0]  io_out_aw_bits_id,
  output [7:0]  io_out_aw_bits_len,
  output [2:0]  io_out_aw_bits_size,
  output [1:0]  io_out_aw_bits_burst,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [7:0]  io_out_w_bits_strb,
  output [63:0] io_out_w_bits_data,
  output        io_out_w_bits_last,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [3:0]  io_out_ar_bits_id,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output [1:0]  io_out_ar_bits_burst,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif
  wire [3:0] io_out_w_bits_strb_numValid = 4'h1 << io_in_req_bits_size;
  wire [3:0] _GEN_5 = {{1'd0}, io_in_req_bits_addr[2:0]};
  wire [3:0] _io_out_w_bits_strb_wmask_0_T_4 = _GEN_5 + io_out_w_bits_strb_numValid;
  wire  io_out_w_bits_strb_wmask_0 = io_in_req_bits_addr[2:0] <= 3'h0 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h0;
  wire  io_out_w_bits_strb_wmask_1 = io_in_req_bits_addr[2:0] <= 3'h1 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h1;
  wire  io_out_w_bits_strb_wmask_2 = io_in_req_bits_addr[2:0] <= 3'h2 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h2;
  wire  io_out_w_bits_strb_wmask_3 = io_in_req_bits_addr[2:0] <= 3'h3 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h3;
  wire  io_out_w_bits_strb_wmask_4 = io_in_req_bits_addr[2:0] <= 3'h4 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h4;
  wire  io_out_w_bits_strb_wmask_5 = io_in_req_bits_addr[2:0] <= 3'h5 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h5;
  wire  io_out_w_bits_strb_wmask_6 = io_in_req_bits_addr[2:0] <= 3'h6 & _io_out_w_bits_strb_wmask_0_T_4 > 4'h6;
  wire  io_out_w_bits_strb_wmask_7 = _io_out_w_bits_strb_wmask_0_T_4 > 4'h7;
  wire [3:0] io_out_w_bits_strb_lo = {io_out_w_bits_strb_wmask_3,io_out_w_bits_strb_wmask_2,io_out_w_bits_strb_wmask_1,
    io_out_w_bits_strb_wmask_0};
  wire [3:0] io_out_w_bits_strb_hi = {io_out_w_bits_strb_wmask_7,io_out_w_bits_strb_wmask_6,io_out_w_bits_strb_wmask_5,
    io_out_w_bits_strb_wmask_4};
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid;
  reg  awAck;
  wire  _GEN_0 = _awAck_T | awAck;
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid;
  reg  wAck;
  wire  wSend = _awAck_T & _wSend_T_1 & io_out_w_bits_last | awAck & wAck;
  wire  _wAck_T_1 = _wSend_T_1 & io_out_w_bits_last;
  wire  _GEN_2 = _wAck_T_1 | wAck;
  wire  _wen_T_2 = io_in_req_bits_cmd == 3'h1 | io_in_req_bits_cmd == 3'h4;
  wire  _wen_T_3 = io_in_req_ready & io_in_req_valid;
  reg  wen;
  wire  _io_out_ar_valid_T_2 = io_in_req_bits_cmd == 3'h0 | io_in_req_bits_cmd == 3'h3;
  wire  _io_out_aw_valid_T_3 = io_in_req_valid & _wen_T_2;
  wire  _io_out_w_valid_T_4 = ~wAck;
  assign io_in_req_ready = _wen_T_2 ? _io_out_w_valid_T_4 & io_out_w_ready : io_out_ar_ready;
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid;
  assign io_in_resp_bits_rdata = io_out_r_bits_data;
  assign io_out_aw_valid = _io_out_aw_valid_T_3 & ~awAck;
  assign io_out_aw_bits_addr = io_out_ar_bits_addr;
  assign io_out_aw_bits_id = io_out_ar_bits_id;
  assign io_out_aw_bits_len = io_out_ar_bits_len;
  assign io_out_aw_bits_size = io_out_ar_bits_size;
  assign io_out_aw_bits_burst = io_out_ar_bits_burst;
  assign io_out_w_valid = _io_out_aw_valid_T_3 & ~wAck;
  assign io_out_w_bits_strb = {io_out_w_bits_strb_hi,io_out_w_bits_strb_lo};
  assign io_out_w_bits_data = io_in_req_bits_wdata;
  assign io_out_w_bits_last = 1'h1;
  assign io_out_b_ready = io_in_resp_ready;
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_2;
  assign io_out_ar_bits_addr = io_in_req_bits_addr;
  assign io_out_ar_bits_id = 4'h0;
  assign io_out_ar_bits_len = 8'h0;
  assign io_out_ar_bits_size = {{1'd0}, io_in_req_bits_size};
  assign io_out_ar_bits_burst = 2'h1;
  assign io_out_r_ready = io_in_resp_ready;
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_3) begin
      wen <= _wen_T_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~1'h1 & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif
  `endif
end
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif
endmodule
module ysyx_040656(
  input          clock,
  input          reset,
  input          io_interrupt,
  input          io_master_arready,
  output         io_master_arvalid,
  output [31:0]  io_master_araddr,
  output [3:0]   io_master_arid,
  output [7:0]   io_master_arlen,
  output [2:0]   io_master_arsize,
  output [1:0]   io_master_arburst,
  output         io_master_rready,
  input          io_master_rvalid,
  input  [1:0]   io_master_rresp,
  input  [63:0]  io_master_rdata,
  input          io_master_rlast,
  input  [3:0]   io_master_rid,
  input          io_master_awready,
  output         io_master_awvalid,
  output [31:0]  io_master_awaddr,
  output [3:0]   io_master_awid,
  output [7:0]   io_master_awlen,
  output [2:0]   io_master_awsize,
  output [1:0]   io_master_awburst,
  input          io_master_wready,
  output         io_master_wvalid,
  output [63:0]  io_master_wdata,
  output [7:0]   io_master_wstrb,
  output         io_master_wlast,
  output         io_master_bready,
  input          io_master_bvalid,
  input  [1:0]   io_master_bresp,
  input  [3:0]   io_master_bid,
  output         io_slave_arready,
  input          io_slave_arvalid,
  input  [31:0]  io_slave_araddr,
  input  [3:0]   io_slave_arid,
  input  [7:0]   io_slave_arlen,
  input  [2:0]   io_slave_arsize,
  input  [1:0]   io_slave_arburst,
  input          io_slave_rready,
  output         io_slave_rvalid,
  output [1:0]   io_slave_rresp,
  output [63:0]  io_slave_rdata,
  output         io_slave_rlast,
  output [3:0]   io_slave_rid,
  output         io_slave_awready,
  input          io_slave_awvalid,
  input  [31:0]  io_slave_awaddr,
  input  [3:0]   io_slave_awid,
  input  [7:0]   io_slave_awlen,
  input  [2:0]   io_slave_awsize,
  input  [1:0]   io_slave_awburst,
  output         io_slave_wready,
  input          io_slave_wvalid,
  input  [63:0]  io_slave_wdata,
  input  [7:0]   io_slave_wstrb,
  input          io_slave_wlast,
  input          io_slave_bready,
  output         io_slave_bvalid,
  output [1:0]   io_slave_bresp,
  output [3:0]   io_slave_bid,
  input  [127:0] io_sram0_rdata,
  output         io_sram0_wen,
  output         io_sram0_cen,
  output [5:0]   io_sram0_addr,
  output [127:0] io_sram0_wdata,
  output [127:0] io_sram0_wmask,
  input  [127:0] io_sram1_rdata,
  output         io_sram1_wen,
  output         io_sram1_cen,
  output [5:0]   io_sram1_addr,
  output [127:0] io_sram1_wdata,
  output [127:0] io_sram1_wmask,
  input  [127:0] io_sram2_rdata,
  output         io_sram2_wen,
  output         io_sram2_cen,
  output [5:0]   io_sram2_addr,
  output [127:0] io_sram2_wdata,
  output [127:0] io_sram2_wmask,
  input  [127:0] io_sram3_rdata,
  output         io_sram3_wen,
  output         io_sram3_cen,
  output [5:0]   io_sram3_addr,
  output [127:0] io_sram3_wdata,
  output [127:0] io_sram3_wmask,
  input  [127:0] io_sram4_rdata,
  output         io_sram4_wen,
  output         io_sram4_cen,
  output [5:0]   io_sram4_addr,
  output [127:0] io_sram4_wdata,
  output [127:0] io_sram4_wmask,
  input  [127:0] io_sram5_rdata,
  output         io_sram5_wen,
  output         io_sram5_cen,
  output [5:0]   io_sram5_addr,
  output [127:0] io_sram5_wdata,
  output [127:0] io_sram5_wmask,
  input  [127:0] io_sram6_rdata,
  output         io_sram6_wen,
  output         io_sram6_cen,
  output [5:0]   io_sram6_addr,
  output [127:0] io_sram6_wdata,
  output [127:0] io_sram6_wmask,
  input  [127:0] io_sram7_rdata,
  output         io_sram7_wen,
  output         io_sram7_cen,
  output [5:0]   io_sram7_addr,
  output [127:0] io_sram7_wdata,
  output [127:0] io_sram7_wmask
);
  wire  overlay_clock;
  wire  overlay_reset;
  wire  overlay_io_imem_req_ready;
  wire  overlay_io_imem_req_valid;
  wire [31:0] overlay_io_imem_req_bits_addr;
  wire [127:0] overlay_io_imem_req_bits_wdata;
  wire [2:0] overlay_io_imem_req_bits_cmd;
  wire  overlay_io_imem_resp_valid;
  wire [127:0] overlay_io_imem_resp_bits_rdata;
  wire  overlay_io_dmem_req_ready;
  wire  overlay_io_dmem_req_valid;
  wire [31:0] overlay_io_dmem_req_bits_addr;
  wire [127:0] overlay_io_dmem_req_bits_wdata;
  wire [2:0] overlay_io_dmem_req_bits_cmd;
  wire  overlay_io_dmem_resp_valid;
  wire [127:0] overlay_io_dmem_resp_bits_rdata;
  wire  overlay_io_link_req_ready;
  wire  overlay_io_link_req_valid;
  wire [31:0] overlay_io_link_req_bits_addr;
  wire [127:0] overlay_io_link_req_bits_wdata;
  wire  overlay_io_link_resp_valid;
  wire [2:0] overlay_io_link_resp_bits_cmd;
  wire [127:0] overlay_io_link_resp_bits_rdata;
  wire  overlay_io_immio_req_ready;
  wire  overlay_io_immio_req_valid;
  wire [31:0] overlay_io_immio_req_bits_addr;
  wire [1:0] overlay_io_immio_req_bits_size;
  wire  overlay_io_immio_resp_valid;
  wire [63:0] overlay_io_immio_resp_bits_rdata;
  wire  overlay_io_dmmio_req_ready;
  wire  overlay_io_dmmio_req_valid;
  wire [31:0] overlay_io_dmmio_req_bits_addr;
  wire [63:0] overlay_io_dmmio_req_bits_wdata;
  wire [1:0] overlay_io_dmmio_req_bits_size;
  wire [2:0] overlay_io_dmmio_req_bits_cmd;
  wire  overlay_io_dmmio_resp_valid;
  wire [63:0] overlay_io_dmmio_resp_bits_rdata;
  wire [127:0] overlay_io_sram0_rdata;
  wire  overlay_io_sram0_wen;
  wire [5:0] overlay_io_sram0_addr;
  wire [127:0] overlay_io_sram0_wdata;
  wire [127:0] overlay_io_sram1_rdata;
  wire  overlay_io_sram1_wen;
  wire [5:0] overlay_io_sram1_addr;
  wire [127:0] overlay_io_sram1_wdata;
  wire [127:0] overlay_io_sram2_rdata;
  wire  overlay_io_sram2_wen;
  wire [5:0] overlay_io_sram2_addr;
  wire [127:0] overlay_io_sram2_wdata;
  wire [127:0] overlay_io_sram3_rdata;
  wire  overlay_io_sram3_wen;
  wire [5:0] overlay_io_sram3_addr;
  wire [127:0] overlay_io_sram3_wdata;
  wire [127:0] overlay_io_sram4_rdata;
  wire  overlay_io_sram4_wen;
  wire [5:0] overlay_io_sram4_addr;
  wire [127:0] overlay_io_sram4_wdata;
  wire [127:0] overlay_io_sram5_rdata;
  wire  overlay_io_sram5_wen;
  wire [5:0] overlay_io_sram5_addr;
  wire [127:0] overlay_io_sram5_wdata;
  wire [127:0] overlay_io_sram6_rdata;
  wire  overlay_io_sram6_wen;
  wire [5:0] overlay_io_sram6_addr;
  wire [127:0] overlay_io_sram6_wdata;
  wire [127:0] overlay_io_sram7_rdata;
  wire  overlay_io_sram7_wen;
  wire [5:0] overlay_io_sram7_addr;
  wire [127:0] overlay_io_sram7_wdata;
  wire  xConnect_clock;
  wire  xConnect_reset;
  wire  xConnect_io_in_req_ready;
  wire  xConnect_io_in_req_valid;
  wire [31:0] xConnect_io_in_req_bits_addr;
  wire [127:0] xConnect_io_in_req_bits_wdata;
  wire [2:0] xConnect_io_in_req_bits_cmd;
  wire  xConnect_io_in_resp_valid;
  wire [127:0] xConnect_io_in_resp_bits_rdata;
  wire  xConnect_io_out_mem_req_ready;
  wire  xConnect_io_out_mem_req_valid;
  wire [31:0] xConnect_io_out_mem_req_bits_addr;
  wire [127:0] xConnect_io_out_mem_req_bits_wdata;
  wire [2:0] xConnect_io_out_mem_req_bits_cmd;
  wire  xConnect_io_out_mem_resp_ready;
  wire  xConnect_io_out_mem_resp_valid;
  wire [2:0] xConnect_io_out_mem_resp_bits_cmd;
  wire [127:0] xConnect_io_out_mem_resp_bits_rdata;
  wire  xConnect_io_out_link_req_ready;
  wire  xConnect_io_out_link_req_valid;
  wire [31:0] xConnect_io_out_link_req_bits_addr;
  wire [127:0] xConnect_io_out_link_req_bits_wdata;
  wire  xConnect_io_out_link_resp_ready;
  wire  xConnect_io_out_link_resp_valid;
  wire [2:0] xConnect_io_out_link_resp_bits_cmd;
  wire [127:0] xConnect_io_out_link_resp_bits_rdata;
  wire  clint_clock;
  wire  clint_reset;
  wire  clint_io_in_aw_ready;
  wire  clint_io_in_aw_valid;
  wire [31:0] clint_io_in_aw_bits_addr;
  wire  clint_io_in_w_ready;
  wire  clint_io_in_w_valid;
  wire [7:0] clint_io_in_w_bits_strb;
  wire [63:0] clint_io_in_w_bits_data;
  wire  clint_io_in_b_ready;
  wire  clint_io_in_b_valid;
  wire  clint_io_in_ar_ready;
  wire  clint_io_in_ar_valid;
  wire [31:0] clint_io_in_ar_bits_addr;
  wire  clint_io_in_r_ready;
  wire  clint_io_in_r_valid;
  wire [63:0] clint_io_in_r_bits_data;
  wire  axi4XBar_clock;
  wire  axi4XBar_reset;
  wire  axi4XBar_io_in_0_aw_ready;
  wire  axi4XBar_io_in_0_aw_valid;
  wire [31:0] axi4XBar_io_in_0_aw_bits_addr;
  wire [2:0] axi4XBar_io_in_0_aw_bits_size;
  wire  axi4XBar_io_in_0_w_ready;
  wire  axi4XBar_io_in_0_w_valid;
  wire [63:0] axi4XBar_io_in_0_w_bits_data;
  wire  axi4XBar_io_in_0_w_bits_last;
  wire  axi4XBar_io_in_0_b_ready;
  wire  axi4XBar_io_in_0_b_valid;
  wire  axi4XBar_io_in_0_ar_ready;
  wire  axi4XBar_io_in_0_ar_valid;
  wire [31:0] axi4XBar_io_in_0_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_0_ar_bits_size;
  wire  axi4XBar_io_in_0_r_ready;
  wire  axi4XBar_io_in_0_r_valid;
  wire [63:0] axi4XBar_io_in_0_r_bits_data;
  wire  axi4XBar_io_in_0_r_bits_last;
  wire  axi4XBar_io_in_1_aw_ready;
  wire  axi4XBar_io_in_1_aw_valid;
  wire [31:0] axi4XBar_io_in_1_aw_bits_addr;
  wire [2:0] axi4XBar_io_in_1_aw_bits_size;
  wire  axi4XBar_io_in_1_w_ready;
  wire  axi4XBar_io_in_1_w_valid;
  wire [63:0] axi4XBar_io_in_1_w_bits_data;
  wire  axi4XBar_io_in_1_w_bits_last;
  wire  axi4XBar_io_in_1_b_ready;
  wire  axi4XBar_io_in_1_b_valid;
  wire  axi4XBar_io_in_1_ar_ready;
  wire  axi4XBar_io_in_1_ar_valid;
  wire [31:0] axi4XBar_io_in_1_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_1_ar_bits_size;
  wire  axi4XBar_io_in_1_r_ready;
  wire  axi4XBar_io_in_1_r_valid;
  wire [63:0] axi4XBar_io_in_1_r_bits_data;
  wire  axi4XBar_io_in_1_r_bits_last;
  wire  axi4XBar_io_in_2_aw_ready;
  wire  axi4XBar_io_in_2_aw_valid;
  wire [31:0] axi4XBar_io_in_2_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_2_aw_bits_id;
  wire [7:0] axi4XBar_io_in_2_aw_bits_len;
  wire [2:0] axi4XBar_io_in_2_aw_bits_size;
  wire [1:0] axi4XBar_io_in_2_aw_bits_burst;
  wire  axi4XBar_io_in_2_w_ready;
  wire  axi4XBar_io_in_2_w_valid;
  wire [7:0] axi4XBar_io_in_2_w_bits_strb;
  wire [63:0] axi4XBar_io_in_2_w_bits_data;
  wire  axi4XBar_io_in_2_b_ready;
  wire  axi4XBar_io_in_2_b_valid;
  wire  axi4XBar_io_in_2_ar_ready;
  wire  axi4XBar_io_in_2_ar_valid;
  wire [31:0] axi4XBar_io_in_2_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_2_ar_bits_size;
  wire  axi4XBar_io_in_2_r_ready;
  wire  axi4XBar_io_in_2_r_valid;
  wire [63:0] axi4XBar_io_in_2_r_bits_data;
  wire  axi4XBar_io_in_2_r_bits_last;
  wire  axi4XBar_io_in_3_aw_ready;
  wire  axi4XBar_io_in_3_aw_valid;
  wire [31:0] axi4XBar_io_in_3_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_3_aw_bits_id;
  wire [7:0] axi4XBar_io_in_3_aw_bits_len;
  wire [2:0] axi4XBar_io_in_3_aw_bits_size;
  wire [1:0] axi4XBar_io_in_3_aw_bits_burst;
  wire  axi4XBar_io_in_3_w_ready;
  wire  axi4XBar_io_in_3_w_valid;
  wire [7:0] axi4XBar_io_in_3_w_bits_strb;
  wire [63:0] axi4XBar_io_in_3_w_bits_data;
  wire  axi4XBar_io_in_3_b_ready;
  wire  axi4XBar_io_in_3_b_valid;
  wire  axi4XBar_io_in_3_ar_ready;
  wire  axi4XBar_io_in_3_ar_valid;
  wire [31:0] axi4XBar_io_in_3_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_3_ar_bits_size;
  wire  axi4XBar_io_in_3_r_ready;
  wire  axi4XBar_io_in_3_r_valid;
  wire [63:0] axi4XBar_io_in_3_r_bits_data;
  wire  axi4XBar_io_in_3_r_bits_last;
  wire  axi4XBar_io_in_4_aw_ready;
  wire  axi4XBar_io_in_4_aw_valid;
  wire [31:0] axi4XBar_io_in_4_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_4_aw_bits_id;
  wire [7:0] axi4XBar_io_in_4_aw_bits_len;
  wire [2:0] axi4XBar_io_in_4_aw_bits_size;
  wire [1:0] axi4XBar_io_in_4_aw_bits_burst;
  wire  axi4XBar_io_in_4_w_ready;
  wire  axi4XBar_io_in_4_w_valid;
  wire [7:0] axi4XBar_io_in_4_w_bits_strb;
  wire [63:0] axi4XBar_io_in_4_w_bits_data;
  wire  axi4XBar_io_in_4_b_ready;
  wire  axi4XBar_io_in_4_b_valid;
  wire  axi4XBar_io_in_4_ar_ready;
  wire  axi4XBar_io_in_4_ar_valid;
  wire [31:0] axi4XBar_io_in_4_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_4_ar_bits_size;
  wire  axi4XBar_io_in_4_r_ready;
  wire  axi4XBar_io_in_4_r_valid;
  wire [63:0] axi4XBar_io_in_4_r_bits_data;
  wire  axi4XBar_io_in_4_r_bits_last;
  wire  axi4XBar_io_in_5_aw_ready;
  wire  axi4XBar_io_in_5_aw_valid;
  wire [31:0] axi4XBar_io_in_5_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_5_aw_bits_id;
  wire [7:0] axi4XBar_io_in_5_aw_bits_len;
  wire [2:0] axi4XBar_io_in_5_aw_bits_size;
  wire [1:0] axi4XBar_io_in_5_aw_bits_burst;
  wire  axi4XBar_io_in_5_w_ready;
  wire  axi4XBar_io_in_5_w_valid;
  wire [7:0] axi4XBar_io_in_5_w_bits_strb;
  wire [63:0] axi4XBar_io_in_5_w_bits_data;
  wire  axi4XBar_io_in_5_b_ready;
  wire  axi4XBar_io_in_5_b_valid;
  wire  axi4XBar_io_in_5_ar_ready;
  wire  axi4XBar_io_in_5_ar_valid;
  wire [31:0] axi4XBar_io_in_5_ar_bits_addr;
  wire [2:0] axi4XBar_io_in_5_ar_bits_size;
  wire  axi4XBar_io_in_5_r_ready;
  wire  axi4XBar_io_in_5_r_valid;
  wire [63:0] axi4XBar_io_in_5_r_bits_data;
  wire  axi4XBar_io_in_5_r_bits_last;
  wire  axi4XBar_io_out_aw_ready;
  wire  axi4XBar_io_out_aw_valid;
  wire [31:0] axi4XBar_io_out_aw_bits_addr;
  wire [3:0] axi4XBar_io_out_aw_bits_id;
  wire [7:0] axi4XBar_io_out_aw_bits_len;
  wire [2:0] axi4XBar_io_out_aw_bits_size;
  wire [1:0] axi4XBar_io_out_aw_bits_burst;
  wire  axi4XBar_io_out_w_ready;
  wire  axi4XBar_io_out_w_valid;
  wire [7:0] axi4XBar_io_out_w_bits_strb;
  wire [63:0] axi4XBar_io_out_w_bits_data;
  wire  axi4XBar_io_out_w_bits_last;
  wire  axi4XBar_io_out_b_ready;
  wire  axi4XBar_io_out_b_valid;
  wire  axi4XBar_io_out_ar_ready;
  wire  axi4XBar_io_out_ar_valid;
  wire [31:0] axi4XBar_io_out_ar_bits_addr;
  wire [7:0] axi4XBar_io_out_ar_bits_len;
  wire [2:0] axi4XBar_io_out_ar_bits_size;
  wire [1:0] axi4XBar_io_out_ar_bits_burst;
  wire  axi4XBar_io_out_r_ready;
  wire  axi4XBar_io_out_r_valid;
  wire [63:0] axi4XBar_io_out_r_bits_data;
  wire  axi4XBar_io_out_r_bits_last;
  wire  mmioXBar_clock;
  wire  mmioXBar_reset;
  wire  mmioXBar_io_in_req_ready;
  wire  mmioXBar_io_in_req_valid;
  wire [31:0] mmioXBar_io_in_req_bits_addr;
  wire [63:0] mmioXBar_io_in_req_bits_wdata;
  wire [1:0] mmioXBar_io_in_req_bits_size;
  wire [2:0] mmioXBar_io_in_req_bits_cmd;
  wire  mmioXBar_io_in_resp_valid;
  wire [63:0] mmioXBar_io_in_resp_bits_rdata;
  wire  mmioXBar_io_out_0_req_ready;
  wire  mmioXBar_io_out_0_req_valid;
  wire [31:0] mmioXBar_io_out_0_req_bits_addr;
  wire [63:0] mmioXBar_io_out_0_req_bits_wdata;
  wire [1:0] mmioXBar_io_out_0_req_bits_size;
  wire [2:0] mmioXBar_io_out_0_req_bits_cmd;
  wire  mmioXBar_io_out_0_resp_ready;
  wire  mmioXBar_io_out_0_resp_valid;
  wire [63:0] mmioXBar_io_out_0_resp_bits_rdata;
  wire  mmioXBar_io_out_1_req_ready;
  wire  mmioXBar_io_out_1_req_valid;
  wire [31:0] mmioXBar_io_out_1_req_bits_addr;
  wire [63:0] mmioXBar_io_out_1_req_bits_wdata;
  wire [1:0] mmioXBar_io_out_1_req_bits_size;
  wire [2:0] mmioXBar_io_out_1_req_bits_cmd;
  wire  mmioXBar_io_out_1_resp_ready;
  wire  mmioXBar_io_out_1_resp_valid;
  wire [63:0] mmioXBar_io_out_1_resp_bits_rdata;
  wire  mmioXBar_io_out_2_req_ready;
  wire  mmioXBar_io_out_2_req_valid;
  wire [31:0] mmioXBar_io_out_2_req_bits_addr;
  wire [63:0] mmioXBar_io_out_2_req_bits_wdata;
  wire [1:0] mmioXBar_io_out_2_req_bits_size;
  wire [2:0] mmioXBar_io_out_2_req_bits_cmd;
  wire  mmioXBar_io_out_2_resp_ready;
  wire  mmioXBar_io_out_2_resp_valid;
  wire [63:0] mmioXBar_io_out_2_resp_bits_rdata;
  wire  mmioXBar_io_out_3_req_ready;
  wire  mmioXBar_io_out_3_req_valid;
  wire [31:0] mmioXBar_io_out_3_req_bits_addr;
  wire [63:0] mmioXBar_io_out_3_req_bits_wdata;
  wire [1:0] mmioXBar_io_out_3_req_bits_size;
  wire [2:0] mmioXBar_io_out_3_req_bits_cmd;
  wire  mmioXBar_io_out_3_resp_ready;
  wire  mmioXBar_io_out_3_resp_valid;
  wire [63:0] mmioXBar_io_out_3_resp_bits_rdata;
  wire  axiBridge_0_clock;
  wire  axiBridge_0_reset;
  wire  axiBridge_0_io_in_req_ready;
  wire  axiBridge_0_io_in_req_valid;
  wire [31:0] axiBridge_0_io_in_req_bits_addr;
  wire [127:0] axiBridge_0_io_in_req_bits_wdata;
  wire [2:0] axiBridge_0_io_in_req_bits_cmd;
  wire  axiBridge_0_io_in_resp_valid;
  wire [2:0] axiBridge_0_io_in_resp_bits_cmd;
  wire [127:0] axiBridge_0_io_in_resp_bits_rdata;
  wire  axiBridge_0_io_out_aw_ready;
  wire  axiBridge_0_io_out_aw_valid;
  wire [31:0] axiBridge_0_io_out_aw_bits_addr;
  wire [2:0] axiBridge_0_io_out_aw_bits_size;
  wire  axiBridge_0_io_out_w_ready;
  wire  axiBridge_0_io_out_w_valid;
  wire [63:0] axiBridge_0_io_out_w_bits_data;
  wire  axiBridge_0_io_out_w_bits_last;
  wire  axiBridge_0_io_out_b_ready;
  wire  axiBridge_0_io_out_b_valid;
  wire  axiBridge_0_io_out_ar_ready;
  wire  axiBridge_0_io_out_ar_valid;
  wire [31:0] axiBridge_0_io_out_ar_bits_addr;
  wire [2:0] axiBridge_0_io_out_ar_bits_size;
  wire  axiBridge_0_io_out_r_ready;
  wire  axiBridge_0_io_out_r_valid;
  wire [63:0] axiBridge_0_io_out_r_bits_data;
  wire  axiBridge_0_io_out_r_bits_last;
  wire  axiBridge_1_clock;
  wire  axiBridge_1_reset;
  wire  axiBridge_1_io_in_req_ready;
  wire  axiBridge_1_io_in_req_valid;
  wire [31:0] axiBridge_1_io_in_req_bits_addr;
  wire [127:0] axiBridge_1_io_in_req_bits_wdata;
  wire [2:0] axiBridge_1_io_in_req_bits_cmd;
  wire  axiBridge_1_io_in_resp_valid;
  wire [2:0] axiBridge_1_io_in_resp_bits_cmd;
  wire [127:0] axiBridge_1_io_in_resp_bits_rdata;
  wire  axiBridge_1_io_out_aw_ready;
  wire  axiBridge_1_io_out_aw_valid;
  wire [31:0] axiBridge_1_io_out_aw_bits_addr;
  wire [2:0] axiBridge_1_io_out_aw_bits_size;
  wire  axiBridge_1_io_out_w_ready;
  wire  axiBridge_1_io_out_w_valid;
  wire [63:0] axiBridge_1_io_out_w_bits_data;
  wire  axiBridge_1_io_out_w_bits_last;
  wire  axiBridge_1_io_out_b_ready;
  wire  axiBridge_1_io_out_b_valid;
  wire  axiBridge_1_io_out_ar_ready;
  wire  axiBridge_1_io_out_ar_valid;
  wire [31:0] axiBridge_1_io_out_ar_bits_addr;
  wire [2:0] axiBridge_1_io_out_ar_bits_size;
  wire  axiBridge_1_io_out_r_ready;
  wire  axiBridge_1_io_out_r_valid;
  wire [63:0] axiBridge_1_io_out_r_bits_data;
  wire  axiBridge_1_io_out_r_bits_last;
  wire  clint_io_in_toAXIbridge_clock;
  wire  clint_io_in_toAXIbridge_reset;
  wire  clint_io_in_toAXIbridge_io_in_req_ready;
  wire  clint_io_in_toAXIbridge_io_in_req_valid;
  wire [31:0] clint_io_in_toAXIbridge_io_in_req_bits_addr;
  wire [63:0] clint_io_in_toAXIbridge_io_in_req_bits_wdata;
  wire [1:0] clint_io_in_toAXIbridge_io_in_req_bits_size;
  wire [2:0] clint_io_in_toAXIbridge_io_in_req_bits_cmd;
  wire  clint_io_in_toAXIbridge_io_in_resp_ready;
  wire  clint_io_in_toAXIbridge_io_in_resp_valid;
  wire [63:0] clint_io_in_toAXIbridge_io_in_resp_bits_rdata;
  wire  clint_io_in_toAXIbridge_io_out_aw_ready;
  wire  clint_io_in_toAXIbridge_io_out_aw_valid;
  wire [31:0] clint_io_in_toAXIbridge_io_out_aw_bits_addr;
  wire  clint_io_in_toAXIbridge_io_out_w_ready;
  wire  clint_io_in_toAXIbridge_io_out_w_valid;
  wire [7:0] clint_io_in_toAXIbridge_io_out_w_bits_strb;
  wire [63:0] clint_io_in_toAXIbridge_io_out_w_bits_data;
  wire  clint_io_in_toAXIbridge_io_out_b_ready;
  wire  clint_io_in_toAXIbridge_io_out_b_valid;
  wire  clint_io_in_toAXIbridge_io_out_ar_ready;
  wire  clint_io_in_toAXIbridge_io_out_ar_valid;
  wire [31:0] clint_io_in_toAXIbridge_io_out_ar_bits_addr;
  wire  clint_io_in_toAXIbridge_io_out_r_ready;
  wire  clint_io_in_toAXIbridge_io_out_r_valid;
  wire [63:0] clint_io_in_toAXIbridge_io_out_r_bits_data;
  wire  axi4XBar_io_in_2_toAXIbridge_clock;
  wire  axi4XBar_io_in_2_toAXIbridge_reset;
  wire  axi4XBar_io_in_2_toAXIbridge_io_in_req_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_in_req_valid;
  wire [31:0] axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_addr;
  wire [63:0] axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_wdata;
  wire [1:0] axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_size;
  wire [2:0] axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_cmd;
  wire  axi4XBar_io_in_2_toAXIbridge_io_in_resp_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_in_resp_valid;
  wire [63:0] axi4XBar_io_in_2_toAXIbridge_io_in_resp_bits_rdata;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_aw_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_aw_valid;
  wire [31:0] axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_id;
  wire [7:0] axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_len;
  wire [2:0] axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_size;
  wire [1:0] axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_burst;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_w_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_w_valid;
  wire [7:0] axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_strb;
  wire [63:0] axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_data;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_last;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_b_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_b_valid;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_ar_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_ar_valid;
  wire [31:0] axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_addr;
  wire [3:0] axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_id;
  wire [7:0] axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_len;
  wire [2:0] axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_size;
  wire [1:0] axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_burst;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_r_ready;
  wire  axi4XBar_io_in_2_toAXIbridge_io_out_r_valid;
  wire [63:0] axi4XBar_io_in_2_toAXIbridge_io_out_r_bits_data;
  wire  axi4XBar_io_in_3_toAXIbridge_clock;
  wire  axi4XBar_io_in_3_toAXIbridge_reset;
  wire  axi4XBar_io_in_3_toAXIbridge_io_in_req_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_in_req_valid;
  wire [31:0] axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_addr;
  wire [63:0] axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_wdata;
  wire [1:0] axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_size;
  wire [2:0] axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_cmd;
  wire  axi4XBar_io_in_3_toAXIbridge_io_in_resp_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_in_resp_valid;
  wire [63:0] axi4XBar_io_in_3_toAXIbridge_io_in_resp_bits_rdata;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_aw_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_aw_valid;
  wire [31:0] axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_id;
  wire [7:0] axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_len;
  wire [2:0] axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_size;
  wire [1:0] axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_burst;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_w_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_w_valid;
  wire [7:0] axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_strb;
  wire [63:0] axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_data;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_last;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_b_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_b_valid;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_ar_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_ar_valid;
  wire [31:0] axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_addr;
  wire [3:0] axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_id;
  wire [7:0] axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_len;
  wire [2:0] axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_size;
  wire [1:0] axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_burst;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_r_ready;
  wire  axi4XBar_io_in_3_toAXIbridge_io_out_r_valid;
  wire [63:0] axi4XBar_io_in_3_toAXIbridge_io_out_r_bits_data;
  wire  axi4XBar_io_in_4_toAXIbridge_clock;
  wire  axi4XBar_io_in_4_toAXIbridge_reset;
  wire  axi4XBar_io_in_4_toAXIbridge_io_in_req_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_in_req_valid;
  wire [31:0] axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_addr;
  wire [63:0] axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_wdata;
  wire [1:0] axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_size;
  wire [2:0] axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_cmd;
  wire  axi4XBar_io_in_4_toAXIbridge_io_in_resp_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_in_resp_valid;
  wire [63:0] axi4XBar_io_in_4_toAXIbridge_io_in_resp_bits_rdata;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_aw_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_aw_valid;
  wire [31:0] axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_id;
  wire [7:0] axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_len;
  wire [2:0] axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_size;
  wire [1:0] axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_burst;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_w_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_w_valid;
  wire [7:0] axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_strb;
  wire [63:0] axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_data;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_last;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_b_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_b_valid;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_ar_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_ar_valid;
  wire [31:0] axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_addr;
  wire [3:0] axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_id;
  wire [7:0] axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_len;
  wire [2:0] axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_size;
  wire [1:0] axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_burst;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_r_ready;
  wire  axi4XBar_io_in_4_toAXIbridge_io_out_r_valid;
  wire [63:0] axi4XBar_io_in_4_toAXIbridge_io_out_r_bits_data;
  wire  axi4XBar_io_in_5_toAXIbridge_clock;
  wire  axi4XBar_io_in_5_toAXIbridge_reset;
  wire  axi4XBar_io_in_5_toAXIbridge_io_in_req_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_in_req_valid;
  wire [31:0] axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_addr;
  wire [63:0] axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_wdata;
  wire [1:0] axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_size;
  wire [2:0] axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_cmd;
  wire  axi4XBar_io_in_5_toAXIbridge_io_in_resp_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_in_resp_valid;
  wire [63:0] axi4XBar_io_in_5_toAXIbridge_io_in_resp_bits_rdata;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_aw_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_aw_valid;
  wire [31:0] axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_addr;
  wire [3:0] axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_id;
  wire [7:0] axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_len;
  wire [2:0] axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_size;
  wire [1:0] axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_burst;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_w_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_w_valid;
  wire [7:0] axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_strb;
  wire [63:0] axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_data;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_last;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_b_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_b_valid;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_ar_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_ar_valid;
  wire [31:0] axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_addr;
  wire [3:0] axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_id;
  wire [7:0] axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_len;
  wire [2:0] axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_size;
  wire [1:0] axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_burst;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_r_ready;
  wire  axi4XBar_io_in_5_toAXIbridge_io_out_r_valid;
  wire [63:0] axi4XBar_io_in_5_toAXIbridge_io_out_r_bits_data;
  ysyx_040656_CoreOverlay overlay (
    .clock(overlay_clock),
    .reset(overlay_reset),
    .io_imem_req_ready(overlay_io_imem_req_ready),
    .io_imem_req_valid(overlay_io_imem_req_valid),
    .io_imem_req_bits_addr(overlay_io_imem_req_bits_addr),
    .io_imem_req_bits_wdata(overlay_io_imem_req_bits_wdata),
    .io_imem_req_bits_cmd(overlay_io_imem_req_bits_cmd),
    .io_imem_resp_valid(overlay_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(overlay_io_imem_resp_bits_rdata),
    .io_dmem_req_ready(overlay_io_dmem_req_ready),
    .io_dmem_req_valid(overlay_io_dmem_req_valid),
    .io_dmem_req_bits_addr(overlay_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(overlay_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_cmd(overlay_io_dmem_req_bits_cmd),
    .io_dmem_resp_valid(overlay_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(overlay_io_dmem_resp_bits_rdata),
    .io_link_req_ready(overlay_io_link_req_ready),
    .io_link_req_valid(overlay_io_link_req_valid),
    .io_link_req_bits_addr(overlay_io_link_req_bits_addr),
    .io_link_req_bits_wdata(overlay_io_link_req_bits_wdata),
    .io_link_resp_valid(overlay_io_link_resp_valid),
    .io_link_resp_bits_cmd(overlay_io_link_resp_bits_cmd),
    .io_link_resp_bits_rdata(overlay_io_link_resp_bits_rdata),
    .io_immio_req_ready(overlay_io_immio_req_ready),
    .io_immio_req_valid(overlay_io_immio_req_valid),
    .io_immio_req_bits_addr(overlay_io_immio_req_bits_addr),
    .io_immio_req_bits_size(overlay_io_immio_req_bits_size),
    .io_immio_resp_valid(overlay_io_immio_resp_valid),
    .io_immio_resp_bits_rdata(overlay_io_immio_resp_bits_rdata),
    .io_dmmio_req_ready(overlay_io_dmmio_req_ready),
    .io_dmmio_req_valid(overlay_io_dmmio_req_valid),
    .io_dmmio_req_bits_addr(overlay_io_dmmio_req_bits_addr),
    .io_dmmio_req_bits_wdata(overlay_io_dmmio_req_bits_wdata),
    .io_dmmio_req_bits_size(overlay_io_dmmio_req_bits_size),
    .io_dmmio_req_bits_cmd(overlay_io_dmmio_req_bits_cmd),
    .io_dmmio_resp_valid(overlay_io_dmmio_resp_valid),
    .io_dmmio_resp_bits_rdata(overlay_io_dmmio_resp_bits_rdata),
    .io_sram0_rdata(overlay_io_sram0_rdata),
    .io_sram0_wen(overlay_io_sram0_wen),
    .io_sram0_addr(overlay_io_sram0_addr),
    .io_sram0_wdata(overlay_io_sram0_wdata),
    .io_sram1_rdata(overlay_io_sram1_rdata),
    .io_sram1_wen(overlay_io_sram1_wen),
    .io_sram1_addr(overlay_io_sram1_addr),
    .io_sram1_wdata(overlay_io_sram1_wdata),
    .io_sram2_rdata(overlay_io_sram2_rdata),
    .io_sram2_wen(overlay_io_sram2_wen),
    .io_sram2_addr(overlay_io_sram2_addr),
    .io_sram2_wdata(overlay_io_sram2_wdata),
    .io_sram3_rdata(overlay_io_sram3_rdata),
    .io_sram3_wen(overlay_io_sram3_wen),
    .io_sram3_addr(overlay_io_sram3_addr),
    .io_sram3_wdata(overlay_io_sram3_wdata),
    .io_sram4_rdata(overlay_io_sram4_rdata),
    .io_sram4_wen(overlay_io_sram4_wen),
    .io_sram4_addr(overlay_io_sram4_addr),
    .io_sram4_wdata(overlay_io_sram4_wdata),
    .io_sram5_rdata(overlay_io_sram5_rdata),
    .io_sram5_wen(overlay_io_sram5_wen),
    .io_sram5_addr(overlay_io_sram5_addr),
    .io_sram5_wdata(overlay_io_sram5_wdata),
    .io_sram6_rdata(overlay_io_sram6_rdata),
    .io_sram6_wen(overlay_io_sram6_wen),
    .io_sram6_addr(overlay_io_sram6_addr),
    .io_sram6_wdata(overlay_io_sram6_wdata),
    .io_sram7_rdata(overlay_io_sram7_rdata),
    .io_sram7_wen(overlay_io_sram7_wen),
    .io_sram7_addr(overlay_io_sram7_addr),
    .io_sram7_wdata(overlay_io_sram7_wdata)
  );
  ysyx_040656_XConnect xConnect (
    .clock(xConnect_clock),
    .reset(xConnect_reset),
    .io_in_req_ready(xConnect_io_in_req_ready),
    .io_in_req_valid(xConnect_io_in_req_valid),
    .io_in_req_bits_addr(xConnect_io_in_req_bits_addr),
    .io_in_req_bits_wdata(xConnect_io_in_req_bits_wdata),
    .io_in_req_bits_cmd(xConnect_io_in_req_bits_cmd),
    .io_in_resp_valid(xConnect_io_in_resp_valid),
    .io_in_resp_bits_rdata(xConnect_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(xConnect_io_out_mem_req_ready),
    .io_out_mem_req_valid(xConnect_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(xConnect_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_wdata(xConnect_io_out_mem_req_bits_wdata),
    .io_out_mem_req_bits_cmd(xConnect_io_out_mem_req_bits_cmd),
    .io_out_mem_resp_ready(xConnect_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(xConnect_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(xConnect_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(xConnect_io_out_mem_resp_bits_rdata),
    .io_out_link_req_ready(xConnect_io_out_link_req_ready),
    .io_out_link_req_valid(xConnect_io_out_link_req_valid),
    .io_out_link_req_bits_addr(xConnect_io_out_link_req_bits_addr),
    .io_out_link_req_bits_wdata(xConnect_io_out_link_req_bits_wdata),
    .io_out_link_resp_ready(xConnect_io_out_link_resp_ready),
    .io_out_link_resp_valid(xConnect_io_out_link_resp_valid),
    .io_out_link_resp_bits_cmd(xConnect_io_out_link_resp_bits_cmd),
    .io_out_link_resp_bits_rdata(xConnect_io_out_link_resp_bits_rdata)
  );
  ysyx_040656_AXI4CLINT clint (
    .clock(clint_clock),
    .reset(clint_reset),
    .io_in_aw_ready(clint_io_in_aw_ready),
    .io_in_aw_valid(clint_io_in_aw_valid),
    .io_in_aw_bits_addr(clint_io_in_aw_bits_addr),
    .io_in_w_ready(clint_io_in_w_ready),
    .io_in_w_valid(clint_io_in_w_valid),
    .io_in_w_bits_strb(clint_io_in_w_bits_strb),
    .io_in_w_bits_data(clint_io_in_w_bits_data),
    .io_in_b_ready(clint_io_in_b_ready),
    .io_in_b_valid(clint_io_in_b_valid),
    .io_in_ar_ready(clint_io_in_ar_ready),
    .io_in_ar_valid(clint_io_in_ar_valid),
    .io_in_ar_bits_addr(clint_io_in_ar_bits_addr),
    .io_in_r_ready(clint_io_in_r_ready),
    .io_in_r_valid(clint_io_in_r_valid),
    .io_in_r_bits_data(clint_io_in_r_bits_data)
  );
  ysyx_040656_AXI4XBar_Nto1 axi4XBar (
    .clock(axi4XBar_clock),
    .reset(axi4XBar_reset),
    .io_in_0_aw_ready(axi4XBar_io_in_0_aw_ready),
    .io_in_0_aw_valid(axi4XBar_io_in_0_aw_valid),
    .io_in_0_aw_bits_addr(axi4XBar_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_size(axi4XBar_io_in_0_aw_bits_size),
    .io_in_0_w_ready(axi4XBar_io_in_0_w_ready),
    .io_in_0_w_valid(axi4XBar_io_in_0_w_valid),
    .io_in_0_w_bits_data(axi4XBar_io_in_0_w_bits_data),
    .io_in_0_w_bits_last(axi4XBar_io_in_0_w_bits_last),
    .io_in_0_b_ready(axi4XBar_io_in_0_b_ready),
    .io_in_0_b_valid(axi4XBar_io_in_0_b_valid),
    .io_in_0_ar_ready(axi4XBar_io_in_0_ar_ready),
    .io_in_0_ar_valid(axi4XBar_io_in_0_ar_valid),
    .io_in_0_ar_bits_addr(axi4XBar_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_size(axi4XBar_io_in_0_ar_bits_size),
    .io_in_0_r_ready(axi4XBar_io_in_0_r_ready),
    .io_in_0_r_valid(axi4XBar_io_in_0_r_valid),
    .io_in_0_r_bits_data(axi4XBar_io_in_0_r_bits_data),
    .io_in_0_r_bits_last(axi4XBar_io_in_0_r_bits_last),
    .io_in_1_aw_ready(axi4XBar_io_in_1_aw_ready),
    .io_in_1_aw_valid(axi4XBar_io_in_1_aw_valid),
    .io_in_1_aw_bits_addr(axi4XBar_io_in_1_aw_bits_addr),
    .io_in_1_aw_bits_size(axi4XBar_io_in_1_aw_bits_size),
    .io_in_1_w_ready(axi4XBar_io_in_1_w_ready),
    .io_in_1_w_valid(axi4XBar_io_in_1_w_valid),
    .io_in_1_w_bits_data(axi4XBar_io_in_1_w_bits_data),
    .io_in_1_w_bits_last(axi4XBar_io_in_1_w_bits_last),
    .io_in_1_b_ready(axi4XBar_io_in_1_b_ready),
    .io_in_1_b_valid(axi4XBar_io_in_1_b_valid),
    .io_in_1_ar_ready(axi4XBar_io_in_1_ar_ready),
    .io_in_1_ar_valid(axi4XBar_io_in_1_ar_valid),
    .io_in_1_ar_bits_addr(axi4XBar_io_in_1_ar_bits_addr),
    .io_in_1_ar_bits_size(axi4XBar_io_in_1_ar_bits_size),
    .io_in_1_r_ready(axi4XBar_io_in_1_r_ready),
    .io_in_1_r_valid(axi4XBar_io_in_1_r_valid),
    .io_in_1_r_bits_data(axi4XBar_io_in_1_r_bits_data),
    .io_in_1_r_bits_last(axi4XBar_io_in_1_r_bits_last),
    .io_in_2_aw_ready(axi4XBar_io_in_2_aw_ready),
    .io_in_2_aw_valid(axi4XBar_io_in_2_aw_valid),
    .io_in_2_aw_bits_addr(axi4XBar_io_in_2_aw_bits_addr),
    .io_in_2_aw_bits_id(axi4XBar_io_in_2_aw_bits_id),
    .io_in_2_aw_bits_len(axi4XBar_io_in_2_aw_bits_len),
    .io_in_2_aw_bits_size(axi4XBar_io_in_2_aw_bits_size),
    .io_in_2_aw_bits_burst(axi4XBar_io_in_2_aw_bits_burst),
    .io_in_2_w_ready(axi4XBar_io_in_2_w_ready),
    .io_in_2_w_valid(axi4XBar_io_in_2_w_valid),
    .io_in_2_w_bits_strb(axi4XBar_io_in_2_w_bits_strb),
    .io_in_2_w_bits_data(axi4XBar_io_in_2_w_bits_data),
    .io_in_2_b_ready(axi4XBar_io_in_2_b_ready),
    .io_in_2_b_valid(axi4XBar_io_in_2_b_valid),
    .io_in_2_ar_ready(axi4XBar_io_in_2_ar_ready),
    .io_in_2_ar_valid(axi4XBar_io_in_2_ar_valid),
    .io_in_2_ar_bits_addr(axi4XBar_io_in_2_ar_bits_addr),
    .io_in_2_ar_bits_size(axi4XBar_io_in_2_ar_bits_size),
    .io_in_2_r_ready(axi4XBar_io_in_2_r_ready),
    .io_in_2_r_valid(axi4XBar_io_in_2_r_valid),
    .io_in_2_r_bits_data(axi4XBar_io_in_2_r_bits_data),
    .io_in_2_r_bits_last(axi4XBar_io_in_2_r_bits_last),
    .io_in_3_aw_ready(axi4XBar_io_in_3_aw_ready),
    .io_in_3_aw_valid(axi4XBar_io_in_3_aw_valid),
    .io_in_3_aw_bits_addr(axi4XBar_io_in_3_aw_bits_addr),
    .io_in_3_aw_bits_id(axi4XBar_io_in_3_aw_bits_id),
    .io_in_3_aw_bits_len(axi4XBar_io_in_3_aw_bits_len),
    .io_in_3_aw_bits_size(axi4XBar_io_in_3_aw_bits_size),
    .io_in_3_aw_bits_burst(axi4XBar_io_in_3_aw_bits_burst),
    .io_in_3_w_ready(axi4XBar_io_in_3_w_ready),
    .io_in_3_w_valid(axi4XBar_io_in_3_w_valid),
    .io_in_3_w_bits_strb(axi4XBar_io_in_3_w_bits_strb),
    .io_in_3_w_bits_data(axi4XBar_io_in_3_w_bits_data),
    .io_in_3_b_ready(axi4XBar_io_in_3_b_ready),
    .io_in_3_b_valid(axi4XBar_io_in_3_b_valid),
    .io_in_3_ar_ready(axi4XBar_io_in_3_ar_ready),
    .io_in_3_ar_valid(axi4XBar_io_in_3_ar_valid),
    .io_in_3_ar_bits_addr(axi4XBar_io_in_3_ar_bits_addr),
    .io_in_3_ar_bits_size(axi4XBar_io_in_3_ar_bits_size),
    .io_in_3_r_ready(axi4XBar_io_in_3_r_ready),
    .io_in_3_r_valid(axi4XBar_io_in_3_r_valid),
    .io_in_3_r_bits_data(axi4XBar_io_in_3_r_bits_data),
    .io_in_3_r_bits_last(axi4XBar_io_in_3_r_bits_last),
    .io_in_4_aw_ready(axi4XBar_io_in_4_aw_ready),
    .io_in_4_aw_valid(axi4XBar_io_in_4_aw_valid),
    .io_in_4_aw_bits_addr(axi4XBar_io_in_4_aw_bits_addr),
    .io_in_4_aw_bits_id(axi4XBar_io_in_4_aw_bits_id),
    .io_in_4_aw_bits_len(axi4XBar_io_in_4_aw_bits_len),
    .io_in_4_aw_bits_size(axi4XBar_io_in_4_aw_bits_size),
    .io_in_4_aw_bits_burst(axi4XBar_io_in_4_aw_bits_burst),
    .io_in_4_w_ready(axi4XBar_io_in_4_w_ready),
    .io_in_4_w_valid(axi4XBar_io_in_4_w_valid),
    .io_in_4_w_bits_strb(axi4XBar_io_in_4_w_bits_strb),
    .io_in_4_w_bits_data(axi4XBar_io_in_4_w_bits_data),
    .io_in_4_b_ready(axi4XBar_io_in_4_b_ready),
    .io_in_4_b_valid(axi4XBar_io_in_4_b_valid),
    .io_in_4_ar_ready(axi4XBar_io_in_4_ar_ready),
    .io_in_4_ar_valid(axi4XBar_io_in_4_ar_valid),
    .io_in_4_ar_bits_addr(axi4XBar_io_in_4_ar_bits_addr),
    .io_in_4_ar_bits_size(axi4XBar_io_in_4_ar_bits_size),
    .io_in_4_r_ready(axi4XBar_io_in_4_r_ready),
    .io_in_4_r_valid(axi4XBar_io_in_4_r_valid),
    .io_in_4_r_bits_data(axi4XBar_io_in_4_r_bits_data),
    .io_in_4_r_bits_last(axi4XBar_io_in_4_r_bits_last),
    .io_in_5_aw_ready(axi4XBar_io_in_5_aw_ready),
    .io_in_5_aw_valid(axi4XBar_io_in_5_aw_valid),
    .io_in_5_aw_bits_addr(axi4XBar_io_in_5_aw_bits_addr),
    .io_in_5_aw_bits_id(axi4XBar_io_in_5_aw_bits_id),
    .io_in_5_aw_bits_len(axi4XBar_io_in_5_aw_bits_len),
    .io_in_5_aw_bits_size(axi4XBar_io_in_5_aw_bits_size),
    .io_in_5_aw_bits_burst(axi4XBar_io_in_5_aw_bits_burst),
    .io_in_5_w_ready(axi4XBar_io_in_5_w_ready),
    .io_in_5_w_valid(axi4XBar_io_in_5_w_valid),
    .io_in_5_w_bits_strb(axi4XBar_io_in_5_w_bits_strb),
    .io_in_5_w_bits_data(axi4XBar_io_in_5_w_bits_data),
    .io_in_5_b_ready(axi4XBar_io_in_5_b_ready),
    .io_in_5_b_valid(axi4XBar_io_in_5_b_valid),
    .io_in_5_ar_ready(axi4XBar_io_in_5_ar_ready),
    .io_in_5_ar_valid(axi4XBar_io_in_5_ar_valid),
    .io_in_5_ar_bits_addr(axi4XBar_io_in_5_ar_bits_addr),
    .io_in_5_ar_bits_size(axi4XBar_io_in_5_ar_bits_size),
    .io_in_5_r_ready(axi4XBar_io_in_5_r_ready),
    .io_in_5_r_valid(axi4XBar_io_in_5_r_valid),
    .io_in_5_r_bits_data(axi4XBar_io_in_5_r_bits_data),
    .io_in_5_r_bits_last(axi4XBar_io_in_5_r_bits_last),
    .io_out_aw_ready(axi4XBar_io_out_aw_ready),
    .io_out_aw_valid(axi4XBar_io_out_aw_valid),
    .io_out_aw_bits_addr(axi4XBar_io_out_aw_bits_addr),
    .io_out_aw_bits_id(axi4XBar_io_out_aw_bits_id),
    .io_out_aw_bits_len(axi4XBar_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi4XBar_io_out_aw_bits_size),
    .io_out_aw_bits_burst(axi4XBar_io_out_aw_bits_burst),
    .io_out_w_ready(axi4XBar_io_out_w_ready),
    .io_out_w_valid(axi4XBar_io_out_w_valid),
    .io_out_w_bits_strb(axi4XBar_io_out_w_bits_strb),
    .io_out_w_bits_data(axi4XBar_io_out_w_bits_data),
    .io_out_w_bits_last(axi4XBar_io_out_w_bits_last),
    .io_out_b_ready(axi4XBar_io_out_b_ready),
    .io_out_b_valid(axi4XBar_io_out_b_valid),
    .io_out_ar_ready(axi4XBar_io_out_ar_ready),
    .io_out_ar_valid(axi4XBar_io_out_ar_valid),
    .io_out_ar_bits_addr(axi4XBar_io_out_ar_bits_addr),
    .io_out_ar_bits_len(axi4XBar_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi4XBar_io_out_ar_bits_size),
    .io_out_ar_bits_burst(axi4XBar_io_out_ar_bits_burst),
    .io_out_r_ready(axi4XBar_io_out_r_ready),
    .io_out_r_valid(axi4XBar_io_out_r_valid),
    .io_out_r_bits_data(axi4XBar_io_out_r_bits_data),
    .io_out_r_bits_last(axi4XBar_io_out_r_bits_last)
  );
  ysyx_040656_CoreLinkXBar mmioXBar (
    .clock(mmioXBar_clock),
    .reset(mmioXBar_reset),
    .io_in_req_ready(mmioXBar_io_in_req_ready),
    .io_in_req_valid(mmioXBar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXBar_io_in_req_bits_addr),
    .io_in_req_bits_wdata(mmioXBar_io_in_req_bits_wdata),
    .io_in_req_bits_size(mmioXBar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXBar_io_in_req_bits_cmd),
    .io_in_resp_valid(mmioXBar_io_in_resp_valid),
    .io_in_resp_bits_rdata(mmioXBar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXBar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXBar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXBar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_wdata(mmioXBar_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_size(mmioXBar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(mmioXBar_io_out_0_req_bits_cmd),
    .io_out_0_resp_ready(mmioXBar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXBar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXBar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXBar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXBar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXBar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_wdata(mmioXBar_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_size(mmioXBar_io_out_1_req_bits_size),
    .io_out_1_req_bits_cmd(mmioXBar_io_out_1_req_bits_cmd),
    .io_out_1_resp_ready(mmioXBar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXBar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXBar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXBar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXBar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXBar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_wdata(mmioXBar_io_out_2_req_bits_wdata),
    .io_out_2_req_bits_size(mmioXBar_io_out_2_req_bits_size),
    .io_out_2_req_bits_cmd(mmioXBar_io_out_2_req_bits_cmd),
    .io_out_2_resp_ready(mmioXBar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXBar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(mmioXBar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(mmioXBar_io_out_3_req_ready),
    .io_out_3_req_valid(mmioXBar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(mmioXBar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_wdata(mmioXBar_io_out_3_req_bits_wdata),
    .io_out_3_req_bits_size(mmioXBar_io_out_3_req_bits_size),
    .io_out_3_req_bits_cmd(mmioXBar_io_out_3_req_bits_cmd),
    .io_out_3_resp_ready(mmioXBar_io_out_3_resp_ready),
    .io_out_3_resp_valid(mmioXBar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(mmioXBar_io_out_3_resp_bits_rdata)
  );
  ysyx_040656_AXI4Bridge axiBridge_0 (
    .clock(axiBridge_0_clock),
    .reset(axiBridge_0_reset),
    .io_in_req_ready(axiBridge_0_io_in_req_ready),
    .io_in_req_valid(axiBridge_0_io_in_req_valid),
    .io_in_req_bits_addr(axiBridge_0_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axiBridge_0_io_in_req_bits_wdata),
    .io_in_req_bits_cmd(axiBridge_0_io_in_req_bits_cmd),
    .io_in_resp_valid(axiBridge_0_io_in_resp_valid),
    .io_in_resp_bits_cmd(axiBridge_0_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(axiBridge_0_io_in_resp_bits_rdata),
    .io_out_aw_ready(axiBridge_0_io_out_aw_ready),
    .io_out_aw_valid(axiBridge_0_io_out_aw_valid),
    .io_out_aw_bits_addr(axiBridge_0_io_out_aw_bits_addr),
    .io_out_aw_bits_size(axiBridge_0_io_out_aw_bits_size),
    .io_out_w_ready(axiBridge_0_io_out_w_ready),
    .io_out_w_valid(axiBridge_0_io_out_w_valid),
    .io_out_w_bits_data(axiBridge_0_io_out_w_bits_data),
    .io_out_w_bits_last(axiBridge_0_io_out_w_bits_last),
    .io_out_b_ready(axiBridge_0_io_out_b_ready),
    .io_out_b_valid(axiBridge_0_io_out_b_valid),
    .io_out_ar_ready(axiBridge_0_io_out_ar_ready),
    .io_out_ar_valid(axiBridge_0_io_out_ar_valid),
    .io_out_ar_bits_addr(axiBridge_0_io_out_ar_bits_addr),
    .io_out_ar_bits_size(axiBridge_0_io_out_ar_bits_size),
    .io_out_r_ready(axiBridge_0_io_out_r_ready),
    .io_out_r_valid(axiBridge_0_io_out_r_valid),
    .io_out_r_bits_data(axiBridge_0_io_out_r_bits_data),
    .io_out_r_bits_last(axiBridge_0_io_out_r_bits_last)
  );
  ysyx_040656_AXI4Bridge axiBridge_1 (
    .clock(axiBridge_1_clock),
    .reset(axiBridge_1_reset),
    .io_in_req_ready(axiBridge_1_io_in_req_ready),
    .io_in_req_valid(axiBridge_1_io_in_req_valid),
    .io_in_req_bits_addr(axiBridge_1_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axiBridge_1_io_in_req_bits_wdata),
    .io_in_req_bits_cmd(axiBridge_1_io_in_req_bits_cmd),
    .io_in_resp_valid(axiBridge_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(axiBridge_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(axiBridge_1_io_in_resp_bits_rdata),
    .io_out_aw_ready(axiBridge_1_io_out_aw_ready),
    .io_out_aw_valid(axiBridge_1_io_out_aw_valid),
    .io_out_aw_bits_addr(axiBridge_1_io_out_aw_bits_addr),
    .io_out_aw_bits_size(axiBridge_1_io_out_aw_bits_size),
    .io_out_w_ready(axiBridge_1_io_out_w_ready),
    .io_out_w_valid(axiBridge_1_io_out_w_valid),
    .io_out_w_bits_data(axiBridge_1_io_out_w_bits_data),
    .io_out_w_bits_last(axiBridge_1_io_out_w_bits_last),
    .io_out_b_ready(axiBridge_1_io_out_b_ready),
    .io_out_b_valid(axiBridge_1_io_out_b_valid),
    .io_out_ar_ready(axiBridge_1_io_out_ar_ready),
    .io_out_ar_valid(axiBridge_1_io_out_ar_valid),
    .io_out_ar_bits_addr(axiBridge_1_io_out_ar_bits_addr),
    .io_out_ar_bits_size(axiBridge_1_io_out_ar_bits_size),
    .io_out_r_ready(axiBridge_1_io_out_r_ready),
    .io_out_r_valid(axiBridge_1_io_out_r_valid),
    .io_out_r_bits_data(axiBridge_1_io_out_r_bits_data),
    .io_out_r_bits_last(axiBridge_1_io_out_r_bits_last)
  );
  ysyx_040656_CoreLink2AXI4 clint_io_in_toAXIbridge (
    .clock(clint_io_in_toAXIbridge_clock),
    .reset(clint_io_in_toAXIbridge_reset),
    .io_in_req_ready(clint_io_in_toAXIbridge_io_in_req_ready),
    .io_in_req_valid(clint_io_in_toAXIbridge_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_toAXIbridge_io_in_req_bits_addr),
    .io_in_req_bits_wdata(clint_io_in_toAXIbridge_io_in_req_bits_wdata),
    .io_in_req_bits_size(clint_io_in_toAXIbridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(clint_io_in_toAXIbridge_io_in_req_bits_cmd),
    .io_in_resp_ready(clint_io_in_toAXIbridge_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_toAXIbridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_toAXIbridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(clint_io_in_toAXIbridge_io_out_aw_ready),
    .io_out_aw_valid(clint_io_in_toAXIbridge_io_out_aw_valid),
    .io_out_aw_bits_addr(clint_io_in_toAXIbridge_io_out_aw_bits_addr),
    .io_out_w_ready(clint_io_in_toAXIbridge_io_out_w_ready),
    .io_out_w_valid(clint_io_in_toAXIbridge_io_out_w_valid),
    .io_out_w_bits_strb(clint_io_in_toAXIbridge_io_out_w_bits_strb),
    .io_out_w_bits_data(clint_io_in_toAXIbridge_io_out_w_bits_data),
    .io_out_b_ready(clint_io_in_toAXIbridge_io_out_b_ready),
    .io_out_b_valid(clint_io_in_toAXIbridge_io_out_b_valid),
    .io_out_ar_ready(clint_io_in_toAXIbridge_io_out_ar_ready),
    .io_out_ar_valid(clint_io_in_toAXIbridge_io_out_ar_valid),
    .io_out_ar_bits_addr(clint_io_in_toAXIbridge_io_out_ar_bits_addr),
    .io_out_r_ready(clint_io_in_toAXIbridge_io_out_r_ready),
    .io_out_r_valid(clint_io_in_toAXIbridge_io_out_r_valid),
    .io_out_r_bits_data(clint_io_in_toAXIbridge_io_out_r_bits_data)
  );
  ysyx_040656_CoreLink2AXI4_1 axi4XBar_io_in_2_toAXIbridge (
    .clock(axi4XBar_io_in_2_toAXIbridge_clock),
    .reset(axi4XBar_io_in_2_toAXIbridge_reset),
    .io_in_req_ready(axi4XBar_io_in_2_toAXIbridge_io_in_req_ready),
    .io_in_req_valid(axi4XBar_io_in_2_toAXIbridge_io_in_req_valid),
    .io_in_req_bits_addr(axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_wdata),
    .io_in_req_bits_size(axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_cmd),
    .io_in_resp_ready(axi4XBar_io_in_2_toAXIbridge_io_in_resp_ready),
    .io_in_resp_valid(axi4XBar_io_in_2_toAXIbridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(axi4XBar_io_in_2_toAXIbridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(axi4XBar_io_in_2_toAXIbridge_io_out_aw_ready),
    .io_out_aw_valid(axi4XBar_io_in_2_toAXIbridge_io_out_aw_valid),
    .io_out_aw_bits_addr(axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_addr),
    .io_out_aw_bits_id(axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_id),
    .io_out_aw_bits_len(axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_burst),
    .io_out_w_ready(axi4XBar_io_in_2_toAXIbridge_io_out_w_ready),
    .io_out_w_valid(axi4XBar_io_in_2_toAXIbridge_io_out_w_valid),
    .io_out_w_bits_strb(axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_strb),
    .io_out_w_bits_data(axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_data),
    .io_out_w_bits_last(axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_last),
    .io_out_b_ready(axi4XBar_io_in_2_toAXIbridge_io_out_b_ready),
    .io_out_b_valid(axi4XBar_io_in_2_toAXIbridge_io_out_b_valid),
    .io_out_ar_ready(axi4XBar_io_in_2_toAXIbridge_io_out_ar_ready),
    .io_out_ar_valid(axi4XBar_io_in_2_toAXIbridge_io_out_ar_valid),
    .io_out_ar_bits_addr(axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_addr),
    .io_out_ar_bits_id(axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_id),
    .io_out_ar_bits_len(axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_burst),
    .io_out_r_ready(axi4XBar_io_in_2_toAXIbridge_io_out_r_ready),
    .io_out_r_valid(axi4XBar_io_in_2_toAXIbridge_io_out_r_valid),
    .io_out_r_bits_data(axi4XBar_io_in_2_toAXIbridge_io_out_r_bits_data)
  );
  ysyx_040656_CoreLink2AXI4_1 axi4XBar_io_in_3_toAXIbridge (
    .clock(axi4XBar_io_in_3_toAXIbridge_clock),
    .reset(axi4XBar_io_in_3_toAXIbridge_reset),
    .io_in_req_ready(axi4XBar_io_in_3_toAXIbridge_io_in_req_ready),
    .io_in_req_valid(axi4XBar_io_in_3_toAXIbridge_io_in_req_valid),
    .io_in_req_bits_addr(axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_wdata),
    .io_in_req_bits_size(axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_cmd),
    .io_in_resp_ready(axi4XBar_io_in_3_toAXIbridge_io_in_resp_ready),
    .io_in_resp_valid(axi4XBar_io_in_3_toAXIbridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(axi4XBar_io_in_3_toAXIbridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(axi4XBar_io_in_3_toAXIbridge_io_out_aw_ready),
    .io_out_aw_valid(axi4XBar_io_in_3_toAXIbridge_io_out_aw_valid),
    .io_out_aw_bits_addr(axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_addr),
    .io_out_aw_bits_id(axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_id),
    .io_out_aw_bits_len(axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_burst),
    .io_out_w_ready(axi4XBar_io_in_3_toAXIbridge_io_out_w_ready),
    .io_out_w_valid(axi4XBar_io_in_3_toAXIbridge_io_out_w_valid),
    .io_out_w_bits_strb(axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_strb),
    .io_out_w_bits_data(axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_data),
    .io_out_w_bits_last(axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_last),
    .io_out_b_ready(axi4XBar_io_in_3_toAXIbridge_io_out_b_ready),
    .io_out_b_valid(axi4XBar_io_in_3_toAXIbridge_io_out_b_valid),
    .io_out_ar_ready(axi4XBar_io_in_3_toAXIbridge_io_out_ar_ready),
    .io_out_ar_valid(axi4XBar_io_in_3_toAXIbridge_io_out_ar_valid),
    .io_out_ar_bits_addr(axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_addr),
    .io_out_ar_bits_id(axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_id),
    .io_out_ar_bits_len(axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_burst),
    .io_out_r_ready(axi4XBar_io_in_3_toAXIbridge_io_out_r_ready),
    .io_out_r_valid(axi4XBar_io_in_3_toAXIbridge_io_out_r_valid),
    .io_out_r_bits_data(axi4XBar_io_in_3_toAXIbridge_io_out_r_bits_data)
  );
  ysyx_040656_CoreLink2AXI4_1 axi4XBar_io_in_4_toAXIbridge (
    .clock(axi4XBar_io_in_4_toAXIbridge_clock),
    .reset(axi4XBar_io_in_4_toAXIbridge_reset),
    .io_in_req_ready(axi4XBar_io_in_4_toAXIbridge_io_in_req_ready),
    .io_in_req_valid(axi4XBar_io_in_4_toAXIbridge_io_in_req_valid),
    .io_in_req_bits_addr(axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_wdata),
    .io_in_req_bits_size(axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_cmd),
    .io_in_resp_ready(axi4XBar_io_in_4_toAXIbridge_io_in_resp_ready),
    .io_in_resp_valid(axi4XBar_io_in_4_toAXIbridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(axi4XBar_io_in_4_toAXIbridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(axi4XBar_io_in_4_toAXIbridge_io_out_aw_ready),
    .io_out_aw_valid(axi4XBar_io_in_4_toAXIbridge_io_out_aw_valid),
    .io_out_aw_bits_addr(axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_addr),
    .io_out_aw_bits_id(axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_id),
    .io_out_aw_bits_len(axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_burst),
    .io_out_w_ready(axi4XBar_io_in_4_toAXIbridge_io_out_w_ready),
    .io_out_w_valid(axi4XBar_io_in_4_toAXIbridge_io_out_w_valid),
    .io_out_w_bits_strb(axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_strb),
    .io_out_w_bits_data(axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_data),
    .io_out_w_bits_last(axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_last),
    .io_out_b_ready(axi4XBar_io_in_4_toAXIbridge_io_out_b_ready),
    .io_out_b_valid(axi4XBar_io_in_4_toAXIbridge_io_out_b_valid),
    .io_out_ar_ready(axi4XBar_io_in_4_toAXIbridge_io_out_ar_ready),
    .io_out_ar_valid(axi4XBar_io_in_4_toAXIbridge_io_out_ar_valid),
    .io_out_ar_bits_addr(axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_addr),
    .io_out_ar_bits_id(axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_id),
    .io_out_ar_bits_len(axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_burst),
    .io_out_r_ready(axi4XBar_io_in_4_toAXIbridge_io_out_r_ready),
    .io_out_r_valid(axi4XBar_io_in_4_toAXIbridge_io_out_r_valid),
    .io_out_r_bits_data(axi4XBar_io_in_4_toAXIbridge_io_out_r_bits_data)
  );
  ysyx_040656_CoreLink2AXI4_1 axi4XBar_io_in_5_toAXIbridge (
    .clock(axi4XBar_io_in_5_toAXIbridge_clock),
    .reset(axi4XBar_io_in_5_toAXIbridge_reset),
    .io_in_req_ready(axi4XBar_io_in_5_toAXIbridge_io_in_req_ready),
    .io_in_req_valid(axi4XBar_io_in_5_toAXIbridge_io_in_req_valid),
    .io_in_req_bits_addr(axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_addr),
    .io_in_req_bits_wdata(axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_wdata),
    .io_in_req_bits_size(axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_cmd),
    .io_in_resp_ready(axi4XBar_io_in_5_toAXIbridge_io_in_resp_ready),
    .io_in_resp_valid(axi4XBar_io_in_5_toAXIbridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(axi4XBar_io_in_5_toAXIbridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(axi4XBar_io_in_5_toAXIbridge_io_out_aw_ready),
    .io_out_aw_valid(axi4XBar_io_in_5_toAXIbridge_io_out_aw_valid),
    .io_out_aw_bits_addr(axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_addr),
    .io_out_aw_bits_id(axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_id),
    .io_out_aw_bits_len(axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_len),
    .io_out_aw_bits_size(axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_size),
    .io_out_aw_bits_burst(axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_burst),
    .io_out_w_ready(axi4XBar_io_in_5_toAXIbridge_io_out_w_ready),
    .io_out_w_valid(axi4XBar_io_in_5_toAXIbridge_io_out_w_valid),
    .io_out_w_bits_strb(axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_strb),
    .io_out_w_bits_data(axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_data),
    .io_out_w_bits_last(axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_last),
    .io_out_b_ready(axi4XBar_io_in_5_toAXIbridge_io_out_b_ready),
    .io_out_b_valid(axi4XBar_io_in_5_toAXIbridge_io_out_b_valid),
    .io_out_ar_ready(axi4XBar_io_in_5_toAXIbridge_io_out_ar_ready),
    .io_out_ar_valid(axi4XBar_io_in_5_toAXIbridge_io_out_ar_valid),
    .io_out_ar_bits_addr(axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_addr),
    .io_out_ar_bits_id(axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_id),
    .io_out_ar_bits_len(axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_size),
    .io_out_ar_bits_burst(axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_burst),
    .io_out_r_ready(axi4XBar_io_in_5_toAXIbridge_io_out_r_ready),
    .io_out_r_valid(axi4XBar_io_in_5_toAXIbridge_io_out_r_valid),
    .io_out_r_bits_data(axi4XBar_io_in_5_toAXIbridge_io_out_r_bits_data)
  );
  assign io_master_arvalid = axi4XBar_io_out_ar_valid;
  assign io_master_araddr = axi4XBar_io_out_ar_bits_addr;
  assign io_master_arid = 4'h0;
  assign io_master_arlen = axi4XBar_io_out_ar_bits_len;
  assign io_master_arsize = axi4XBar_io_out_ar_bits_size;
  assign io_master_arburst = axi4XBar_io_out_ar_bits_burst;
  assign io_master_rready = axi4XBar_io_out_r_ready;
  assign io_master_awvalid = axi4XBar_io_out_aw_valid;
  assign io_master_awaddr = axi4XBar_io_out_aw_bits_addr;
  assign io_master_awid = axi4XBar_io_out_aw_bits_id;
  assign io_master_awlen = axi4XBar_io_out_aw_bits_len;
  assign io_master_awsize = axi4XBar_io_out_aw_bits_size;
  assign io_master_awburst = axi4XBar_io_out_aw_bits_burst;
  assign io_master_wvalid = axi4XBar_io_out_w_valid;
  assign io_master_wdata = axi4XBar_io_out_w_bits_data;
  assign io_master_wstrb = axi4XBar_io_out_w_bits_strb;
  assign io_master_wlast = axi4XBar_io_out_w_bits_last;
  assign io_master_bready = axi4XBar_io_out_b_ready;
  assign io_slave_arready = 1'h0;
  assign io_slave_rvalid = 1'h0;
  assign io_slave_rresp = 2'h0;
  assign io_slave_rdata = 64'h0;
  assign io_slave_rlast = 1'h0;
  assign io_slave_rid = 4'h0;
  assign io_slave_awready = 1'h0;
  assign io_slave_wready = 1'h0;
  assign io_slave_bvalid = 1'h0;
  assign io_slave_bresp = 2'h0;
  assign io_slave_bid = 4'h0;
  assign io_sram0_wen = overlay_io_sram0_wen;
  assign io_sram0_cen = 1'h0;
  assign io_sram0_addr = overlay_io_sram0_addr;
  assign io_sram0_wdata = overlay_io_sram0_wdata;
  assign io_sram0_wmask = 128'h0;
  assign io_sram1_wen = overlay_io_sram1_wen;
  assign io_sram1_cen = 1'h0;
  assign io_sram1_addr = overlay_io_sram1_addr;
  assign io_sram1_wdata = overlay_io_sram1_wdata;
  assign io_sram1_wmask = 128'h0;
  assign io_sram2_wen = overlay_io_sram2_wen;
  assign io_sram2_cen = 1'h0;
  assign io_sram2_addr = overlay_io_sram2_addr;
  assign io_sram2_wdata = overlay_io_sram2_wdata;
  assign io_sram2_wmask = 128'h0;
  assign io_sram3_wen = overlay_io_sram3_wen;
  assign io_sram3_cen = 1'h0;
  assign io_sram3_addr = overlay_io_sram3_addr;
  assign io_sram3_wdata = overlay_io_sram3_wdata;
  assign io_sram3_wmask = 128'h0;
  assign io_sram4_wen = overlay_io_sram4_wen;
  assign io_sram4_cen = 1'h0;
  assign io_sram4_addr = overlay_io_sram4_addr;
  assign io_sram4_wdata = overlay_io_sram4_wdata;
  assign io_sram4_wmask = 128'h0;
  assign io_sram5_wen = overlay_io_sram5_wen;
  assign io_sram5_cen = 1'h0;
  assign io_sram5_addr = overlay_io_sram5_addr;
  assign io_sram5_wdata = overlay_io_sram5_wdata;
  assign io_sram5_wmask = 128'h0;
  assign io_sram6_wen = overlay_io_sram6_wen;
  assign io_sram6_cen = 1'h0;
  assign io_sram6_addr = overlay_io_sram6_addr;
  assign io_sram6_wdata = overlay_io_sram6_wdata;
  assign io_sram6_wmask = 128'h0;
  assign io_sram7_wen = overlay_io_sram7_wen;
  assign io_sram7_cen = 1'h0;
  assign io_sram7_addr = overlay_io_sram7_addr;
  assign io_sram7_wdata = overlay_io_sram7_wdata;
  assign io_sram7_wmask = 128'h0;
  assign overlay_clock = clock;
  assign overlay_reset = reset;
  assign overlay_io_imem_req_ready = xConnect_io_in_req_ready;
  assign overlay_io_imem_resp_valid = xConnect_io_in_resp_valid;
  assign overlay_io_imem_resp_bits_rdata = xConnect_io_in_resp_bits_rdata;
  assign overlay_io_dmem_req_ready = axiBridge_1_io_in_req_ready;
  assign overlay_io_dmem_resp_valid = axiBridge_1_io_in_resp_valid;
  assign overlay_io_dmem_resp_bits_rdata = axiBridge_1_io_in_resp_bits_rdata;
  assign overlay_io_link_req_valid = xConnect_io_out_link_req_valid;
  assign overlay_io_link_req_bits_addr = xConnect_io_out_link_req_bits_addr;
  assign overlay_io_link_req_bits_wdata = xConnect_io_out_link_req_bits_wdata;
  assign overlay_io_immio_req_ready = axi4XBar_io_in_2_toAXIbridge_io_in_req_ready;
  assign overlay_io_immio_resp_valid = axi4XBar_io_in_2_toAXIbridge_io_in_resp_valid;
  assign overlay_io_immio_resp_bits_rdata = axi4XBar_io_in_2_toAXIbridge_io_in_resp_bits_rdata;
  assign overlay_io_dmmio_req_ready = mmioXBar_io_in_req_ready;
  assign overlay_io_dmmio_resp_valid = mmioXBar_io_in_resp_valid;
  assign overlay_io_dmmio_resp_bits_rdata = mmioXBar_io_in_resp_bits_rdata;
  assign overlay_io_sram0_rdata = io_sram0_rdata;
  assign overlay_io_sram1_rdata = io_sram1_rdata;
  assign overlay_io_sram2_rdata = io_sram2_rdata;
  assign overlay_io_sram3_rdata = io_sram3_rdata;
  assign overlay_io_sram4_rdata = io_sram4_rdata;
  assign overlay_io_sram5_rdata = io_sram5_rdata;
  assign overlay_io_sram6_rdata = io_sram6_rdata;
  assign overlay_io_sram7_rdata = io_sram7_rdata;
  assign xConnect_clock = clock;
  assign xConnect_reset = reset;
  assign xConnect_io_in_req_valid = overlay_io_imem_req_valid;
  assign xConnect_io_in_req_bits_addr = overlay_io_imem_req_bits_addr;
  assign xConnect_io_in_req_bits_wdata = overlay_io_imem_req_bits_wdata;
  assign xConnect_io_in_req_bits_cmd = overlay_io_imem_req_bits_cmd;
  assign xConnect_io_out_mem_req_ready = axiBridge_0_io_in_req_ready;
  assign xConnect_io_out_mem_resp_valid = axiBridge_0_io_in_resp_valid;
  assign xConnect_io_out_mem_resp_bits_cmd = axiBridge_0_io_in_resp_bits_cmd;
  assign xConnect_io_out_mem_resp_bits_rdata = axiBridge_0_io_in_resp_bits_rdata;
  assign xConnect_io_out_link_req_ready = overlay_io_link_req_ready;
  assign xConnect_io_out_link_resp_valid = overlay_io_link_resp_valid;
  assign xConnect_io_out_link_resp_bits_cmd = overlay_io_link_resp_bits_cmd;
  assign xConnect_io_out_link_resp_bits_rdata = overlay_io_link_resp_bits_rdata;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_in_aw_valid = clint_io_in_toAXIbridge_io_out_aw_valid;
  assign clint_io_in_aw_bits_addr = clint_io_in_toAXIbridge_io_out_aw_bits_addr;
  assign clint_io_in_w_valid = clint_io_in_toAXIbridge_io_out_w_valid;
  assign clint_io_in_w_bits_strb = clint_io_in_toAXIbridge_io_out_w_bits_strb;
  assign clint_io_in_w_bits_data = clint_io_in_toAXIbridge_io_out_w_bits_data;
  assign clint_io_in_b_ready = clint_io_in_toAXIbridge_io_out_b_ready;
  assign clint_io_in_ar_valid = clint_io_in_toAXIbridge_io_out_ar_valid;
  assign clint_io_in_ar_bits_addr = clint_io_in_toAXIbridge_io_out_ar_bits_addr;
  assign clint_io_in_r_ready = clint_io_in_toAXIbridge_io_out_r_ready;
  assign axi4XBar_clock = clock;
  assign axi4XBar_reset = reset;
  assign axi4XBar_io_in_0_aw_valid = axiBridge_0_io_out_aw_valid;
  assign axi4XBar_io_in_0_aw_bits_addr = axiBridge_0_io_out_aw_bits_addr;
  assign axi4XBar_io_in_0_aw_bits_size = axiBridge_0_io_out_aw_bits_size;
  assign axi4XBar_io_in_0_w_valid = axiBridge_0_io_out_w_valid;
  assign axi4XBar_io_in_0_w_bits_data = axiBridge_0_io_out_w_bits_data;
  assign axi4XBar_io_in_0_w_bits_last = axiBridge_0_io_out_w_bits_last;
  assign axi4XBar_io_in_0_b_ready = axiBridge_0_io_out_b_ready;
  assign axi4XBar_io_in_0_ar_valid = axiBridge_0_io_out_ar_valid;
  assign axi4XBar_io_in_0_ar_bits_addr = axiBridge_0_io_out_ar_bits_addr;
  assign axi4XBar_io_in_0_ar_bits_size = axiBridge_0_io_out_ar_bits_size;
  assign axi4XBar_io_in_0_r_ready = axiBridge_0_io_out_r_ready;
  assign axi4XBar_io_in_1_aw_valid = axiBridge_1_io_out_aw_valid;
  assign axi4XBar_io_in_1_aw_bits_addr = axiBridge_1_io_out_aw_bits_addr;
  assign axi4XBar_io_in_1_aw_bits_size = axiBridge_1_io_out_aw_bits_size;
  assign axi4XBar_io_in_1_w_valid = axiBridge_1_io_out_w_valid;
  assign axi4XBar_io_in_1_w_bits_data = axiBridge_1_io_out_w_bits_data;
  assign axi4XBar_io_in_1_w_bits_last = axiBridge_1_io_out_w_bits_last;
  assign axi4XBar_io_in_1_b_ready = axiBridge_1_io_out_b_ready;
  assign axi4XBar_io_in_1_ar_valid = axiBridge_1_io_out_ar_valid;
  assign axi4XBar_io_in_1_ar_bits_addr = axiBridge_1_io_out_ar_bits_addr;
  assign axi4XBar_io_in_1_ar_bits_size = axiBridge_1_io_out_ar_bits_size;
  assign axi4XBar_io_in_1_r_ready = axiBridge_1_io_out_r_ready;
  assign axi4XBar_io_in_2_aw_valid = axi4XBar_io_in_2_toAXIbridge_io_out_aw_valid;
  assign axi4XBar_io_in_2_aw_bits_addr = axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_addr;
  assign axi4XBar_io_in_2_aw_bits_id = axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_id;
  assign axi4XBar_io_in_2_aw_bits_len = axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_len;
  assign axi4XBar_io_in_2_aw_bits_size = axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_size;
  assign axi4XBar_io_in_2_aw_bits_burst = axi4XBar_io_in_2_toAXIbridge_io_out_aw_bits_burst;
  assign axi4XBar_io_in_2_w_valid = axi4XBar_io_in_2_toAXIbridge_io_out_w_valid;
  assign axi4XBar_io_in_2_w_bits_strb = axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_strb;
  assign axi4XBar_io_in_2_w_bits_data = axi4XBar_io_in_2_toAXIbridge_io_out_w_bits_data;
  assign axi4XBar_io_in_2_b_ready = axi4XBar_io_in_2_toAXIbridge_io_out_b_ready;
  assign axi4XBar_io_in_2_ar_valid = axi4XBar_io_in_2_toAXIbridge_io_out_ar_valid;
  assign axi4XBar_io_in_2_ar_bits_addr = axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_addr;
  assign axi4XBar_io_in_2_ar_bits_size = axi4XBar_io_in_2_toAXIbridge_io_out_ar_bits_size;
  assign axi4XBar_io_in_2_r_ready = axi4XBar_io_in_2_toAXIbridge_io_out_r_ready;
  assign axi4XBar_io_in_3_aw_valid = axi4XBar_io_in_3_toAXIbridge_io_out_aw_valid;
  assign axi4XBar_io_in_3_aw_bits_addr = axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_addr;
  assign axi4XBar_io_in_3_aw_bits_id = axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_id;
  assign axi4XBar_io_in_3_aw_bits_len = axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_len;
  assign axi4XBar_io_in_3_aw_bits_size = axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_size;
  assign axi4XBar_io_in_3_aw_bits_burst = axi4XBar_io_in_3_toAXIbridge_io_out_aw_bits_burst;
  assign axi4XBar_io_in_3_w_valid = axi4XBar_io_in_3_toAXIbridge_io_out_w_valid;
  assign axi4XBar_io_in_3_w_bits_strb = axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_strb;
  assign axi4XBar_io_in_3_w_bits_data = axi4XBar_io_in_3_toAXIbridge_io_out_w_bits_data;
  assign axi4XBar_io_in_3_b_ready = axi4XBar_io_in_3_toAXIbridge_io_out_b_ready;
  assign axi4XBar_io_in_3_ar_valid = axi4XBar_io_in_3_toAXIbridge_io_out_ar_valid;
  assign axi4XBar_io_in_3_ar_bits_addr = axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_addr;
  assign axi4XBar_io_in_3_ar_bits_size = axi4XBar_io_in_3_toAXIbridge_io_out_ar_bits_size;
  assign axi4XBar_io_in_3_r_ready = axi4XBar_io_in_3_toAXIbridge_io_out_r_ready;
  assign axi4XBar_io_in_4_aw_valid = axi4XBar_io_in_4_toAXIbridge_io_out_aw_valid;
  assign axi4XBar_io_in_4_aw_bits_addr = axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_addr;
  assign axi4XBar_io_in_4_aw_bits_id = axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_id;
  assign axi4XBar_io_in_4_aw_bits_len = axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_len;
  assign axi4XBar_io_in_4_aw_bits_size = axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_size;
  assign axi4XBar_io_in_4_aw_bits_burst = axi4XBar_io_in_4_toAXIbridge_io_out_aw_bits_burst;
  assign axi4XBar_io_in_4_w_valid = axi4XBar_io_in_4_toAXIbridge_io_out_w_valid;
  assign axi4XBar_io_in_4_w_bits_strb = axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_strb;
  assign axi4XBar_io_in_4_w_bits_data = axi4XBar_io_in_4_toAXIbridge_io_out_w_bits_data;
  assign axi4XBar_io_in_4_b_ready = axi4XBar_io_in_4_toAXIbridge_io_out_b_ready;
  assign axi4XBar_io_in_4_ar_valid = axi4XBar_io_in_4_toAXIbridge_io_out_ar_valid;
  assign axi4XBar_io_in_4_ar_bits_addr = axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_addr;
  assign axi4XBar_io_in_4_ar_bits_size = axi4XBar_io_in_4_toAXIbridge_io_out_ar_bits_size;
  assign axi4XBar_io_in_4_r_ready = axi4XBar_io_in_4_toAXIbridge_io_out_r_ready;
  assign axi4XBar_io_in_5_aw_valid = axi4XBar_io_in_5_toAXIbridge_io_out_aw_valid;
  assign axi4XBar_io_in_5_aw_bits_addr = axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_addr;
  assign axi4XBar_io_in_5_aw_bits_id = axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_id;
  assign axi4XBar_io_in_5_aw_bits_len = axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_len;
  assign axi4XBar_io_in_5_aw_bits_size = axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_size;
  assign axi4XBar_io_in_5_aw_bits_burst = axi4XBar_io_in_5_toAXIbridge_io_out_aw_bits_burst;
  assign axi4XBar_io_in_5_w_valid = axi4XBar_io_in_5_toAXIbridge_io_out_w_valid;
  assign axi4XBar_io_in_5_w_bits_strb = axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_strb;
  assign axi4XBar_io_in_5_w_bits_data = axi4XBar_io_in_5_toAXIbridge_io_out_w_bits_data;
  assign axi4XBar_io_in_5_b_ready = axi4XBar_io_in_5_toAXIbridge_io_out_b_ready;
  assign axi4XBar_io_in_5_ar_valid = axi4XBar_io_in_5_toAXIbridge_io_out_ar_valid;
  assign axi4XBar_io_in_5_ar_bits_addr = axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_addr;
  assign axi4XBar_io_in_5_ar_bits_size = axi4XBar_io_in_5_toAXIbridge_io_out_ar_bits_size;
  assign axi4XBar_io_in_5_r_ready = axi4XBar_io_in_5_toAXIbridge_io_out_r_ready;
  assign axi4XBar_io_out_aw_ready = io_master_awready;
  assign axi4XBar_io_out_w_ready = io_master_wready;
  assign axi4XBar_io_out_b_valid = io_master_bvalid;
  assign axi4XBar_io_out_ar_ready = io_master_arready;
  assign axi4XBar_io_out_r_valid = io_master_rvalid;
  assign axi4XBar_io_out_r_bits_data = io_master_rdata;
  assign axi4XBar_io_out_r_bits_last = io_master_rlast;
  assign mmioXBar_clock = clock;
  assign mmioXBar_reset = reset;
  assign mmioXBar_io_in_req_valid = overlay_io_dmmio_req_valid;
  assign mmioXBar_io_in_req_bits_addr = overlay_io_dmmio_req_bits_addr;
  assign mmioXBar_io_in_req_bits_wdata = overlay_io_dmmio_req_bits_wdata;
  assign mmioXBar_io_in_req_bits_size = overlay_io_dmmio_req_bits_size;
  assign mmioXBar_io_in_req_bits_cmd = overlay_io_dmmio_req_bits_cmd;
  assign mmioXBar_io_out_0_req_ready = axi4XBar_io_in_3_toAXIbridge_io_in_req_ready;
  assign mmioXBar_io_out_0_resp_valid = axi4XBar_io_in_3_toAXIbridge_io_in_resp_valid;
  assign mmioXBar_io_out_0_resp_bits_rdata = axi4XBar_io_in_3_toAXIbridge_io_in_resp_bits_rdata;
  assign mmioXBar_io_out_1_req_ready = clint_io_in_toAXIbridge_io_in_req_ready;
  assign mmioXBar_io_out_1_resp_valid = clint_io_in_toAXIbridge_io_in_resp_valid;
  assign mmioXBar_io_out_1_resp_bits_rdata = clint_io_in_toAXIbridge_io_in_resp_bits_rdata;
  assign mmioXBar_io_out_2_req_ready = axi4XBar_io_in_4_toAXIbridge_io_in_req_ready;
  assign mmioXBar_io_out_2_resp_valid = axi4XBar_io_in_4_toAXIbridge_io_in_resp_valid;
  assign mmioXBar_io_out_2_resp_bits_rdata = axi4XBar_io_in_4_toAXIbridge_io_in_resp_bits_rdata;
  assign mmioXBar_io_out_3_req_ready = axi4XBar_io_in_5_toAXIbridge_io_in_req_ready;
  assign mmioXBar_io_out_3_resp_valid = axi4XBar_io_in_5_toAXIbridge_io_in_resp_valid;
  assign mmioXBar_io_out_3_resp_bits_rdata = axi4XBar_io_in_5_toAXIbridge_io_in_resp_bits_rdata;
  assign axiBridge_0_clock = clock;
  assign axiBridge_0_reset = reset;
  assign axiBridge_0_io_in_req_valid = xConnect_io_out_mem_req_valid;
  assign axiBridge_0_io_in_req_bits_addr = xConnect_io_out_mem_req_bits_addr;
  assign axiBridge_0_io_in_req_bits_wdata = xConnect_io_out_mem_req_bits_wdata;
  assign axiBridge_0_io_in_req_bits_cmd = xConnect_io_out_mem_req_bits_cmd;
  assign axiBridge_0_io_out_aw_ready = axi4XBar_io_in_0_aw_ready;
  assign axiBridge_0_io_out_w_ready = axi4XBar_io_in_0_w_ready;
  assign axiBridge_0_io_out_b_valid = axi4XBar_io_in_0_b_valid;
  assign axiBridge_0_io_out_ar_ready = axi4XBar_io_in_0_ar_ready;
  assign axiBridge_0_io_out_r_valid = axi4XBar_io_in_0_r_valid;
  assign axiBridge_0_io_out_r_bits_data = axi4XBar_io_in_0_r_bits_data;
  assign axiBridge_0_io_out_r_bits_last = axi4XBar_io_in_0_r_bits_last;
  assign axiBridge_1_clock = clock;
  assign axiBridge_1_reset = reset;
  assign axiBridge_1_io_in_req_valid = overlay_io_dmem_req_valid;
  assign axiBridge_1_io_in_req_bits_addr = overlay_io_dmem_req_bits_addr;
  assign axiBridge_1_io_in_req_bits_wdata = overlay_io_dmem_req_bits_wdata;
  assign axiBridge_1_io_in_req_bits_cmd = overlay_io_dmem_req_bits_cmd;
  assign axiBridge_1_io_out_aw_ready = axi4XBar_io_in_1_aw_ready;
  assign axiBridge_1_io_out_w_ready = axi4XBar_io_in_1_w_ready;
  assign axiBridge_1_io_out_b_valid = axi4XBar_io_in_1_b_valid;
  assign axiBridge_1_io_out_ar_ready = axi4XBar_io_in_1_ar_ready;
  assign axiBridge_1_io_out_r_valid = axi4XBar_io_in_1_r_valid;
  assign axiBridge_1_io_out_r_bits_data = axi4XBar_io_in_1_r_bits_data;
  assign axiBridge_1_io_out_r_bits_last = axi4XBar_io_in_1_r_bits_last;
  assign clint_io_in_toAXIbridge_clock = clock;
  assign clint_io_in_toAXIbridge_reset = reset;
  assign clint_io_in_toAXIbridge_io_in_req_valid = mmioXBar_io_out_1_req_valid;
  assign clint_io_in_toAXIbridge_io_in_req_bits_addr = mmioXBar_io_out_1_req_bits_addr;
  assign clint_io_in_toAXIbridge_io_in_req_bits_wdata = mmioXBar_io_out_1_req_bits_wdata;
  assign clint_io_in_toAXIbridge_io_in_req_bits_size = mmioXBar_io_out_1_req_bits_size;
  assign clint_io_in_toAXIbridge_io_in_req_bits_cmd = mmioXBar_io_out_1_req_bits_cmd;
  assign clint_io_in_toAXIbridge_io_in_resp_ready = mmioXBar_io_out_1_resp_ready;
  assign clint_io_in_toAXIbridge_io_out_aw_ready = clint_io_in_aw_ready;
  assign clint_io_in_toAXIbridge_io_out_w_ready = clint_io_in_w_ready;
  assign clint_io_in_toAXIbridge_io_out_b_valid = clint_io_in_b_valid;
  assign clint_io_in_toAXIbridge_io_out_ar_ready = clint_io_in_ar_ready;
  assign clint_io_in_toAXIbridge_io_out_r_valid = clint_io_in_r_valid;
  assign clint_io_in_toAXIbridge_io_out_r_bits_data = clint_io_in_r_bits_data;
  assign axi4XBar_io_in_2_toAXIbridge_clock = clock;
  assign axi4XBar_io_in_2_toAXIbridge_reset = reset;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_req_valid = overlay_io_immio_req_valid;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_addr = overlay_io_immio_req_bits_addr;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_wdata = 64'h0;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_size = overlay_io_immio_req_bits_size;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_req_bits_cmd = 3'h0;
  assign axi4XBar_io_in_2_toAXIbridge_io_in_resp_ready = 1'h1;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_aw_ready = axi4XBar_io_in_2_aw_ready;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_w_ready = axi4XBar_io_in_2_w_ready;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_b_valid = axi4XBar_io_in_2_b_valid;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_ar_ready = axi4XBar_io_in_2_ar_ready;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_r_valid = axi4XBar_io_in_2_r_valid;
  assign axi4XBar_io_in_2_toAXIbridge_io_out_r_bits_data = axi4XBar_io_in_2_r_bits_data;
  assign axi4XBar_io_in_3_toAXIbridge_clock = clock;
  assign axi4XBar_io_in_3_toAXIbridge_reset = reset;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_req_valid = mmioXBar_io_out_0_req_valid;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_addr = mmioXBar_io_out_0_req_bits_addr;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_wdata = mmioXBar_io_out_0_req_bits_wdata;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_size = mmioXBar_io_out_0_req_bits_size;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_req_bits_cmd = mmioXBar_io_out_0_req_bits_cmd;
  assign axi4XBar_io_in_3_toAXIbridge_io_in_resp_ready = mmioXBar_io_out_0_resp_ready;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_aw_ready = axi4XBar_io_in_3_aw_ready;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_w_ready = axi4XBar_io_in_3_w_ready;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_b_valid = axi4XBar_io_in_3_b_valid;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_ar_ready = axi4XBar_io_in_3_ar_ready;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_r_valid = axi4XBar_io_in_3_r_valid;
  assign axi4XBar_io_in_3_toAXIbridge_io_out_r_bits_data = axi4XBar_io_in_3_r_bits_data;
  assign axi4XBar_io_in_4_toAXIbridge_clock = clock;
  assign axi4XBar_io_in_4_toAXIbridge_reset = reset;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_req_valid = mmioXBar_io_out_2_req_valid;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_addr = mmioXBar_io_out_2_req_bits_addr;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_wdata = mmioXBar_io_out_2_req_bits_wdata;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_size = mmioXBar_io_out_2_req_bits_size;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_req_bits_cmd = mmioXBar_io_out_2_req_bits_cmd;
  assign axi4XBar_io_in_4_toAXIbridge_io_in_resp_ready = mmioXBar_io_out_2_resp_ready;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_aw_ready = axi4XBar_io_in_4_aw_ready;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_w_ready = axi4XBar_io_in_4_w_ready;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_b_valid = axi4XBar_io_in_4_b_valid;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_ar_ready = axi4XBar_io_in_4_ar_ready;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_r_valid = axi4XBar_io_in_4_r_valid;
  assign axi4XBar_io_in_4_toAXIbridge_io_out_r_bits_data = axi4XBar_io_in_4_r_bits_data;
  assign axi4XBar_io_in_5_toAXIbridge_clock = clock;
  assign axi4XBar_io_in_5_toAXIbridge_reset = reset;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_req_valid = mmioXBar_io_out_3_req_valid;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_addr = mmioXBar_io_out_3_req_bits_addr;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_wdata = mmioXBar_io_out_3_req_bits_wdata;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_size = mmioXBar_io_out_3_req_bits_size;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_req_bits_cmd = mmioXBar_io_out_3_req_bits_cmd;
  assign axi4XBar_io_in_5_toAXIbridge_io_in_resp_ready = mmioXBar_io_out_3_resp_ready;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_aw_ready = axi4XBar_io_in_5_aw_ready;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_w_ready = axi4XBar_io_in_5_w_ready;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_b_valid = axi4XBar_io_in_5_b_valid;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_ar_ready = axi4XBar_io_in_5_ar_ready;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_r_valid = axi4XBar_io_in_5_r_valid;
  assign axi4XBar_io_in_5_toAXIbridge_io_out_r_bits_data = axi4XBar_io_in_5_r_bits_data;
endmodule
