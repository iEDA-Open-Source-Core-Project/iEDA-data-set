module ysyx_22040886_alu(
  input  [15:0] io_ctrl,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_result,
  output        io_overflow,
  input         io_data_w
);
  wire [5:0] sa = io_in2[5:0]; // @[alu.scala 23:28]
  wire [4:0] sa_for_32bit = io_in2[4:0]; // @[alu.scala 24:30]
  wire [63:0] answer_and = io_in1 & io_in2; // @[alu.scala 26:32]
  wire [63:0] answer_or = io_in1 | io_in2; // @[alu.scala 27:32]
  wire [63:0] answer_xor = io_in1 ^ io_in2; // @[alu.scala 28:32]
  wire [63:0] answer_nor = ~answer_or; // @[alu.scala 29:25]
  wire  answer_slt = $signed(io_in1) < $signed(io_in2); // @[alu.scala 31:43]
  wire  answer_sltu = io_in1 < io_in2; // @[alu.scala 32:36]
  wire [126:0] _GEN_20 = {{63'd0}, io_in1}; // @[alu.scala 33:31]
  wire [126:0] answer_sll = _GEN_20 << sa; // @[alu.scala 33:31]
  wire [63:0] answer_srl = io_in1 >> sa; // @[alu.scala 35:31]
  wire [31:0] answer_srlw = io_in1[31:0] >> sa_for_32bit; // @[alu.scala 36:37]
  wire [63:0] answer_sra = $signed(io_in1) >>> sa; // @[alu.scala 37:46]
  wire [31:0] _answer_sraw_T_1 = io_in1[31:0]; // @[alu.scala 38:38]
  wire [31:0] answer_sraw = $signed(_answer_sraw_T_1) >>> sa_for_32bit; // @[alu.scala 38:62]
  wire [31:0] _answer_lui_T_1 = {io_in2[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [7:0] answer_lui_lo_lo = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] answer_lui_lo = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],answer_lui_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _answer_lui_T_34 = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],answer_lui_lo_lo,answer_lui_lo}; // @[Cat.scala 31:58]
  wire [63:0] answer_lui = {_answer_lui_T_34,io_in2[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [64:0] in1_extend = {io_in1[63],io_in1}; // @[Cat.scala 31:58]
  wire [64:0] in2_extend = {io_in2[63],io_in2}; // @[Cat.scala 31:58]
  wire [64:0] answer_add = in1_extend + in2_extend; // @[alu.scala 45:35]
  wire [64:0] answer_sub = in1_extend - in2_extend; // @[alu.scala 46:35]
  wire [15:0] _normal_result_T = {{1'd0}, io_ctrl[15:1]}; // @[alu.scala 49:16]
  wire [15:0] _normal_result_T_3 = {{2'd0}, io_ctrl[15:2]}; // @[alu.scala 50:16]
  wire [15:0] _normal_result_T_6 = {{3'd0}, io_ctrl[15:3]}; // @[alu.scala 51:16]
  wire [15:0] _normal_result_T_9 = {{6'd0}, io_ctrl[15:6]}; // @[alu.scala 52:16]
  wire [15:0] _normal_result_T_12 = {{8'd0}, io_ctrl[15:8]}; // @[alu.scala 53:16]
  wire [15:0] _normal_result_T_15 = {{9'd0}, io_ctrl[15:9]}; // @[alu.scala 54:16]
  wire [15:0] _normal_result_T_18 = {{4'd0}, io_ctrl[15:4]}; // @[alu.scala 55:16]
  wire [15:0] _normal_result_T_20 = {{11'd0}, io_ctrl[15:11]}; // @[alu.scala 56:16]
  wire [15:0] _normal_result_T_22 = {{10'd0}, io_ctrl[15:10]}; // @[alu.scala 57:16]
  wire [15:0] _normal_result_T_26 = {{7'd0}, io_ctrl[15:7]}; // @[alu.scala 59:16]
  wire [15:0] _normal_result_T_28 = {{12'd0}, io_ctrl[15:12]}; // @[alu.scala 60:16]
  wire [15:0] _normal_result_T_30 = {{13'd0}, io_ctrl[15:13]}; // @[alu.scala 61:16]
  wire [15:0] _normal_result_T_32 = {{15'd0}, io_ctrl[15]}; // @[alu.scala 62:16]
  wire [63:0] _normal_result_T_34 = io_data_w ? {{32'd0}, answer_sraw} : answer_sra; // @[alu.scala 62:35]
  wire [15:0] _normal_result_T_35 = {{5'd0}, io_ctrl[15:5]}; // @[alu.scala 63:16]
  wire [63:0] _normal_result_T_37 = io_data_w ? {{32'd0}, answer_srlw} : answer_srl; // @[alu.scala 63:35]
  wire [15:0] _normal_result_T_38 = {{14'd0}, io_ctrl[15:14]}; // @[alu.scala 64:16]
  wire [63:0] _normal_result_T_40 = _normal_result_T[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_41 = _normal_result_T_3[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_42 = _normal_result_T_6[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_43 = _normal_result_T_9[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_44 = _normal_result_T_12[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_45 = _normal_result_T_15[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_46 = _normal_result_T_18[0] ? answer_and : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_47 = _normal_result_T_20[0] ? answer_or : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_48 = _normal_result_T_22[0] ? answer_nor : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_49 = io_ctrl[0] ? answer_xor : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_50 = _normal_result_T_26[0] ? answer_lui : 64'h0; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_51 = _normal_result_T_28[0] ? answer_sll : 127'h0; // @[Mux.scala 27:73]
  wire  _normal_result_T_52 = _normal_result_T_30[0] & answer_slt; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_53 = _normal_result_T_32[0] ? _normal_result_T_34 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_54 = _normal_result_T_35[0] ? _normal_result_T_37 : 64'h0; // @[Mux.scala 27:73]
  wire  _normal_result_T_55 = _normal_result_T_38[0] & answer_sltu; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_56 = _normal_result_T_40 | _normal_result_T_41; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_57 = _normal_result_T_56 | _normal_result_T_42; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_58 = _normal_result_T_57 | _normal_result_T_43; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_59 = _normal_result_T_58 | _normal_result_T_44; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_60 = _normal_result_T_59 | _normal_result_T_45; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_61 = _normal_result_T_60 | _normal_result_T_46; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_62 = _normal_result_T_61 | _normal_result_T_47; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_63 = _normal_result_T_62 | _normal_result_T_48; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_64 = _normal_result_T_63 | _normal_result_T_49; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_65 = _normal_result_T_64 | _normal_result_T_50; // @[Mux.scala 27:73]
  wire [126:0] _GEN_15 = {{63'd0}, _normal_result_T_65}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_66 = _GEN_15 | _normal_result_T_51; // @[Mux.scala 27:73]
  wire [126:0] _GEN_16 = {{126'd0}, _normal_result_T_52}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_67 = _normal_result_T_66 | _GEN_16; // @[Mux.scala 27:73]
  wire [126:0] _GEN_17 = {{63'd0}, _normal_result_T_53}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_68 = _normal_result_T_67 | _GEN_17; // @[Mux.scala 27:73]
  wire [126:0] _GEN_18 = {{63'd0}, _normal_result_T_54}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_69 = _normal_result_T_68 | _GEN_18; // @[Mux.scala 27:73]
  wire [126:0] _GEN_19 = {{126'd0}, _normal_result_T_55}; // @[Mux.scala 27:73]
  wire [126:0] normal_result = _normal_result_T_69 | _GEN_19; // @[Mux.scala 27:73]
  wire [7:0] io_result_lo_lo = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[31
    ],normal_result[31],normal_result[31],normal_result[31]}; // @[Cat.scala 31:58]
  wire [15:0] io_result_lo = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[31],
    normal_result[31],normal_result[31],normal_result[31],io_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _io_result_T_33 = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[
    31],normal_result[31],normal_result[31],normal_result[31],io_result_lo_lo,io_result_lo}; // @[Cat.scala 31:58]
  wire [63:0] _io_result_T_35 = {_io_result_T_33,normal_result[31:0]}; // @[Cat.scala 31:58]
  wire [126:0] _io_result_T_36 = io_data_w ? {{63'd0}, _io_result_T_35} : normal_result; // @[alu.scala 67:21]
  assign io_result = _io_result_T_36[63:0]; // @[alu.scala 67:15]
  assign io_overflow = _normal_result_T_3[0] & answer_add[64] != answer_add[63] | _normal_result_T_12[0] & answer_sub[64
    ] != answer_sub[63]; // @[alu.scala 68:101]
endmodule
module ysyx_22040886_br(
  input         reset,
  input  [63:0] io_r1,
  input  [63:0] io_r2,
  input  [5:0]  io_branch,
  output        io_exe
);
  wire  _result_T = io_r1 >= io_r2; // @[br.scala 24:38]
  wire  _result_T_1 = io_r1 < io_r2; // @[br.scala 25:37]
  wire  _result_T_4 = $signed(io_r1) >= $signed(io_r2); // @[br.scala 26:37]
  wire  _result_T_7 = $signed(io_r1) < $signed(io_r2); // @[br.scala 27:37]
  wire  _result_T_8 = io_r1 != io_r2; // @[br.scala 28:30]
  wire  _result_T_9 = io_r1 == io_r2; // @[br.scala 29:30]
  wire [5:0] result = {_result_T,_result_T_1,_result_T_4,_result_T_7,_result_T_8,_result_T_9}; // @[Cat.scala 31:58]
  wire [5:0] _io_exe_T_4 = result & io_branch; // @[br.scala 30:57]
  assign io_exe = ~reset & _io_exe_T_4 != 6'h0; // @[br.scala 30:45]
endmodule
module ysyx_22040886_cfu(
  input         reset,
  input         io_Inst_Fifo_Empty,
  input         io_dmem_calD,
  input         io_BranchD_Flag,
  input         io_JRD,
  input         io_CanBranchD,
  input         io_DivPendingE,
  input         io_DataPendingM,
  input         io_InException,
  input  [4:0]  io_WriteRegE,
  input         io_RegWriteE,
  input         io_csrToRegE,
  input  [4:0]  io_WriteRegM,
  input         io_MemToRegM,
  input         io_RegWriteM,
  input         io_csrWriteM,
  input  [4:0]  io_WriteRegM2,
  input         io_MemToRegM2,
  input         io_RegWriteM2,
  input         io_csrWriteM2,
  input  [4:0]  io_WriteRegW,
  input         io_RegWriteW,
  input  [11:0] io_ReadcsrAddrE,
  input  [11:0] io_WritecsrAddrM,
  input  [11:0] io_WritecsrAddrM2,
  input  [4:0]  io_R2D,
  input  [4:0]  io_R1D,
  input  [4:0]  io_R2E,
  input  [4:0]  io_R1E,
  output        io_StallF,
  output        io_StallD,
  output        io_StallE,
  output        io_StallM,
  output        io_StallM2,
  output        io_StallW,
  output        io_FlushD,
  output        io_FlushE,
  output        io_FlushM,
  output        io_FlushM2,
  output        io_FlushW,
  output [1:0]  io_Forward1E,
  output [1:0]  io_Forward2E,
  output [1:0]  io_Forward1D,
  output [1:0]  io_Forward2D,
  output [1:0]  io_ForwardcsrE
);
  wire  _io_Forward2D_T_3 = io_R2D == io_WriteRegM & io_RegWriteM; // @[cfu.scala 94:73]
  wire  _io_Forward2D_T_5 = ~io_MemToRegM; // @[cfu.scala 94:99]
  wire  _io_Forward2D_T_9 = io_R2D == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 95:34]
  wire  _io_Forward2D_T_11 = ~io_MemToRegM2; // @[cfu.scala 95:61]
  wire  _io_Forward2D_T_12 = io_R2D == io_WriteRegM2 & io_RegWriteM2 & ~io_MemToRegM2; // @[cfu.scala 95:58]
  wire [1:0] _io_Forward2D_T_13 = _io_Forward2D_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 94:131]
  wire [1:0] _io_Forward2D_T_14 = io_R2D == io_WriteRegM & io_RegWriteM & ~io_MemToRegM ? 2'h1 : _io_Forward2D_T_13; // @[cfu.scala 94:48]
  wire  _io_Forward1D_T_3 = io_R1D == io_WriteRegM & io_RegWriteM; // @[cfu.scala 96:73]
  wire  _io_Forward1D_T_9 = io_R1D == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 97:34]
  wire  _io_Forward1D_T_12 = io_R1D == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 97:58]
  wire [1:0] _io_Forward1D_T_13 = _io_Forward1D_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 96:131]
  wire [1:0] _io_Forward1D_T_14 = io_R1D == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5 ? 2'h1 : _io_Forward1D_T_13; // @[cfu.scala 96:48]
  wire  _io_Forward2E_T_3 = io_R2E == io_WriteRegM & io_RegWriteM; // @[cfu.scala 103:34]
  wire  _io_Forward2E_T_6 = io_R2E == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5; // @[cfu.scala 103:57]
  wire  _io_Forward2E_T_9 = io_R2E == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 104:35]
  wire  _io_Forward2E_T_12 = io_R2E == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 104:59]
  wire  _io_Forward2E_T_15 = io_R2E == io_WriteRegW & io_RegWriteW; // @[cfu.scala 105:34]
  wire [1:0] _io_Forward2E_T_17 = _io_Forward2E_T_12 ? 2'h3 : {{1'd0}, _io_Forward2E_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_Forward2E_T_18 = _io_Forward2E_T_6 ? 2'h2 : _io_Forward2E_T_17; // @[Mux.scala 101:16]
  wire  _io_Forward1E_T_3 = io_R1E == io_WriteRegM & io_RegWriteM; // @[cfu.scala 110:34]
  wire  _io_Forward1E_T_6 = io_R1E == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5; // @[cfu.scala 110:57]
  wire  _io_Forward1E_T_9 = io_R1E == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 111:35]
  wire  _io_Forward1E_T_12 = io_R1E == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 111:59]
  wire  _io_Forward1E_T_15 = io_R1E == io_WriteRegW & io_RegWriteW; // @[cfu.scala 112:34]
  wire [1:0] _io_Forward1E_T_17 = _io_Forward1E_T_12 ? 2'h3 : {{1'd0}, _io_Forward1E_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_Forward1E_T_18 = _io_Forward1E_T_6 ? 2'h2 : _io_Forward1E_T_17; // @[Mux.scala 101:16]
  wire  _io_ForwardcsrE_T_3 = io_ReadcsrAddrE == io_WritecsrAddrM & io_csrWriteM; // @[cfu.scala 118:59]
  wire  _io_ForwardcsrE_T_6 = io_ReadcsrAddrE == io_WritecsrAddrM2 & io_csrWriteM2; // @[cfu.scala 119:60]
  wire [1:0] _io_ForwardcsrE_T_7 = _io_ForwardcsrE_T_6 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardcsrE_T_8 = _io_ForwardcsrE_T_3 ? 2'h1 : _io_ForwardcsrE_T_7; // @[Mux.scala 101:16]
  wire  _br_Stall_T_5 = io_WriteRegE == io_R1D; // @[cfu.scala 125:75]
  wire  _br_Stall_T_10 = io_WriteRegM == io_R1D; // @[cfu.scala 126:74]
  wire  _br_Stall_T_12 = io_MemToRegM & (io_WriteRegM == io_R2D | io_WriteRegM == io_R1D); // @[cfu.scala 126:30]
  wire  _br_Stall_T_13 = io_RegWriteE & (io_WriteRegE == io_R2D | io_WriteRegE == io_R1D) | _br_Stall_T_12; // @[cfu.scala 125:88]
  wire  _br_Stall_T_16 = io_WriteRegM2 == io_R1D; // @[cfu.scala 127:77]
  wire  _br_Stall_T_18 = io_MemToRegM2 & (io_WriteRegM2 == io_R2D | io_WriteRegM2 == io_R1D); // @[cfu.scala 127:31]
  wire  _br_Stall_T_19 = _br_Stall_T_13 | _br_Stall_T_18; // @[cfu.scala 126:87]
  wire  _br_Stall_T_20 = io_CanBranchD & io_BranchD_Flag & _br_Stall_T_19; // @[cfu.scala 124:71]
  wire  _br_Stall_T_22 = ~io_InException; // @[cfu.scala 127:95]
  wire  br_Stall = _br_Stall_T_20 & ~io_InException; // @[cfu.scala 127:92]
  wire  _jr_Stall_T_8 = io_MemToRegM & _br_Stall_T_10; // @[cfu.scala 130:30]
  wire  _jr_Stall_T_9 = io_RegWriteE & _br_Stall_T_5 | _jr_Stall_T_8; // @[cfu.scala 129:61]
  wire  _jr_Stall_T_12 = io_MemToRegM2 & _br_Stall_T_16; // @[cfu.scala 131:31]
  wire  _jr_Stall_T_13 = _jr_Stall_T_9 | _jr_Stall_T_12; // @[cfu.scala 130:62]
  wire  _jr_Stall_T_14 = (io_JRD | io_dmem_calD) & _jr_Stall_T_13; // @[cfu.scala 128:60]
  wire  dmem_addr_cal_Stall = _jr_Stall_T_14 & _br_Stall_T_22; // @[cfu.scala 131:65]
  wire  _mem2regM_Stall_T_9 = _io_Forward1E_T_3 & io_MemToRegM; // @[cfu.scala 142:87]
  wire  _mem2regM_Stall_T_10 = _io_Forward2E_T_3 & io_MemToRegM | _mem2regM_Stall_T_9; // @[cfu.scala 141:120]
  wire  _mem2regM_Stall_T_15 = _io_Forward2D_T_3 & io_MemToRegM; // @[cfu.scala 143:87]
  wire  _mem2regM_Stall_T_16 = _mem2regM_Stall_T_10 | _mem2regM_Stall_T_15; // @[cfu.scala 142:111]
  wire  _mem2regM_Stall_T_21 = _io_Forward1D_T_3 & io_MemToRegM; // @[cfu.scala 144:87]
  wire  _mem2regM_Stall_T_22 = _mem2regM_Stall_T_16 | _mem2regM_Stall_T_21; // @[cfu.scala 143:111]
  wire  _mem2regM_Stall_T_27 = _io_Forward2E_T_9 & io_MemToRegM2; // @[cfu.scala 145:89]
  wire  _mem2regM_Stall_T_28 = _mem2regM_Stall_T_22 | _mem2regM_Stall_T_27; // @[cfu.scala 144:111]
  wire  _mem2regM_Stall_T_33 = _io_Forward1E_T_9 & io_MemToRegM2; // @[cfu.scala 146:89]
  wire  _mem2regM_Stall_T_34 = _mem2regM_Stall_T_28 | _mem2regM_Stall_T_33; // @[cfu.scala 145:114]
  wire  _mem2regM_Stall_T_39 = _io_Forward2D_T_9 & io_MemToRegM2; // @[cfu.scala 147:89]
  wire  _mem2regM_Stall_T_40 = _mem2regM_Stall_T_34 | _mem2regM_Stall_T_39; // @[cfu.scala 146:114]
  wire  _mem2regM_Stall_T_45 = _io_Forward1D_T_9 & io_MemToRegM2; // @[cfu.scala 148:89]
  wire  mem2regM_Stall = _mem2regM_Stall_T_40 | _mem2regM_Stall_T_45; // @[cfu.scala 147:114]
  wire  _has_Stall_T = br_Stall | dmem_addr_cal_Stall; // @[cfu.scala 155:44]
  wire  _io_StallF_T_5 = _has_Stall_T | io_DivPendingE | io_DataPendingM | mem2regM_Stall; // @[cfu.scala 160:133]
  wire  _io_StallM_T_1 = ~io_DataPendingM; // @[cfu.scala 163:39]
  assign io_StallF = reset | ~(_has_Stall_T | io_DivPendingE | io_DataPendingM | mem2regM_Stall | io_Inst_Fifo_Empty); // @[cfu.scala 160:21]
  assign io_StallD = reset | ~_io_StallF_T_5; // @[cfu.scala 161:21]
  assign io_StallE = reset | ~(io_DivPendingE | io_DataPendingM | mem2regM_Stall); // @[cfu.scala 162:21]
  assign io_StallM = reset | ~io_DataPendingM; // @[cfu.scala 163:21]
  assign io_StallM2 = reset | _io_StallM_T_1; // @[cfu.scala 164:22]
  assign io_StallW = reset | _io_StallM_T_1; // @[cfu.scala 165:21]
  assign io_FlushD = reset ? 1'h0 : io_InException; // @[cfu.scala 167:21]
  assign io_FlushE = reset ? 1'h0 : io_StallE & _has_Stall_T | io_InException; // @[cfu.scala 168:21]
  assign io_FlushM = reset ? 1'h0 : io_StallM & (io_DivPendingE | mem2regM_Stall) | io_InException; // @[cfu.scala 169:21]
  assign io_FlushM2 = reset ? 1'h0 : io_InException; // @[cfu.scala 170:22]
  assign io_FlushW = reset ? 1'h0 : io_StallW & (io_DataPendingM | io_InException); // @[cfu.scala 171:21]
  assign io_Forward1E = io_R1E == 5'h0 ? 2'h0 : _io_Forward1E_T_18; // @[cfu.scala 109:24]
  assign io_Forward2E = io_R2E == 5'h0 ? 2'h0 : _io_Forward2E_T_18; // @[cfu.scala 102:24]
  assign io_Forward1D = io_R1D == 5'h0 ? 2'h0 : _io_Forward1D_T_14; // @[cfu.scala 96:24]
  assign io_Forward2D = io_R2D == 5'h0 ? 2'h0 : _io_Forward2D_T_14; // @[cfu.scala 94:24]
  assign io_ForwardcsrE = io_csrToRegE ? _io_ForwardcsrE_T_8 : 2'h0; // @[cfu.scala 117:26]
endmodule
module ysyx_22040886_csr(
  input         clock,
  input         reset,
  input  [11:0] io_csr_read_addr,
  input  [11:0] io_csr_write_addr,
  input  [63:0] io_csr_write_data,
  input         io_csr_write_en,
  input  [63:0] io_pc,
  input  [30:0] io_exception_type_i,
  output [63:0] io_return_pc,
  output        io_exception,
  output [63:0] io_csr_read_data,
  output        io_icache_tags_flush,
  input         io_int_type_timer,
  input         io_int_type_out_int,
  input  [63:0] io_stageW_pc,
  output        io_Int_able,
  output        io_int_type_able_timer,
  output        io_int_type_able_out_int
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] csr_cause; // @[csr.scala 61:28]
  reg [63:0] csr_status; // @[csr.scala 62:25]
  wire  _csr_status_to_be_T_3 = io_csr_write_en & io_csr_write_addr == 12'h300; // @[csr.scala 183:33]
  wire  csr_status_to_vec_63 = csr_status[63]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_62 = csr_status[62]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_61 = csr_status[61]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_60 = csr_status[60]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_59 = csr_status[59]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_58 = csr_status[58]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_57 = csr_status[57]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_56 = csr_status[56]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_55 = csr_status[55]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_54 = csr_status[54]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_53 = csr_status[53]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_52 = csr_status[52]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_51 = csr_status[51]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_50 = csr_status[50]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_49 = csr_status[49]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_48 = csr_status[48]; // @[csr.scala 175:28]
  wire [7:0] csr_status_to_be_hi_hi_lo = {csr_status_to_vec_55,csr_status_to_vec_54,csr_status_to_vec_53,
    csr_status_to_vec_52,csr_status_to_vec_51,csr_status_to_vec_50,csr_status_to_vec_49,csr_status_to_vec_48}; // @[csr.scala 182:53]
  wire  csr_status_to_vec_47 = csr_status[47]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_46 = csr_status[46]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_45 = csr_status[45]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_44 = csr_status[44]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_43 = csr_status[43]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_42 = csr_status[42]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_41 = csr_status[41]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_40 = csr_status[40]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_39 = csr_status[39]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_38 = csr_status[38]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_37 = csr_status[37]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_36 = csr_status[36]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_35 = csr_status[35]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_34 = csr_status[34]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_33 = csr_status[33]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_32 = csr_status[32]; // @[csr.scala 175:28]
  wire [7:0] csr_status_to_be_hi_lo_lo = {csr_status_to_vec_39,csr_status_to_vec_38,csr_status_to_vec_37,
    csr_status_to_vec_36,csr_status_to_vec_35,csr_status_to_vec_34,csr_status_to_vec_33,csr_status_to_vec_32}; // @[csr.scala 182:53]
  wire [15:0] csr_status_to_be_hi_lo = {csr_status_to_vec_47,csr_status_to_vec_46,csr_status_to_vec_45,
    csr_status_to_vec_44,csr_status_to_vec_43,csr_status_to_vec_42,csr_status_to_vec_41,csr_status_to_vec_40,
    csr_status_to_be_hi_lo_lo}; // @[csr.scala 182:53]
  wire [31:0] csr_status_to_be_hi = {csr_status_to_vec_63,csr_status_to_vec_62,csr_status_to_vec_61,csr_status_to_vec_60
    ,csr_status_to_vec_59,csr_status_to_vec_58,csr_status_to_vec_57,csr_status_to_vec_56,csr_status_to_be_hi_hi_lo,
    csr_status_to_be_hi_lo}; // @[csr.scala 182:53]
  wire  csr_status_to_vec_31 = csr_status[31]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_30 = csr_status[30]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_29 = csr_status[29]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_28 = csr_status[28]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_27 = csr_status[27]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_26 = csr_status[26]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_25 = csr_status[25]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_24 = csr_status[24]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_23 = csr_status[23]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_22 = csr_status[22]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_21 = csr_status[21]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_20 = csr_status[20]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_19 = csr_status[19]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_18 = csr_status[18]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_17 = csr_status[17]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_16 = csr_status[16]; // @[csr.scala 175:28]
  wire [7:0] csr_status_to_be_lo_hi_lo = {csr_status_to_vec_23,csr_status_to_vec_22,csr_status_to_vec_21,
    csr_status_to_vec_20,csr_status_to_vec_19,csr_status_to_vec_18,csr_status_to_vec_17,csr_status_to_vec_16}; // @[csr.scala 182:53]
  wire  csr_status_to_vec_15 = csr_status[15]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_14 = csr_status[14]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_13 = csr_status[13]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_12 = csr_status[12]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_11 = csr_status[11]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_10 = csr_status[10]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_9 = csr_status[9]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_8 = csr_status[8]; // @[csr.scala 175:28]
  reg [63:0] csr_mie; // @[csr.scala 73:28]
  wire  _commit_int_T_3 = io_int_type_out_int & csr_mie[11]; // @[csr.scala 89:44]
  wire  _commit_int_T_4 = io_int_type_timer & csr_mie[7] | _commit_int_T_3; // @[csr.scala 88:60]
  wire  commit_int = _commit_int_T_4 & csr_status[3] & io_stageW_pc != 64'h0; // @[csr.scala 89:92]
  wire [31:0] exception_type = {io_exception_type_i,commit_int}; // @[Cat.scala 31:58]
  wire  commit_eret = exception_type[31]; // @[csr.scala 94:38]
  wire  csr_status_to_vec_7 = commit_eret | csr_status[7]; // @[csr.scala 173:21]
  wire  csr_status_to_vec_6 = csr_status[6]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_5 = csr_status[5]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_4 = csr_status[4]; // @[csr.scala 175:28]
  wire  _csr_status_to_vec_3_T_3 = commit_eret ? csr_status[7] : csr_status[3]; // @[csr.scala 171:20]
  wire  csr_status_to_vec_3 = commit_int ? 1'h0 : _csr_status_to_vec_3_T_3; // @[csr.scala 170:21]
  wire  csr_status_to_vec_2 = csr_status[2]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_1 = csr_status[1]; // @[csr.scala 175:28]
  wire  csr_status_to_vec_0 = csr_status[0]; // @[csr.scala 175:28]
  wire [7:0] csr_status_to_be_lo_lo_lo = {csr_status_to_vec_7,csr_status_to_vec_6,csr_status_to_vec_5,
    csr_status_to_vec_4,csr_status_to_vec_3,csr_status_to_vec_2,csr_status_to_vec_1,csr_status_to_vec_0}; // @[csr.scala 182:53]
  wire [15:0] csr_status_to_be_lo_lo = {csr_status_to_vec_15,csr_status_to_vec_14,csr_status_to_vec_13,
    csr_status_to_vec_12,csr_status_to_vec_11,csr_status_to_vec_10,csr_status_to_vec_9,csr_status_to_vec_8,
    csr_status_to_be_lo_lo_lo}; // @[csr.scala 182:53]
  wire [31:0] csr_status_to_be_lo = {csr_status_to_vec_31,csr_status_to_vec_30,csr_status_to_vec_29,csr_status_to_vec_28
    ,csr_status_to_vec_27,csr_status_to_vec_26,csr_status_to_vec_25,csr_status_to_vec_24,csr_status_to_be_lo_hi_lo,
    csr_status_to_be_lo_lo}; // @[csr.scala 182:53]
  wire [63:0] _csr_status_to_be_T = {csr_status_to_be_hi,csr_status_to_be_lo}; // @[csr.scala 182:53]
  reg [63:0] csr_epc; // @[csr.scala 65:26]
  reg [63:0] csr_mtvec; // @[csr.scala 66:28]
  reg [63:0] csr_mip; // @[csr.scala 74:28]
  wire [31:0] _commit_exception_T_2 = {{24'd0}, exception_type[31:24]}; // @[csr.scala 93:76]
  wire  commit_exception = exception_type[30:0] != 31'h0 & ~_commit_exception_T_2[0]; // @[csr.scala 93:58]
  wire [63:0] _csr_read_data_Wire_T_1 = 12'h341 == io_csr_read_addr ? csr_epc : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_3 = 12'h342 == io_csr_read_addr ? csr_cause : _csr_read_data_Wire_T_1; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_5 = 12'h305 == io_csr_read_addr ? csr_mtvec : _csr_read_data_Wire_T_3; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_7 = 12'h300 == io_csr_read_addr ? csr_status : _csr_read_data_Wire_T_5; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_9 = 12'h344 == io_csr_read_addr ? csr_mip : _csr_read_data_Wire_T_7; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_11 = 12'h304 == io_csr_read_addr ? csr_mie : _csr_read_data_Wire_T_9; // @[Mux.scala 81:58]
  wire [63:0] csr_read_data_Wire = 12'hf14 == io_csr_read_addr ? 64'h0 : _csr_read_data_Wire_T_11; // @[Mux.scala 81:58]
  wire [63:0] _io_return_pc_T_2 = io_pc + 64'h4; // @[csr.scala 109:38]
  wire [63:0] _io_return_pc_T_3 = _commit_exception_T_2[0] ? _io_return_pc_T_2 : csr_mtvec; // @[Mux.scala 101:16]
  wire [62:0] _int_code_T = io_int_type_timer ? 63'h7 : 63'h0; // @[Mux.scala 27:73]
  wire [62:0] _int_code_T_1 = io_int_type_out_int ? 63'hb : 63'h0; // @[Mux.scala 27:73]
  wire [62:0] int_code = _int_code_T | _int_code_T_1; // @[Mux.scala 27:73]
  wire [63:0] _cause_exccode_T_2 = {1'h1,int_code}; // @[Cat.scala 31:58]
  wire [31:0] _cause_exccode_T_3 = {{8'd0}, exception_type[31:8]}; // @[csr.scala 123:23]
  wire [63:0] _cause_exccode_T_5 = exception_type[0] ? _cause_exccode_T_2 : 64'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_T_6 = _cause_exccode_T_3[0] ? 4'hb : 4'h0; // @[Mux.scala 27:73]
  wire [63:0] _GEN_3 = {{60'd0}, _cause_exccode_T_6}; // @[Mux.scala 27:73]
  wire [63:0] cause_exccode = _cause_exccode_T_5 | _GEN_3; // @[Mux.scala 27:73]
  wire  _csr_epc_T_3 = io_csr_write_en & io_csr_write_addr == 12'h341; // @[csr.scala 180:32]
  wire  _csr_mtvec_T_2 = io_csr_write_en & io_csr_write_addr == 12'h305; // @[csr.scala 187:33]
  wire  _csr_cause_T_2 = io_csr_write_en & io_csr_write_addr == 12'h342; // @[csr.scala 191:33]
  wire  _csr_mie_T_2 = io_csr_write_en & io_csr_write_addr == 12'h304; // @[csr.scala 195:33]
  wire  csr_mip_to_be_7 = commit_int ? io_int_type_timer : csr_mip[7]; // @[csr.scala 202:36]
  wire  csr_mip_to_be_11 = commit_int ? io_int_type_out_int : csr_mip[11]; // @[csr.scala 203:42]
  wire [63:0] _csr_mip_T = {32'h0,16'h0,4'h0,csr_mip_to_be_11,1'h0,2'h0,csr_mip_to_be_7,1'h0,2'h0,4'h0}; // @[csr.scala 206:42]
  wire  _csr_mip_T_3 = io_csr_write_en & io_csr_write_addr == 12'h344; // @[csr.scala 207:33]
  assign io_return_pc = commit_eret ? csr_epc : _io_return_pc_T_3; // @[Mux.scala 101:16]
  assign io_exception = commit_exception | commit_eret; // @[csr.scala 96:43]
  assign io_csr_read_data = reset ? 64'h0 : csr_read_data_Wire; // @[csr.scala 103:29]
  assign io_icache_tags_flush = _commit_exception_T_2[0]; // @[csr.scala 95:40]
  assign io_Int_able = csr_status[3]; // @[csr.scala 164:30]
  assign io_int_type_able_timer = csr_mie[7]; // @[csr.scala 198:38]
  assign io_int_type_able_out_int = csr_mie[11]; // @[csr.scala 199:40]
  always @(posedge clock) begin
    if (reset) begin // @[csr.scala 61:28]
      csr_cause <= 64'h400000; // @[csr.scala 61:28]
    end else if (_csr_cause_T_2) begin // @[Mux.scala 101:16]
      csr_cause <= io_csr_write_data;
    end else if (commit_exception) begin // @[Mux.scala 101:16]
      csr_cause <= cause_exccode;
    end
    if (reset) begin // @[csr.scala 64:22]
      csr_status <= 64'ha00001800;
    end else if (_csr_status_to_be_T_3) begin // @[Mux.scala 101:16]
      csr_status <= io_csr_write_data;
    end else begin
      csr_status <= _csr_status_to_be_T;
    end
    if (reset) begin // @[csr.scala 73:28]
      csr_mie <= 64'h0; // @[csr.scala 73:28]
    end else if (_csr_mie_T_2) begin // @[Mux.scala 101:16]
      csr_mie <= io_csr_write_data;
    end
    if (reset) begin // @[csr.scala 65:26]
      csr_epc <= 64'h0; // @[csr.scala 65:26]
    end else if (commit_exception) begin // @[Mux.scala 101:16]
      csr_epc <= io_pc;
    end else if (_csr_epc_T_3) begin // @[Mux.scala 101:16]
      csr_epc <= io_csr_write_data;
    end
    if (reset) begin // @[csr.scala 66:28]
      csr_mtvec <= 64'h0; // @[csr.scala 66:28]
    end else if (_csr_mtvec_T_2) begin // @[Mux.scala 101:16]
      csr_mtvec <= io_csr_write_data;
    end
    if (reset) begin // @[csr.scala 74:28]
      csr_mip <= 64'h0; // @[csr.scala 74:28]
    end else if (_csr_mip_T_3) begin // @[Mux.scala 101:16]
      csr_mip <= io_csr_write_data;
    end else begin
      csr_mip <= _csr_mip_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  csr_cause = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  csr_status = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  csr_mie = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  csr_epc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  csr_mtvec = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  csr_mip = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_cu(
  input  [31:0] io1_InstrD,
  output        io1_BadInstrD,
  output        io1_SysCallD,
  output        io1_EretD,
  output        io1_dmem_addr_cal,
  output        io_RegWriteD,
  output        io_MemToRegD,
  output        io_MemWriteD,
  output [15:0] io_ALUCtrlD,
  output        io_ALUSrcD_0,
  output        io_ALUSrcD_1,
  output [4:0]  io_RegDstD,
  output        io_LinkD,
  output        io_csrWriteD,
  output        io_csrToRegD,
  output        io_LoadUnsignedD,
  output [1:0]  io_MemWidthD,
  output [63:0] io_ImmD,
  output        io_data_wD,
  output [23:0] io_muldiv_control,
  output        io_muldiv_cal,
  output        io_alu_cal,
  output [2:0]  io_csr_control,
  output        io_csr_Imm,
  output        io_fence_i_control
);
  wire [6:0] OpD = io1_InstrD[6:0]; // @[cu.scala 63:25]
  wire [2:0] Funct3D = io1_InstrD[14:12]; // @[cu.scala 64:29]
  wire [6:0] Funct7D = io1_InstrD[31:25]; // @[cu.scala 65:29]
  wire [5:0] Funct6D = io1_InstrD[31:26]; // @[cu.scala 66:29]
  wire [5:0] immI_lo_lo_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31]}
    ; // @[Cat.scala 31:58]
  wire [12:0] immI_lo_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] immI_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo,immI_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _immI_T_53 = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo,immI_lo_lo,immI_lo}; // @[Cat.scala 31:58]
  wire [63:0] immI = {_immI_T_53,io1_InstrD[31:20]}; // @[Cat.scala 31:58]
  wire [11:0] _immS_T_2 = {Funct7D,io1_InstrD[11:7]}; // @[Cat.scala 31:58]
  wire [5:0] immS_lo_lo_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11]}; // @[Cat.scala 31:58]
  wire [12:0] immS_lo_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],
    _immS_T_2[11],immS_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] immS_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[
    11],immS_lo_lo_lo,immS_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _immS_T_55 = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],
    _immS_T_2[11],immS_lo_lo_lo,immS_lo_lo,immS_lo}; // @[Cat.scala 31:58]
  wire [63:0] immS = {_immS_T_55,Funct7D,io1_InstrD[11:7]}; // @[Cat.scala 31:58]
  wire [31:0] _immU_T_1 = {io1_InstrD[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [7:0] immU_lo_lo = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1
    [31],_immU_T_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] immU_lo = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[
    31],_immU_T_1[31],immU_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _immU_T_34 = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],
    _immU_T_1[31],_immU_T_1[31],immU_lo_lo,immU_lo}; // @[Cat.scala 31:58]
  wire [63:0] immU = {_immU_T_34,io1_InstrD[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [12:0] _immSB_T_4 = {io1_InstrD[31],io1_InstrD[7],io1_InstrD[30:25],io1_InstrD[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [5:0] immSB_lo_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12]
    }; // @[Cat.scala 31:58]
  wire [11:0] immSB_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [12:0] immSB_lo_hi = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [24:0] immSB_lo_1 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_lo}; // @[Cat.scala 31:58]
  wire [50:0] _immSB_T_56 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_hi,immSB_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] immSB = {_immSB_T_56,io1_InstrD[31],io1_InstrD[7],io1_InstrD[30:25],io1_InstrD[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] immUJ = {io1_InstrD[31],io1_InstrD[19:12],io1_InstrD[20],io1_InstrD[30:21]}; // @[Cat.scala 31:58]
  wire [3:0] _inst_code_type_T_2 = 7'h0 == Funct7D ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_4 = 6'h0 == Funct6D ? 5'h13 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_6 = 6'h10 == Funct6D ? 5'h14 : _inst_code_type_T_4; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_8 = 3'h2 == Funct3D ? 4'hd : 4'h4; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_10 = 3'h3 == Funct3D ? 4'he : _inst_code_type_T_8; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_12 = 3'h4 == Funct3D ? 5'h17 : {{1'd0}, _inst_code_type_T_10}; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_14 = 3'h6 == Funct3D ? 5'h16 : _inst_code_type_T_12; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_16 = 3'h7 == Funct3D ? 5'h15 : _inst_code_type_T_14; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_18 = 3'h1 == Funct3D ? {{1'd0}, _inst_code_type_T_2} : _inst_code_type_T_16; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_20 = 3'h1 == Funct3D ? 5'hf : _inst_code_type_T_18; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_22 = 3'h5 == Funct3D ? _inst_code_type_T_6 : _inst_code_type_T_20; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_23 = {_inst_code_type_T_22,3'h2}; // @[Cat.scala 31:58]
  wire [5:0] _inst_code_type_T_25 = 7'h20 == Funct7D ? 6'h36 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_27 = 7'h0 == Funct7D ? 6'h30 : _inst_code_type_T_25; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_29 = 7'h1 == Funct7D ? 6'h2c : _inst_code_type_T_27; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_31 = 7'h0 == Funct7D ? 6'h31 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_33 = 7'h1 == Funct7D ? 6'h2d : _inst_code_type_T_31; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_35 = 7'h1 == Funct7D ? 6'h2f : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_37 = 7'h0 == Funct7D ? 6'h34 : _inst_code_type_T_35; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_39 = 7'h0 == Funct7D ? 6'h35 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_41 = 7'h1 == Funct7D ? 6'h2e : _inst_code_type_T_39; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_43 = 7'h0 == Funct7D ? 7'h41 : 7'h0; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_45 = 7'h1 == Funct7D ? 7'h24 : _inst_code_type_T_43; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_47 = 7'h0 == Funct7D ? 6'h32 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_49 = 7'h1 == Funct7D ? 6'h23 : _inst_code_type_T_47; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_51 = 7'h20 == Funct7D ? 6'h33 : _inst_code_type_T_49; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_53 = 7'h0 == Funct7D ? 6'h38 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_55 = 7'h1 == Funct7D ? 6'h26 : _inst_code_type_T_53; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_57 = 7'h0 == Funct7D ? 6'h37 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_59 = 7'h1 == Funct7D ? 6'h25 : _inst_code_type_T_57; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_61 = 3'h1 == Funct3D ? _inst_code_type_T_33 : _inst_code_type_T_29; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_63 = 3'h2 == Funct3D ? _inst_code_type_T_37 : _inst_code_type_T_61; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_65 = 3'h3 == Funct3D ? _inst_code_type_T_41 : _inst_code_type_T_63; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_67 = 3'h4 == Funct3D ? _inst_code_type_T_45 : {{1'd0}, _inst_code_type_T_65}; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_69 = 3'h5 == Funct3D ? {{1'd0}, _inst_code_type_T_51} : _inst_code_type_T_67; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_71 = 3'h6 == Funct3D ? {{1'd0}, _inst_code_type_T_55} : _inst_code_type_T_69; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_73 = 3'h7 == Funct3D ? {{1'd0}, _inst_code_type_T_59} : _inst_code_type_T_71; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_74 = {_inst_code_type_T_73,3'h5}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_76 = 3'h0 == Funct3D ? 5'h1c : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_78 = 3'h1 == Funct3D ? 5'h1d : _inst_code_type_T_76; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_80 = 3'h4 == Funct3D ? 6'h20 : {{1'd0}, _inst_code_type_T_78}; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_82 = 3'h5 == Funct3D ? 6'h1e : _inst_code_type_T_80; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_84 = 3'h6 == Funct3D ? 6'h21 : _inst_code_type_T_82; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_86 = 3'h7 == Funct3D ? 6'h1f : _inst_code_type_T_84; // @[Mux.scala 81:58]
  wire [8:0] _inst_code_type_T_87 = {_inst_code_type_T_86,3'h4}; // @[Cat.scala 31:58]
  wire [3:0] _inst_code_type_T_93 = 3'h0 == Funct3D ? 4'h8 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_95 = 3'h1 == Funct3D ? 4'ha : _inst_code_type_T_93; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_97 = 3'h2 == Funct3D ? 4'hc : _inst_code_type_T_95; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_99 = 3'h4 == Funct3D ? 4'h7 : _inst_code_type_T_97; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_101 = 3'h5 == Funct3D ? 4'h9 : _inst_code_type_T_99; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_103 = 3'h6 == Funct3D ? 4'hb : _inst_code_type_T_101; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_105 = 3'h3 == Funct3D ? 4'h6 : _inst_code_type_T_103; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_106 = {_inst_code_type_T_105,3'h2}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_108 = 3'h0 == Funct3D ? 5'h18 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_110 = 3'h1 == Funct3D ? 5'h19 : _inst_code_type_T_108; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_112 = 3'h2 == Funct3D ? 5'h1a : _inst_code_type_T_110; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_114 = 3'h3 == Funct3D ? 5'h1b : _inst_code_type_T_112; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_115 = {_inst_code_type_T_114,3'h3}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_117 = 7'h0 == Funct7D ? 5'h11 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_119 = 7'h20 == Funct7D ? 5'h12 : _inst_code_type_T_117; // @[Mux.scala 81:58]
  wire [2:0] _inst_code_type_T_121 = 3'h0 == Funct3D ? 3'h5 : 3'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_123 = 3'h1 == Funct3D ? 5'h10 : {{2'd0}, _inst_code_type_T_121}; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_125 = 3'h5 == Funct3D ? _inst_code_type_T_119 : _inst_code_type_T_123; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_126 = {_inst_code_type_T_125,3'h2}; // @[Cat.scala 31:58]
  wire [5:0] _inst_code_type_T_128 = 7'h0 == Funct7D ? 6'h3c : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_130 = 7'h20 == Funct7D ? 6'h3d : _inst_code_type_T_128; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_132 = 7'h1 == Funct7D ? 6'h2b : _inst_code_type_T_130; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_134 = 7'h0 == Funct7D ? 6'h39 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_136 = 7'h0 == Funct7D ? 6'h3a : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_138 = 7'h20 == Funct7D ? 6'h3b : _inst_code_type_T_136; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_140 = 7'h1 == Funct7D ? 6'h28 : _inst_code_type_T_138; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_142 = 3'h0 == Funct3D ? _inst_code_type_T_132 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_144 = 3'h1 == Funct3D ? _inst_code_type_T_134 : _inst_code_type_T_142; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_146 = 3'h5 == Funct3D ? _inst_code_type_T_140 : _inst_code_type_T_144; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_148 = 3'h6 == Funct3D ? 6'h29 : _inst_code_type_T_146; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_150 = 3'h7 == Funct3D ? 6'h2a : _inst_code_type_T_148; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_152 = 3'h4 == Funct3D ? 6'h27 : _inst_code_type_T_150; // @[Mux.scala 81:58]
  wire [8:0] _inst_code_type_T_153 = {_inst_code_type_T_152,3'h5}; // @[Cat.scala 31:58]
  wire [6:0] _inst_code_type_T_156 = 7'h0 == Funct7D ? 7'h4c : 7'h0; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_158 = 7'h18 == Funct7D ? 7'h4d : _inst_code_type_T_156; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_159 = {_inst_code_type_T_158,3'h0}; // @[Cat.scala 31:58]
  wire [9:0] _inst_code_type_T_167 = 3'h0 == Funct3D ? _inst_code_type_T_159 : 10'h0; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_169 = 3'h1 == Funct3D ? 10'h25a : _inst_code_type_T_167; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_171 = 3'h2 == Funct3D ? 10'h252 : _inst_code_type_T_169; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_173 = 3'h3 == Funct3D ? 10'h24a : _inst_code_type_T_171; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_175 = 3'h5 == Funct3D ? 10'h242 : _inst_code_type_T_173; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_177 = 3'h6 == Funct3D ? 10'h23a : _inst_code_type_T_175; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_179 = 3'h7 == Funct3D ? 10'h232 : _inst_code_type_T_177; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_182 = 3'h1 == Funct3D ? 10'h277 : 10'h0; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_184 = 7'h13 == OpD ? _inst_code_type_T_23 : 8'h0; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_186 = 7'h33 == OpD ? _inst_code_type_T_74 : {{2'd0}, _inst_code_type_T_184}; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_188 = 7'h63 == OpD ? {{1'd0}, _inst_code_type_T_87} : _inst_code_type_T_186; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_190 = 7'h6f == OpD ? 10'h16 : _inst_code_type_T_188; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_192 = 7'h67 == OpD ? 10'h1a : _inst_code_type_T_190; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_194 = 7'h37 == OpD ? 10'h9 : _inst_code_type_T_192; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_196 = 7'h17 == OpD ? 10'h201 : _inst_code_type_T_194; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_198 = 7'h3 == OpD ? {{3'd0}, _inst_code_type_T_106} : _inst_code_type_T_196; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_200 = 7'h23 == OpD ? {{2'd0}, _inst_code_type_T_115} : _inst_code_type_T_198; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_202 = 7'h1b == OpD ? {{2'd0}, _inst_code_type_T_126} : _inst_code_type_T_200; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_204 = 7'h3b == OpD ? {{1'd0}, _inst_code_type_T_153} : _inst_code_type_T_202; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_206 = 7'h0 == OpD ? 10'h282 : _inst_code_type_T_204; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_208 = 7'h73 == OpD ? _inst_code_type_T_179 : _inst_code_type_T_206; // @[Mux.scala 81:58]
  wire [9:0] inst_code_type = 7'hf == OpD ? _inst_code_type_T_182 : _inst_code_type_T_208; // @[Mux.scala 81:58]
  wire [6:0] ins_code = inst_code_type[9:3]; // @[cu.scala 195:35]
  wire [2:0] inst_type = inst_code_type[2:0]; // @[cu.scala 196:35]
  wire [3:0] _io_csr_control_T_7 = 7'h4b == ins_code ? 4'h4 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_9 = 7'h48 == ins_code ? 4'h4 : _io_csr_control_T_7; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_11 = 7'h49 == ins_code ? 4'h2 : _io_csr_control_T_9; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_13 = 7'h46 == ins_code ? 4'h2 : _io_csr_control_T_11; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_15 = 7'h4a == ins_code ? 4'h1 : _io_csr_control_T_13; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_17 = 7'h47 == ins_code ? 4'h1 : _io_csr_control_T_15; // @[Mux.scala 81:58]
  wire  _io_ImmD_T = inst_type == 3'h1; // @[cu.scala 236:20]
  wire  _io_ImmD_T_1 = inst_type == 3'h2; // @[cu.scala 237:20]
  wire  _io_ImmD_T_2 = inst_type == 3'h3; // @[cu.scala 238:20]
  wire  _io_ImmD_T_3 = inst_type == 3'h4; // @[cu.scala 239:20]
  wire  _io_ImmD_T_4 = inst_type == 3'h6; // @[cu.scala 240:20]
  wire [63:0] _io_ImmD_T_5 = _io_ImmD_T ? immU : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_6 = _io_ImmD_T_1 ? immI : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_7 = _io_ImmD_T_2 ? immS : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_8 = _io_ImmD_T_3 ? immSB : 64'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_ImmD_T_9 = _io_ImmD_T_4 ? immUJ : 20'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_10 = _io_ImmD_T_5 | _io_ImmD_T_6; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_11 = _io_ImmD_T_10 | _io_ImmD_T_7; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_12 = _io_ImmD_T_11 | _io_ImmD_T_8; // @[Mux.scala 27:73]
  wire [63:0] _GEN_0 = {{44'd0}, _io_ImmD_T_9}; // @[Mux.scala 27:73]
  wire  _io_RegWriteD_T_29 = 7'h30 == ins_code | (7'h2b == ins_code | (7'h2f == ins_code | (7'h2e == ins_code | (7'h2d
     == ins_code | (7'h2c == ins_code | (7'h2b == ins_code | (7'h2a == ins_code | (7'h29 == ins_code | (7'h28 ==
    ins_code | (7'h27 == ins_code | (7'h26 == ins_code | (7'h25 == ins_code | (7'h24 == ins_code | 7'h23 == ins_code))))
    ))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_59 = 7'h2 == ins_code | (7'h3 == ins_code | (7'h3d == ins_code | (7'h3c == ins_code | (7'h3b ==
    ins_code | (7'h3a == ins_code | (7'h39 == ins_code | (7'h38 == ins_code | (7'h37 == ins_code | (7'h36 == ins_code |
    (7'h35 == ins_code | (7'h34 == ins_code | (7'h33 == ins_code | (7'h32 == ins_code | (7'h31 == ins_code |
    _io_RegWriteD_T_29)))))))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_89 = 7'h10 == ins_code | (7'hf == ins_code | (7'he == ins_code | (7'hd == ins_code | (7'h9 ==
    ins_code | (7'h7 == ins_code | (7'hc == ins_code | (7'hb == ins_code | (7'ha == ins_code | (7'h9 == ins_code | (7'h8
     == ins_code | (7'h7 == ins_code | (7'h6 == ins_code | (7'h5 == ins_code | (7'h4 == ins_code | _io_RegWriteD_T_59)))
    ))))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_119 = 7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a == ins_code | (7'h49
     == ins_code | (7'h1 == ins_code | (7'h40 == ins_code | (7'h41 == ins_code | (7'h17 == ins_code | (7'h16 == ins_code
     | (7'h15 == ins_code | (7'h14 == ins_code | (7'h13 == ins_code | (7'h12 == ins_code | (7'h11 == ins_code |
    _io_RegWriteD_T_89)))))))))))))); // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_33 = 7'h40 == ins_code ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_35 = 7'h30 == ins_code ? 2'h2 : _io_ALUCtrlD_T_33; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_37 = 7'h5 == ins_code ? 2'h2 : _io_ALUCtrlD_T_35; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_39 = 7'h4 == ins_code ? 2'h2 : _io_ALUCtrlD_T_37; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_41 = 7'h3c == ins_code ? 2'h2 : _io_ALUCtrlD_T_39; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_43 = 7'hd == ins_code ? 16'h2000 : {{14'd0}, _io_ALUCtrlD_T_41}; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_45 = 7'he == ins_code ? 16'h4000 : _io_ALUCtrlD_T_43; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_47 = 7'hf == ins_code ? 16'h1000 : _io_ALUCtrlD_T_45; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_49 = 7'h10 == ins_code ? 16'h1000 : _io_ALUCtrlD_T_47; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_51 = 7'h11 == ins_code ? 16'h20 : _io_ALUCtrlD_T_49; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_53 = 7'h12 == ins_code ? 16'h8000 : _io_ALUCtrlD_T_51; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_55 = 7'h13 == ins_code ? 16'h20 : _io_ALUCtrlD_T_53; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_57 = 7'h14 == ins_code ? 16'h8000 : _io_ALUCtrlD_T_55; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_59 = 7'h15 == ins_code ? 16'h10 : _io_ALUCtrlD_T_57; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_61 = 7'h16 == ins_code ? 16'h800 : _io_ALUCtrlD_T_59; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_63 = 7'h17 == ins_code ? 16'h1 : _io_ALUCtrlD_T_61; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_65 = 7'h1 == ins_code ? 16'h80 : _io_ALUCtrlD_T_63; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_67 = 7'h30 == ins_code ? 16'h2 : _io_ALUCtrlD_T_65; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_69 = 7'h31 == ins_code ? 16'h1000 : _io_ALUCtrlD_T_67; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_71 = 7'h32 == ins_code ? 16'h20 : _io_ALUCtrlD_T_69; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_73 = 7'h33 == ins_code ? 16'h8000 : _io_ALUCtrlD_T_71; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_75 = 7'h34 == ins_code ? 16'h2000 : _io_ALUCtrlD_T_73; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_77 = 7'h35 == ins_code ? 16'h4000 : _io_ALUCtrlD_T_75; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_79 = 7'h36 == ins_code ? 16'h40 : _io_ALUCtrlD_T_77; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_81 = 7'h37 == ins_code ? 16'h10 : _io_ALUCtrlD_T_79; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_83 = 7'h38 == ins_code ? 16'h800 : _io_ALUCtrlD_T_81; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_85 = 7'h39 == ins_code ? 16'h1000 : _io_ALUCtrlD_T_83; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_87 = 7'h3a == ins_code ? 16'h20 : _io_ALUCtrlD_T_85; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_89 = 7'h3b == ins_code ? 16'h8000 : _io_ALUCtrlD_T_87; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_91 = 7'h3c == ins_code ? 16'h2 : _io_ALUCtrlD_T_89; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_93 = 7'h3d == ins_code ? 16'h40 : _io_ALUCtrlD_T_91; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_5 = 3'h2 == Funct3D ? 2'h2 : {{1'd0}, 3'h1 == Funct3D}; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_7 = 3'h4 == Funct3D ? 2'h0 : _io_MemWidthD_T_5; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_9 = 3'h5 == Funct3D ? 2'h1 : _io_MemWidthD_T_7; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_11 = 3'h6 == Funct3D ? 2'h2 : _io_MemWidthD_T_9; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_13 = 3'h3 == Funct3D ? 2'h3 : _io_MemWidthD_T_11; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_21 = 3'h3 == Funct3D ? 2'h3 : _io_MemWidthD_T_5; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_23 = 7'h3 == OpD ? _io_MemWidthD_T_13 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_muldiv_control_T_14 = 7'h24 == ins_code ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_muldiv_control_T_16 = 7'h23 == ins_code ? 2'h1 : _io_muldiv_control_T_14; // @[Mux.scala 81:58]
  wire [3:0] _io_muldiv_control_T_18 = 7'h25 == ins_code ? 4'h4 : {{2'd0}, _io_muldiv_control_T_16}; // @[Mux.scala 81:58]
  wire [3:0] _io_muldiv_control_T_20 = 7'h26 == ins_code ? 4'h8 : _io_muldiv_control_T_18; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_22 = 7'h27 == ins_code ? 8'h10 : {{4'd0}, _io_muldiv_control_T_20}; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_24 = 7'h28 == ins_code ? 8'h20 : _io_muldiv_control_T_22; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_26 = 7'h29 == ins_code ? 8'h40 : _io_muldiv_control_T_24; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_28 = 7'h2a == ins_code ? 8'h80 : _io_muldiv_control_T_26; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_30 = 7'h2b == ins_code ? 16'h100 : {{8'd0}, _io_muldiv_control_T_28}; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_32 = 7'h2c == ins_code ? 16'h200 : _io_muldiv_control_T_30; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_34 = 7'h2d == ins_code ? 16'h400 : _io_muldiv_control_T_32; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_36 = 7'h2f == ins_code ? 16'h1000 : _io_muldiv_control_T_34; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_38 = 7'h2e == ins_code ? 16'h800 : _io_muldiv_control_T_36; // @[Mux.scala 81:58]
  assign io1_BadInstrD = ins_code == 7'h0; // @[cu.scala 260:31]
  assign io1_SysCallD = ins_code == 7'h4c; // @[cu.scala 261:31]
  assign io1_EretD = ins_code == 7'h4d; // @[cu.scala 262:31]
  assign io1_dmem_addr_cal = 7'h23 == OpD ? 3'h3 == Funct3D | (3'h2 == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D)) : 7'h3
     == OpD & (3'h3 == Funct3D | (3'h6 == Funct3D | (3'h5 == Funct3D | (3'h4 == Funct3D | (3'h2 == Funct3D | (3'h1 ==
    Funct3D | 3'h0 == Funct3D)))))); // @[Mux.scala 81:58]
  assign io_RegWriteD = 7'h46 == ins_code | _io_RegWriteD_T_119; // @[Mux.scala 81:58]
  assign io_MemToRegD = 7'h3 == OpD & (3'h3 == Funct3D | (3'h6 == Funct3D | (3'h5 == Funct3D | (3'h4 == Funct3D | (3'h2
     == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D)))))); // @[Mux.scala 81:58]
  assign io_MemWriteD = 7'h23 == OpD & (3'h3 == Funct3D | (3'h2 == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D))); // @[Mux.scala 81:58]
  assign io_ALUCtrlD = 7'h41 == ins_code ? 16'h1 : _io_ALUCtrlD_T_93; // @[Mux.scala 81:58]
  assign io_ALUSrcD_0 = ins_code == 7'h40; // @[cu.scala 362:32]
  assign io_ALUSrcD_1 = _io_ImmD_T_1 | _io_ImmD_T_4 | _io_ImmD_T; // @[cu.scala 364:79]
  assign io_RegDstD = io1_InstrD[11:7]; // @[cu.scala 76:29]
  assign io_LinkD = ins_code == 7'h3 | ins_code == 7'h2; // @[cu.scala 242:38]
  assign io_csrWriteD = 7'h46 == ins_code | (7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a ==
    ins_code | 7'h49 == ins_code)))); // @[Mux.scala 81:58]
  assign io_csrToRegD = 7'h46 == ins_code | (7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a ==
    ins_code | 7'h49 == ins_code)))); // @[Mux.scala 81:58]
  assign io_LoadUnsignedD = 7'h3 == OpD & (3'h6 == Funct3D | (3'h5 == Funct3D | 3'h4 == Funct3D)); // @[Mux.scala 81:58]
  assign io_MemWidthD = 7'h23 == OpD ? _io_MemWidthD_T_21 : _io_MemWidthD_T_23; // @[Mux.scala 81:58]
  assign io_ImmD = _io_ImmD_T_12 | _GEN_0; // @[Mux.scala 27:73]
  assign io_data_wD = 7'h12 == ins_code | (7'h11 == ins_code | (7'h10 == ins_code | (7'h5 == ins_code | (7'h3d ==
    ins_code | (7'h3c == ins_code | (7'h3b == ins_code | (7'h3a == ins_code | (7'h39 == ins_code | (7'h2b == ins_code |
    (7'h2b == ins_code | (7'h2a == ins_code | (7'h29 == ins_code | (7'h28 == ins_code | 7'h27 == ins_code))))))))))))); // @[Mux.scala 81:58]
  assign io_muldiv_control = {{8'd0}, _io_muldiv_control_T_38}; // @[cu.scala 475:23]
  assign io_muldiv_cal = io_muldiv_control != 24'h0; // @[cu.scala 491:40]
  assign io_alu_cal = io_ALUCtrlD != 16'h0; // @[cu.scala 492:34]
  assign io_csr_control = _io_csr_control_T_17[2:0]; // @[cu.scala 217:20]
  assign io_csr_Imm = ins_code == 7'h48 | ins_code == 7'h46 | ins_code == 7'h47; // @[cu.scala 225:72]
  assign io_fence_i_control = io1_InstrD == 32'h100f; // @[cu.scala 198:39]
endmodule
module ysyx_22040886_dmem(
  input         io_data_ok,
  input  [63:0] io_rdata,
  input  [2:0]  io_Physisc_Address,
  input  [1:0]  io_WIDTH,
  input         io_SIGN,
  output [63:0] io_RD,
  output        io_data_pending
);
  wire [1:0] ra = io_Physisc_Address[1:0]; // @[dmem.scala 39:32]
  wire  third_ra = io_Physisc_Address[2]; // @[dmem.scala 40:38]
  wire [2:0] _io_RD_T_1 = {ra,io_SIGN}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39
    ]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo,io_RD_lo_lo}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_59 = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo,io_RD_lo_lo,io_RD_lo}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_61 = {_io_RD_T_59,io_rdata[39:32]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_64 = {1'h0,io_rdata[39:32]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[
    47]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47
    ],io_RD_lo_lo_lo_1}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_1,io_RD_lo_lo_1}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_122 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47]
    ,io_RD_lo_lo_lo_1,io_RD_lo_lo_1,io_RD_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_124 = {_io_RD_T_122,io_rdata[47:40]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_127 = {1'h0,io_rdata[47:40]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[
    55]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55
    ],io_RD_lo_lo_lo_2}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],
    io_RD_lo_lo_lo_2,io_RD_lo_lo_2}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_185 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55]
    ,io_RD_lo_lo_lo_2,io_RD_lo_lo_2,io_RD_lo_2}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_187 = {_io_RD_T_185,io_rdata[55:48]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_190 = {1'h0,io_rdata[55:48]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[
    63]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63
    ],io_RD_lo_lo_lo_3}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_3,io_RD_lo_lo_3}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_248 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]
    ,io_RD_lo_lo_lo_3,io_RD_lo_lo_3,io_RD_lo_3}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_250 = {_io_RD_T_248,io_rdata[63:56]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_253 = {1'h0,io_rdata[63:56]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_255 = 3'h0 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_64} : _io_RD_T_61; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_257 = 3'h3 == _io_RD_T_1 ? _io_RD_T_124 : _io_RD_T_255; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_259 = 3'h2 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_127} : _io_RD_T_257; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_261 = 3'h5 == _io_RD_T_1 ? _io_RD_T_187 : _io_RD_T_259; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_263 = 3'h4 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_190} : _io_RD_T_261; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_265 = 3'h7 == _io_RD_T_1 ? _io_RD_T_250 : _io_RD_T_263; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_267 = 3'h6 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_253} : _io_RD_T_265; // @[Mux.scala 81:58]
  wire [6:0] io_RD_lo_lo_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4,io_RD_lo_lo_4}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_327 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4,io_RD_lo_lo_4,io_RD_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_329 = {_io_RD_T_327,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_332 = {1'h0,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[
    15]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15
    ],io_RD_lo_lo_lo_5}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_5,io_RD_lo_lo_5}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_390 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]
    ,io_RD_lo_lo_lo_5,io_RD_lo_lo_5,io_RD_lo_5}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_392 = {_io_RD_T_390,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_395 = {1'h0,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[
    23]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23
    ],io_RD_lo_lo_lo_6}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],
    io_RD_lo_lo_lo_6,io_RD_lo_lo_6}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_453 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23]
    ,io_RD_lo_lo_lo_6,io_RD_lo_lo_6,io_RD_lo_6}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_455 = {_io_RD_T_453,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_458 = {1'h0,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[
    31]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31
    ],io_RD_lo_lo_lo_7}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_7,io_RD_lo_lo_7}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_516 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]
    ,io_RD_lo_lo_lo_7,io_RD_lo_lo_7,io_RD_lo_7}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_518 = {_io_RD_T_516,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_521 = {1'h0,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_523 = 3'h0 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_332} : _io_RD_T_329; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_525 = 3'h3 == _io_RD_T_1 ? _io_RD_T_392 : _io_RD_T_523; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_527 = 3'h2 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_395} : _io_RD_T_525; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_529 = 3'h5 == _io_RD_T_1 ? _io_RD_T_455 : _io_RD_T_527; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_531 = 3'h4 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_458} : _io_RD_T_529; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_533 = 3'h7 == _io_RD_T_1 ? _io_RD_T_518 : _io_RD_T_531; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_535 = 3'h6 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_521} : _io_RD_T_533; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_536 = third_ra ? _io_RD_T_267 : _io_RD_T_535; // @[dmem.scala 72:19]
  wire [5:0] io_RD_lo_lo_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8,io_RD_lo_lo_8}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_590 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8,io_RD_lo_lo_8,io_RD_lo_8,io_rdata[47:32]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_593 = {1'h0,io_rdata[47:32]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9,io_RD_lo_lo_9}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_645 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9,io_RD_lo_lo_9,io_RD_lo_9,io_rdata[63:48]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_648 = {1'h0,io_rdata[63:48]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_650 = 3'h1 == _io_RD_T_1 ? _io_RD_T_590 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_652 = 3'h0 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_593} : _io_RD_T_650; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_654 = 3'h5 == _io_RD_T_1 ? _io_RD_T_645 : _io_RD_T_652; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_656 = 3'h4 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_648} : _io_RD_T_654; // @[Mux.scala 81:58]
  wire [5:0] io_RD_lo_lo_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10,io_RD_lo_lo_10}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_710 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10,io_RD_lo_lo_10,io_RD_lo_10,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_713 = {1'h0,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11,io_RD_lo_lo_11}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_765 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11,io_RD_lo_lo_11,io_RD_lo_11,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_768 = {1'h0,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_770 = 3'h1 == _io_RD_T_1 ? _io_RD_T_710 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_772 = 3'h0 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_713} : _io_RD_T_770; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_774 = 3'h5 == _io_RD_T_1 ? _io_RD_T_765 : _io_RD_T_772; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_776 = 3'h4 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_768} : _io_RD_T_774; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_777 = third_ra ? _io_RD_T_656 : _io_RD_T_776; // @[dmem.scala 73:19]
  wire [7:0] io_RD_lo_lo_12 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63
    ],io_rdata[63]}; // @[Cat.scala 31:58]
  wire [15:0] io_RD_lo_12 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_rdata[63],io_RD_lo_lo_12}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_812 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]
    ,io_rdata[63],io_RD_lo_lo_12,io_RD_lo_12}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_814 = {_io_RD_T_812,io_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [32:0] _io_RD_T_816 = {1'h0,io_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_817 = io_SIGN ? _io_RD_T_814 : {{31'd0}, _io_RD_T_816}; // @[dmem.scala 65:12]
  wire [7:0] io_RD_lo_lo_13 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31
    ],io_rdata[31]}; // @[Cat.scala 31:58]
  wire [15:0] io_RD_lo_13 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_rdata[31],io_RD_lo_lo_13}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_852 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]
    ,io_rdata[31],io_RD_lo_lo_13,io_RD_lo_13}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_854 = {_io_RD_T_852,io_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [32:0] _io_RD_T_856 = {1'h0,io_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_857 = io_SIGN ? _io_RD_T_854 : {{31'd0}, _io_RD_T_856}; // @[dmem.scala 65:12]
  wire [63:0] _io_RD_T_858 = third_ra ? _io_RD_T_817 : _io_RD_T_857; // @[dmem.scala 74:19]
  wire [63:0] _io_RD_T_860 = 2'h1 == io_WIDTH ? _io_RD_T_777 : _io_RD_T_536; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_862 = 2'h2 == io_WIDTH ? _io_RD_T_858 : _io_RD_T_860; // @[Mux.scala 81:58]
  assign io_RD = 2'h3 == io_WIDTH ? io_rdata : _io_RD_T_862; // @[Mux.scala 81:58]
  assign io_data_pending = ~io_data_ok; // @[dmem.scala 36:24]
endmodule
module ysyx_22040886_dmemreq(
  input         io_en,
  input         io_MemWriteE,
  input         io_MemToRegE,
  input  [1:0]  io_MemWidthE,
  input  [31:0] io_VAddrE,
  input  [63:0] io_WriteDataE,
  output        io_req,
  output        io_wr,
  output [1:0]  io_size,
  output [31:0] io_addr,
  output [63:0] io_wdata,
  output [7:0]  io_wstrb
);
  wire [2:0] ra = io_VAddrE[2:0]; // @[dmemreq.scala 98:23]
  wire [1:0] _io_wstrb_T_1 = 3'h1 == ra ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _io_wstrb_T_3 = 3'h2 == ra ? 3'h4 : {{1'd0}, _io_wstrb_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_5 = 3'h3 == ra ? 4'h8 : {{1'd0}, _io_wstrb_T_3}; // @[Mux.scala 81:58]
  wire [4:0] _io_wstrb_T_7 = 3'h4 == ra ? 5'h10 : {{1'd0}, _io_wstrb_T_5}; // @[Mux.scala 81:58]
  wire [5:0] _io_wstrb_T_9 = 3'h5 == ra ? 6'h20 : {{1'd0}, _io_wstrb_T_7}; // @[Mux.scala 81:58]
  wire [6:0] _io_wstrb_T_11 = 3'h6 == ra ? 7'h40 : {{1'd0}, _io_wstrb_T_9}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_13 = 3'h7 == ra ? 8'h80 : {{1'd0}, _io_wstrb_T_11}; // @[Mux.scala 81:58]
  wire [1:0] _io_wstrb_T_15 = 3'h0 == ra ? 2'h3 : 2'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_17 = 3'h2 == ra ? 4'hc : {{2'd0}, _io_wstrb_T_15}; // @[Mux.scala 81:58]
  wire [5:0] _io_wstrb_T_19 = 3'h4 == ra ? 6'h30 : {{2'd0}, _io_wstrb_T_17}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_21 = 3'h6 == ra ? 8'hc0 : {{2'd0}, _io_wstrb_T_19}; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_23 = 3'h0 == ra ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_25 = 3'h4 == ra ? 8'hf0 : {{4'd0}, _io_wstrb_T_23}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_27 = 3'h0 == ra ? 8'hff : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_29 = 2'h1 == io_MemWidthE ? _io_wstrb_T_21 : _io_wstrb_T_13; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_31 = 2'h2 == io_MemWidthE ? _io_wstrb_T_25 : _io_wstrb_T_29; // @[Mux.scala 81:58]
  wire  _io_wdata_T_1 = io_VAddrE[31:29] == 3'h4; // @[macros.scala 487:55]
  wire [8:0] _io_wdata_T_5 = {1'h0,io_WriteDataE[7:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_9 = {1'h0,io_WriteDataE[7:0],8'h0}; // @[Cat.scala 31:58]
  wire [24:0] _io_wdata_T_13 = {1'h0,io_WriteDataE[7:0],16'h0}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_17 = {1'h0,io_WriteDataE[7:0],24'h0}; // @[Cat.scala 31:58]
  wire [40:0] _io_wdata_T_21 = {1'h0,io_WriteDataE[7:0],32'h0}; // @[Cat.scala 31:58]
  wire [48:0] _io_wdata_T_25 = {1'h0,io_WriteDataE[7:0],40'h0}; // @[Cat.scala 31:58]
  wire [56:0] _io_wdata_T_29 = {1'h0,io_WriteDataE[7:0],48'h0}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_33 = {1'h0,io_WriteDataE[7:0],56'h0}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_35 = 3'h1 == ra ? _io_wdata_T_9 : {{8'd0}, _io_wdata_T_5}; // @[Mux.scala 81:58]
  wire [24:0] _io_wdata_T_37 = 3'h2 == ra ? _io_wdata_T_13 : {{8'd0}, _io_wdata_T_35}; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_39 = 3'h3 == ra ? _io_wdata_T_17 : {{8'd0}, _io_wdata_T_37}; // @[Mux.scala 81:58]
  wire [40:0] _io_wdata_T_41 = 3'h4 == ra ? _io_wdata_T_21 : {{8'd0}, _io_wdata_T_39}; // @[Mux.scala 81:58]
  wire [48:0] _io_wdata_T_43 = 3'h5 == ra ? _io_wdata_T_25 : {{8'd0}, _io_wdata_T_41}; // @[Mux.scala 81:58]
  wire [56:0] _io_wdata_T_45 = 3'h6 == ra ? _io_wdata_T_29 : {{8'd0}, _io_wdata_T_43}; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_47 = 3'h7 == ra ? _io_wdata_T_33 : {{8'd0}, _io_wdata_T_45}; // @[Mux.scala 81:58]
  wire [16:0] _io_wdata_T_50 = {1'h0,io_WriteDataE[15:0]}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_54 = {1'h0,io_WriteDataE[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [48:0] _io_wdata_T_58 = {1'h0,io_WriteDataE[15:0],32'h0}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_62 = {1'h0,io_WriteDataE[15:0],48'h0}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_64 = 3'h0 == ra ? _io_wdata_T_50 : 17'h0; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_66 = 3'h2 == ra ? _io_wdata_T_54 : {{16'd0}, _io_wdata_T_64}; // @[Mux.scala 81:58]
  wire [48:0] _io_wdata_T_68 = 3'h4 == ra ? _io_wdata_T_58 : {{16'd0}, _io_wdata_T_66}; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_70 = 3'h6 == ra ? _io_wdata_T_62 : {{16'd0}, _io_wdata_T_68}; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_73 = {1'h0,io_WriteDataE[31:0]}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_77 = {1'h0,io_WriteDataE[31:0],32'h0}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_79 = 3'h0 == ra ? _io_wdata_T_73 : 33'h0; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_81 = 3'h4 == ra ? _io_wdata_T_77 : {{32'd0}, _io_wdata_T_79}; // @[Mux.scala 81:58]
  wire [63:0] _io_wdata_T_83 = ra == 3'h0 ? io_WriteDataE : 64'h0; // @[dmemreq.scala 67:23]
  wire [64:0] _io_wdata_T_85 = 2'h1 == io_MemWidthE ? _io_wdata_T_70 : _io_wdata_T_47; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_87 = 2'h2 == io_MemWidthE ? _io_wdata_T_81 : _io_wdata_T_85; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_89 = 2'h3 == io_MemWidthE ? {{1'd0}, _io_wdata_T_83} : _io_wdata_T_87; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_90 = _io_wdata_T_1 ? _io_wdata_T_89 : {{1'd0}, io_WriteDataE}; // @[dmemreq.scala 113:23]
  assign io_req = io_en & (io_MemToRegE | io_MemWriteE); // @[dmemreq.scala 114:33]
  assign io_wr = io_MemWriteE; // @[dmemreq.scala 100:17]
  assign io_size = io_MemWidthE; // @[dmemreq.scala 110:17]
  assign io_addr = io_VAddrE; // @[dmemreq.scala 111:17]
  assign io_wdata = _io_wdata_T_90[63:0]; // @[dmemreq.scala 113:17]
  assign io_wstrb = 2'h3 == io_MemWidthE ? _io_wstrb_T_27 : _io_wstrb_T_31; // @[Mux.scala 81:58]
endmodule
module ysyx_22040886_ex2mem(
  input         clock,
  input         reset,
  input         io1_RegWriteE,
  input         io1_MemToRegE,
  input         io1_LoadUnsignedE,
  input  [1:0]  io1_MemWidthE,
  input         io1_csrWriteE,
  input  [11:0] io1_WritecsrAddrE,
  input  [63:0] io1_PCE,
  input         io1_BranchJump_JrE,
  input         io_en,
  input         io_clr,
  input  [63:0] io_WriteDataE,
  input  [4:0]  io_WriteRegE,
  input  [63:0] io_PhyAddrE,
  input  [63:0] io_CsrWritedataE,
  input  [31:0] io_ExceptionTypeE,
  output        io_RegWriteM,
  output        io_MemToRegM,
  output [63:0] io_WriteDataM,
  output [4:0]  io_WriteRegM,
  output        io_LoadUnsignedM,
  output [1:0]  io_MemWidthM,
  output [63:0] io_PhyAddrM,
  output        io_csrWriteM,
  output [11:0] io_WritecsrAddrM,
  output [63:0] io_PCM,
  output [31:0] io_ExceptionTypeM_Out,
  output        io_BranchJump_JrM,
  output [63:0] io_CsrWritedataM
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg  RegWrite_Reg; // @[ex2mem.scala 58:38]
  reg  MemToReg_Reg; // @[ex2mem.scala 59:38]
  reg [63:0] WriteData_Reg; // @[ex2mem.scala 62:39]
  reg [4:0] WriteReg_Reg; // @[ex2mem.scala 63:38]
  reg  LoadUnsigned_Reg; // @[ex2mem.scala 66:42]
  reg [1:0] MemWidth_Reg; // @[ex2mem.scala 67:38]
  reg [63:0] PhyAddr_Reg; // @[ex2mem.scala 68:37]
  reg  csrWrite_Reg; // @[ex2mem.scala 72:38]
  reg [11:0] WritecsrAddr_Reg; // @[ex2mem.scala 74:42]
  reg [63:0] PC_Reg; // @[ex2mem.scala 77:32]
  reg [31:0] ExceptionType_Reg; // @[ex2mem.scala 79:41]
  reg  BranchJump_JrM_Reg; // @[ex2mem.scala 81:43]
  reg [63:0] CsrWritedataReg; // @[ex2mem.scala 86:43]
  assign io_RegWriteM = RegWrite_Reg; // @[ex2mem.scala 122:30]
  assign io_MemToRegM = MemToReg_Reg; // @[ex2mem.scala 123:30]
  assign io_WriteDataM = WriteData_Reg; // @[ex2mem.scala 126:30]
  assign io_WriteRegM = WriteReg_Reg; // @[ex2mem.scala 127:30]
  assign io_LoadUnsignedM = LoadUnsigned_Reg; // @[ex2mem.scala 130:30]
  assign io_MemWidthM = MemWidth_Reg; // @[ex2mem.scala 131:30]
  assign io_PhyAddrM = PhyAddr_Reg; // @[ex2mem.scala 132:30]
  assign io_csrWriteM = csrWrite_Reg; // @[ex2mem.scala 135:30]
  assign io_WritecsrAddrM = WritecsrAddr_Reg; // @[ex2mem.scala 137:30]
  assign io_PCM = PC_Reg; // @[ex2mem.scala 140:30]
  assign io_ExceptionTypeM_Out = ExceptionType_Reg; // @[ex2mem.scala 142:30]
  assign io_BranchJump_JrM = BranchJump_JrM_Reg; // @[ex2mem.scala 144:30]
  assign io_CsrWritedataM = CsrWritedataReg; // @[ex2mem.scala 149:30]
  always @(posedge clock) begin
    if (reset) begin // @[ex2mem.scala 58:38]
      RegWrite_Reg <= 1'h0; // @[ex2mem.scala 58:38]
    end else if (io_clr) begin // @[ex2mem.scala 91:38]
      RegWrite_Reg <= 1'h0;
    end else if (io_en) begin // @[ex2mem.scala 91:61]
      RegWrite_Reg <= io1_RegWriteE;
    end
    if (reset) begin // @[ex2mem.scala 59:38]
      MemToReg_Reg <= 1'h0; // @[ex2mem.scala 59:38]
    end else if (io_clr) begin // @[ex2mem.scala 110:38]
      MemToReg_Reg <= 1'h0;
    end else if (io_en) begin // @[ex2mem.scala 110:61]
      MemToReg_Reg <= io1_MemToRegE;
    end
    if (reset) begin // @[ex2mem.scala 62:39]
      WriteData_Reg <= 64'h0; // @[ex2mem.scala 62:39]
    end else if (io_clr) begin // @[ex2mem.scala 94:38]
      WriteData_Reg <= 64'h0;
    end else if (io_en) begin // @[ex2mem.scala 94:61]
      WriteData_Reg <= io_WriteDataE;
    end
    if (reset) begin // @[ex2mem.scala 63:38]
      WriteReg_Reg <= 5'h0; // @[ex2mem.scala 63:38]
    end else if (io_clr) begin // @[ex2mem.scala 95:38]
      WriteReg_Reg <= 5'h0;
    end else if (io_en) begin // @[ex2mem.scala 95:61]
      WriteReg_Reg <= io_WriteRegE;
    end
    if (reset) begin // @[ex2mem.scala 66:42]
      LoadUnsigned_Reg <= 1'h0; // @[ex2mem.scala 66:42]
    end else if (io_clr) begin // @[ex2mem.scala 98:38]
      LoadUnsigned_Reg <= 1'h0;
    end else if (io_en) begin // @[ex2mem.scala 98:61]
      LoadUnsigned_Reg <= io1_LoadUnsignedE;
    end
    if (reset) begin // @[ex2mem.scala 67:38]
      MemWidth_Reg <= 2'h0; // @[ex2mem.scala 67:38]
    end else if (io_clr) begin // @[ex2mem.scala 99:38]
      MemWidth_Reg <= 2'h0;
    end else if (io_en) begin // @[ex2mem.scala 99:61]
      MemWidth_Reg <= io1_MemWidthE;
    end
    if (reset) begin // @[ex2mem.scala 68:37]
      PhyAddr_Reg <= 64'h0; // @[ex2mem.scala 68:37]
    end else if (io_clr) begin // @[ex2mem.scala 100:38]
      PhyAddr_Reg <= 64'h0;
    end else if (io_en) begin // @[ex2mem.scala 100:61]
      PhyAddr_Reg <= io_PhyAddrE;
    end
    if (reset) begin // @[ex2mem.scala 72:38]
      csrWrite_Reg <= 1'h0; // @[ex2mem.scala 72:38]
    end else if (io_clr) begin // @[ex2mem.scala 102:38]
      csrWrite_Reg <= 1'h0;
    end else if (io_en) begin // @[ex2mem.scala 102:61]
      csrWrite_Reg <= io1_csrWriteE;
    end
    if (reset) begin // @[ex2mem.scala 74:42]
      WritecsrAddr_Reg <= 12'h0; // @[ex2mem.scala 74:42]
    end else if (io_clr) begin // @[ex2mem.scala 104:38]
      WritecsrAddr_Reg <= 12'h0;
    end else if (io_en) begin // @[ex2mem.scala 104:61]
      WritecsrAddr_Reg <= io1_WritecsrAddrE;
    end
    if (reset) begin // @[ex2mem.scala 77:32]
      PC_Reg <= 64'h0; // @[ex2mem.scala 77:32]
    end else if (io_clr) begin // @[ex2mem.scala 107:38]
      PC_Reg <= 64'h0;
    end else if (io_en) begin // @[ex2mem.scala 107:61]
      PC_Reg <= io1_PCE;
    end
    if (reset) begin // @[ex2mem.scala 79:41]
      ExceptionType_Reg <= 32'h0; // @[ex2mem.scala 79:41]
    end else if (io_clr) begin // @[ex2mem.scala 109:38]
      ExceptionType_Reg <= 32'h0;
    end else if (io_en) begin // @[ex2mem.scala 109:61]
      ExceptionType_Reg <= io_ExceptionTypeE;
    end
    if (reset) begin // @[ex2mem.scala 81:43]
      BranchJump_JrM_Reg <= 1'h0; // @[ex2mem.scala 81:43]
    end else if (io_clr) begin // @[ex2mem.scala 113:38]
      BranchJump_JrM_Reg <= 1'h0;
    end else if (io_en) begin // @[ex2mem.scala 113:60]
      BranchJump_JrM_Reg <= io1_BranchJump_JrE;
    end
    if (reset) begin // @[ex2mem.scala 86:43]
      CsrWritedataReg <= 64'h0; // @[ex2mem.scala 86:43]
    end else if (io_clr) begin // @[ex2mem.scala 118:38]
      CsrWritedataReg <= 64'h0;
    end else if (io_en) begin // @[ex2mem.scala 118:60]
      CsrWritedataReg <= io_CsrWritedataE;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWrite_Reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  MemToReg_Reg = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  WriteData_Reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  WriteReg_Reg = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  LoadUnsigned_Reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  MemWidth_Reg = _RAND_5[1:0];
  _RAND_6 = {2{`RANDOM}};
  PhyAddr_Reg = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  csrWrite_Reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  WritecsrAddr_Reg = _RAND_8[11:0];
  _RAND_9 = {2{`RANDOM}};
  PC_Reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  ExceptionType_Reg = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  BranchJump_JrM_Reg = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  CsrWritedataReg = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_id2ex(
  input         clock,
  input         reset,
  input         io1_RegWriteD,
  input         io1_MemToRegD,
  input         io1_MemWriteD,
  input  [15:0] io1_ALUCtrlD,
  input         io1_ALUSrcD_0,
  input         io1_ALUSrcD_1,
  input  [4:0]  io1_RegDstD,
  input         io1_LinkD,
  input         io1_csrWriteD,
  input         io1_csrToRegD,
  input         io1_LoadUnsignedD,
  input  [1:0]  io1_MemWidthD,
  input         io1_data_wD,
  input  [23:0] io1_muldiv_control,
  input         io1_muldiv_cal,
  input         io1_alu_cal,
  input  [2:0]  io1_csr_control,
  input         io1_csr_Imm,
  input         io1_fence_i_control,
  output        io2_RegWriteE,
  output        io2_MemToRegE,
  output        io2_MemWriteE,
  output [15:0] io2_ALUCtrlE,
  output        io2_ALUSrcE_0,
  output        io2_ALUSrcE_1,
  output [4:0]  io2_RegDstE,
  output        io2_LinkE,
  output [63:0] io2_PCPlus4E,
  output        io2_LoadUnsignedE,
  output [1:0]  io2_MemWidthE,
  output        io2_csrWriteE,
  output [11:0] io2_WritecsrAddrE,
  output [11:0] io2_ReadcsrAddrE,
  output [63:0] io2_PCE,
  output        io2_BranchJump_JrE,
  input         io_en,
  input         io_clr,
  output        io_csrToRegE_Out,
  input  [63:0] io_RD1D,
  input  [63:0] io_RD2D,
  input  [4:0]  io_R2D,
  input  [4:0]  io_R1D,
  input  [63:0] io_ImmD,
  input  [63:0] io_PCPlus4D,
  input  [11:0] io_WritecsrAddrD,
  input  [11:0] io_ReadcsrAddrD,
  input  [63:0] io_PCD,
  input  [31:0] io_ExceptionTypeD,
  input         io_BranchJump_JrD,
  output [63:0] io_RD1E,
  output [63:0] io_RD2E,
  output [4:0]  io_R2E,
  output [4:0]  io_R1E,
  output [63:0] io_ImmE,
  output        io_data_wE,
  output [23:0] io_muldiv_control,
  output        io_alu_calE,
  output        io_muldiv_calE,
  output [31:0] io_ExceptionTypeE_Out,
  output [2:0]  io_csr_controlE,
  output        io_csr_ImmE,
  output        io_fence_i_controlE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] RD1E_Reg; // @[id2ex.scala 99:30]
  reg [63:0] RD2E_Reg; // @[id2ex.scala 100:30]
  reg [4:0] R2E_Reg; // @[id2ex.scala 101:29]
  reg [4:0] R1E_Reg; // @[id2ex.scala 102:29]
  reg [63:0] ImmE_Reg; // @[id2ex.scala 104:30]
  reg [63:0] PCPlus4E_Reg; // @[id2ex.scala 106:34]
  reg [11:0] WritecsrAddrE_Reg; // @[id2ex.scala 112:39]
  reg [11:0] ReadcsrAddrE_Reg; // @[id2ex.scala 113:38]
  reg [63:0] PCE_Reg; // @[id2ex.scala 114:29]
  reg [31:0] ExceptionTypeE_Reg; // @[id2ex.scala 115:40]
  reg  BranchJump_JrE_Reg; // @[id2ex.scala 117:40]
  reg  decoder_port_reg_RegWriteD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_MemToRegD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_MemWriteD; // @[id2ex.scala 126:38]
  reg [15:0] decoder_port_reg_ALUCtrlD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_ALUSrcD_0; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_ALUSrcD_1; // @[id2ex.scala 126:38]
  reg [4:0] decoder_port_reg_RegDstD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_LinkD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_csrWriteD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_csrToRegD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_LoadUnsignedD; // @[id2ex.scala 126:38]
  reg [1:0] decoder_port_reg_MemWidthD; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_data_wD; // @[id2ex.scala 126:38]
  reg [23:0] decoder_port_reg_muldiv_control; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_muldiv_cal; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_alu_cal; // @[id2ex.scala 126:38]
  reg [2:0] decoder_port_reg_csr_control; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_csr_Imm; // @[id2ex.scala 126:38]
  reg  decoder_port_reg_fence_i_control; // @[id2ex.scala 126:38]
  assign io2_RegWriteE = decoder_port_reg_RegWriteD; // @[id2ex.scala 150:23]
  assign io2_MemToRegE = decoder_port_reg_MemToRegD; // @[id2ex.scala 151:23]
  assign io2_MemWriteE = decoder_port_reg_MemWriteD; // @[id2ex.scala 152:23]
  assign io2_ALUCtrlE = decoder_port_reg_ALUCtrlD; // @[id2ex.scala 153:23]
  assign io2_ALUSrcE_0 = decoder_port_reg_ALUSrcD_0; // @[id2ex.scala 154:23]
  assign io2_ALUSrcE_1 = decoder_port_reg_ALUSrcD_1; // @[id2ex.scala 154:23]
  assign io2_RegDstE = decoder_port_reg_RegDstD; // @[id2ex.scala 155:23]
  assign io2_LinkE = decoder_port_reg_LinkD; // @[id2ex.scala 162:23]
  assign io2_PCPlus4E = PCPlus4E_Reg; // @[id2ex.scala 163:23]
  assign io2_LoadUnsignedE = decoder_port_reg_LoadUnsignedD; // @[id2ex.scala 164:23]
  assign io2_MemWidthE = decoder_port_reg_MemWidthD; // @[id2ex.scala 165:23]
  assign io2_csrWriteE = decoder_port_reg_csrWriteD; // @[id2ex.scala 166:23]
  assign io2_WritecsrAddrE = WritecsrAddrE_Reg; // @[id2ex.scala 168:23]
  assign io2_ReadcsrAddrE = ReadcsrAddrE_Reg; // @[id2ex.scala 169:23]
  assign io2_PCE = PCE_Reg; // @[id2ex.scala 170:23]
  assign io2_BranchJump_JrE = BranchJump_JrE_Reg; // @[id2ex.scala 173:24]
  assign io_csrToRegE_Out = decoder_port_reg_csrToRegD; // @[id2ex.scala 167:26]
  assign io_RD1E = RD1E_Reg; // @[id2ex.scala 156:23]
  assign io_RD2E = RD2E_Reg; // @[id2ex.scala 157:23]
  assign io_R2E = R2E_Reg; // @[id2ex.scala 158:23]
  assign io_R1E = R1E_Reg; // @[id2ex.scala 159:23]
  assign io_ImmE = ImmE_Reg; // @[id2ex.scala 161:23]
  assign io_data_wE = decoder_port_reg_data_wD; // @[id2ex.scala 177:27]
  assign io_muldiv_control = decoder_port_reg_muldiv_control; // @[id2ex.scala 181:27]
  assign io_alu_calE = decoder_port_reg_alu_cal; // @[id2ex.scala 149:23]
  assign io_muldiv_calE = decoder_port_reg_muldiv_cal; // @[id2ex.scala 148:23]
  assign io_ExceptionTypeE_Out = ExceptionTypeE_Reg; // @[id2ex.scala 172:26]
  assign io_csr_controlE = decoder_port_reg_csr_control; // @[id2ex.scala 183:27]
  assign io_csr_ImmE = decoder_port_reg_csr_Imm; // @[id2ex.scala 184:27]
  assign io_fence_i_controlE = decoder_port_reg_fence_i_control; // @[id2ex.scala 179:27]
  always @(posedge clock) begin
    if (reset) begin // @[id2ex.scala 99:30]
      RD1E_Reg <= 64'h0; // @[id2ex.scala 99:30]
    end else if (io_clr) begin // @[id2ex.scala 129:42]
      RD1E_Reg <= 64'h0;
    end else if (io_en) begin // @[id2ex.scala 129:64]
      RD1E_Reg <= io_RD1D;
    end
    if (reset) begin // @[id2ex.scala 100:30]
      RD2E_Reg <= 64'h0; // @[id2ex.scala 100:30]
    end else if (io_clr) begin // @[id2ex.scala 130:42]
      RD2E_Reg <= 64'h0;
    end else if (io_en) begin // @[id2ex.scala 130:64]
      RD2E_Reg <= io_RD2D;
    end
    if (reset) begin // @[id2ex.scala 101:29]
      R2E_Reg <= 5'h0; // @[id2ex.scala 101:29]
    end else if (io_clr) begin // @[id2ex.scala 131:42]
      R2E_Reg <= 5'h0;
    end else if (io_en) begin // @[id2ex.scala 131:64]
      R2E_Reg <= io_R2D;
    end
    if (reset) begin // @[id2ex.scala 102:29]
      R1E_Reg <= 5'h0; // @[id2ex.scala 102:29]
    end else if (io_clr) begin // @[id2ex.scala 132:42]
      R1E_Reg <= 5'h0;
    end else if (io_en) begin // @[id2ex.scala 132:64]
      R1E_Reg <= io_R1D;
    end
    if (reset) begin // @[id2ex.scala 104:30]
      ImmE_Reg <= 64'h0; // @[id2ex.scala 104:30]
    end else if (io_clr) begin // @[id2ex.scala 134:42]
      ImmE_Reg <= 64'h0;
    end else if (io_en) begin // @[id2ex.scala 134:64]
      ImmE_Reg <= io_ImmD;
    end
    if (reset) begin // @[id2ex.scala 106:34]
      PCPlus4E_Reg <= 64'h0; // @[id2ex.scala 106:34]
    end else if (io_clr) begin // @[id2ex.scala 135:42]
      PCPlus4E_Reg <= 64'h0;
    end else if (io_en) begin // @[id2ex.scala 135:64]
      PCPlus4E_Reg <= io_PCPlus4D;
    end
    if (reset) begin // @[id2ex.scala 112:39]
      WritecsrAddrE_Reg <= 12'h0; // @[id2ex.scala 112:39]
    end else if (io_clr) begin // @[id2ex.scala 136:42]
      WritecsrAddrE_Reg <= 12'h0;
    end else if (io_en) begin // @[id2ex.scala 136:64]
      WritecsrAddrE_Reg <= io_WritecsrAddrD;
    end
    if (reset) begin // @[id2ex.scala 113:38]
      ReadcsrAddrE_Reg <= 12'h0; // @[id2ex.scala 113:38]
    end else if (io_clr) begin // @[id2ex.scala 138:42]
      ReadcsrAddrE_Reg <= 12'h0;
    end else if (io_en) begin // @[id2ex.scala 138:64]
      ReadcsrAddrE_Reg <= io_ReadcsrAddrD;
    end
    if (reset) begin // @[id2ex.scala 114:29]
      PCE_Reg <= 64'h0; // @[id2ex.scala 114:29]
    end else if (io_clr) begin // @[id2ex.scala 140:42]
      PCE_Reg <= 64'h0;
    end else if (io_en) begin // @[id2ex.scala 140:64]
      PCE_Reg <= io_PCD;
    end
    if (reset) begin // @[id2ex.scala 115:40]
      ExceptionTypeE_Reg <= 32'h0; // @[id2ex.scala 115:40]
    end else if (io_clr) begin // @[id2ex.scala 141:42]
      ExceptionTypeE_Reg <= 32'h0;
    end else if (io_en) begin // @[id2ex.scala 141:64]
      ExceptionTypeE_Reg <= io_ExceptionTypeD;
    end
    if (reset) begin // @[id2ex.scala 117:40]
      BranchJump_JrE_Reg <= 1'h0; // @[id2ex.scala 117:40]
    end else if (io_clr) begin // @[id2ex.scala 142:42]
      BranchJump_JrE_Reg <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 142:64]
      BranchJump_JrE_Reg <= io_BranchJump_JrD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_RegWriteD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_RegWriteD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_RegWriteD <= io1_RegWriteD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_MemToRegD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_MemToRegD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_MemToRegD <= io1_MemToRegD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_MemWriteD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_MemWriteD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_MemWriteD <= io1_MemWriteD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_ALUCtrlD <= 16'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_ALUCtrlD <= 16'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_ALUCtrlD <= io1_ALUCtrlD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_ALUSrcD_0 <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_ALUSrcD_0 <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_ALUSrcD_0 <= io1_ALUSrcD_0;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_ALUSrcD_1 <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_ALUSrcD_1 <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_ALUSrcD_1 <= io1_ALUSrcD_1;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_RegDstD <= 5'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_RegDstD <= 5'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_RegDstD <= io1_RegDstD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_LinkD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_LinkD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_LinkD <= io1_LinkD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_csrWriteD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_csrWriteD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_csrWriteD <= io1_csrWriteD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_csrToRegD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_csrToRegD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_csrToRegD <= io1_csrToRegD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_LoadUnsignedD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_LoadUnsignedD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_LoadUnsignedD <= io1_LoadUnsignedD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_MemWidthD <= 2'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_MemWidthD <= 2'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_MemWidthD <= io1_MemWidthD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_data_wD <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_data_wD <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_data_wD <= io1_data_wD;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_muldiv_control <= 24'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_muldiv_control <= 24'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_muldiv_control <= io1_muldiv_control;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_muldiv_cal <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_muldiv_cal <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_muldiv_cal <= io1_muldiv_cal;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_alu_cal <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_alu_cal <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_alu_cal <= io1_alu_cal;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_csr_control <= 3'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_csr_control <= 3'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_csr_control <= io1_csr_control;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_csr_Imm <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_csr_Imm <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_csr_Imm <= io1_csr_Imm;
    end
    if (reset) begin // @[id2ex.scala 126:38]
      decoder_port_reg_fence_i_control <= 1'h0; // @[id2ex.scala 126:38]
    end else if (io_clr) begin // @[id2ex.scala 127:28]
      decoder_port_reg_fence_i_control <= 1'h0;
    end else if (io_en) begin // @[id2ex.scala 127:77]
      decoder_port_reg_fence_i_control <= io1_fence_i_control;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  RD1E_Reg = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  RD2E_Reg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  R2E_Reg = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  R1E_Reg = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  ImmE_Reg = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  PCPlus4E_Reg = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  WritecsrAddrE_Reg = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  ReadcsrAddrE_Reg = _RAND_7[11:0];
  _RAND_8 = {2{`RANDOM}};
  PCE_Reg = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  ExceptionTypeE_Reg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  BranchJump_JrE_Reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  decoder_port_reg_RegWriteD = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  decoder_port_reg_MemToRegD = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  decoder_port_reg_MemWriteD = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  decoder_port_reg_ALUCtrlD = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  decoder_port_reg_ALUSrcD_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  decoder_port_reg_ALUSrcD_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  decoder_port_reg_RegDstD = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  decoder_port_reg_LinkD = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  decoder_port_reg_csrWriteD = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  decoder_port_reg_csrToRegD = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  decoder_port_reg_LoadUnsignedD = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  decoder_port_reg_MemWidthD = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  decoder_port_reg_data_wD = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  decoder_port_reg_muldiv_control = _RAND_24[23:0];
  _RAND_25 = {1{`RANDOM}};
  decoder_port_reg_muldiv_cal = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  decoder_port_reg_alu_cal = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  decoder_port_reg_csr_control = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  decoder_port_reg_csr_Imm = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  decoder_port_reg_fence_i_control = _RAND_29[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_if2id(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input  [31:0] io_InstrF,
  input  [63:0] io_PCPlus4F,
  input  [63:0] io_PCF,
  input  [1:0]  io_ExceptionTypeF,
  output [31:0] io_InstrD,
  output [63:0] io_PCPlus4D,
  output [63:0] io_PCD,
  output [1:0]  io_ExceptionTypeD_Out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] InstrD_Reg; // @[if2id.scala 30:29]
  reg [63:0] PCPlus4D_Reg; // @[if2id.scala 31:31]
  reg [63:0] PCD_Reg; // @[if2id.scala 33:26]
  reg [1:0] ExceptionTypeD_Reg; // @[if2id.scala 34:37]
  assign io_InstrD = InstrD_Reg; // @[if2id.scala 38:15]
  assign io_PCPlus4D = PCPlus4D_Reg; // @[if2id.scala 39:17]
  assign io_PCD = PCD_Reg; // @[if2id.scala 42:13]
  assign io_ExceptionTypeD_Out = ExceptionTypeD_Reg; // @[if2id.scala 41:27]
  always @(posedge clock) begin
    if (reset) begin // @[if2id.scala 30:29]
      InstrD_Reg <= 32'h13; // @[if2id.scala 30:29]
    end else if (io_clr) begin // @[if2id.scala 45:35]
      InstrD_Reg <= 32'h0;
    end else if (io_en) begin // @[if2id.scala 45:57]
      InstrD_Reg <= io_InstrF;
    end
    if (reset) begin // @[if2id.scala 31:31]
      PCPlus4D_Reg <= 64'h0; // @[if2id.scala 31:31]
    end else if (io_clr) begin // @[if2id.scala 46:35]
      PCPlus4D_Reg <= 64'h0;
    end else if (io_en) begin // @[if2id.scala 46:57]
      PCPlus4D_Reg <= io_PCPlus4F;
    end
    if (reset) begin // @[if2id.scala 33:26]
      PCD_Reg <= 64'h0; // @[if2id.scala 33:26]
    end else if (io_clr) begin // @[if2id.scala 48:39]
      PCD_Reg <= 64'h0;
    end else if (io_en) begin // @[if2id.scala 48:61]
      PCD_Reg <= io_PCF;
    end
    if (reset) begin // @[if2id.scala 34:37]
      ExceptionTypeD_Reg <= 2'h0; // @[if2id.scala 34:37]
    end else if (io_clr) begin // @[if2id.scala 49:39]
      ExceptionTypeD_Reg <= 2'h0;
    end else if (io_en) begin // @[if2id.scala 49:61]
      ExceptionTypeD_Reg <= io_ExceptionTypeF;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InstrD_Reg = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  PCPlus4D_Reg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  PCD_Reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  ExceptionTypeD_Reg = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_mem2wb(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input         io_RegWriteM,
  input  [63:0] io_ResultM,
  input  [4:0]  io_WriteRegM,
  input         io_csrWriteM,
  input  [11:0] io_WritecsrAddrM,
  input  [63:0] io_CsrWritedataM,
  input  [63:0] io_PCM,
  input  [30:0] io_ExceptionTypeM,
  input         io_BranchJump_JrM,
  output        io_RegWriteW_Out,
  output [63:0] io_ResultW,
  output [4:0]  io_WriteRegW,
  output        io_csrWriteW,
  output [11:0] io_WritecsrAddrW,
  output [63:0] io_PCW,
  output [30:0] io_ExceptionTypeW_Out,
  output        io_BranchJump_JrW,
  output [63:0] io_CsrWritedataW
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  RegWriteW; // @[mem2wb.scala 51:34]
  reg [63:0] ResultW; // @[mem2wb.scala 54:32]
  reg [4:0] WriteRegW; // @[mem2wb.scala 55:34]
  reg  csrWriteW; // @[mem2wb.scala 57:34]
  reg [11:0] WritecsrAddrW; // @[mem2wb.scala 58:38]
  reg [63:0] PCW; // @[mem2wb.scala 60:28]
  reg [30:0] ExceptionTypeW; // @[mem2wb.scala 62:39]
  reg  BranchJump_JrW_Reg; // @[mem2wb.scala 64:43]
  reg [63:0] CsrWritedataReg; // @[mem2wb.scala 69:40]
  assign io_RegWriteW_Out = RegWriteW; // @[mem2wb.scala 71:36]
  assign io_ResultW = ResultW; // @[mem2wb.scala 74:32]
  assign io_WriteRegW = WriteRegW; // @[mem2wb.scala 75:32]
  assign io_csrWriteW = csrWriteW; // @[mem2wb.scala 76:32]
  assign io_WritecsrAddrW = WritecsrAddrW; // @[mem2wb.scala 77:32]
  assign io_PCW = PCW; // @[mem2wb.scala 79:32]
  assign io_ExceptionTypeW_Out = ExceptionTypeW; // @[mem2wb.scala 81:32]
  assign io_BranchJump_JrW = BranchJump_JrW_Reg; // @[mem2wb.scala 82:32]
  assign io_CsrWritedataW = CsrWritedataReg; // @[mem2wb.scala 108:28]
  always @(posedge clock) begin
    if (reset) begin // @[mem2wb.scala 51:34]
      RegWriteW <= 1'h0; // @[mem2wb.scala 51:34]
    end else if (io_clr) begin // @[mem2wb.scala 88:34]
      RegWriteW <= 1'h0;
    end else if (io_en) begin // @[mem2wb.scala 88:56]
      RegWriteW <= io_RegWriteM;
    end
    if (reset) begin // @[mem2wb.scala 54:32]
      ResultW <= 64'h0; // @[mem2wb.scala 54:32]
    end else if (io_clr) begin // @[mem2wb.scala 91:34]
      ResultW <= 64'h0;
    end else if (io_en) begin // @[mem2wb.scala 91:56]
      ResultW <= io_ResultM;
    end
    if (reset) begin // @[mem2wb.scala 55:34]
      WriteRegW <= 5'h0; // @[mem2wb.scala 55:34]
    end else if (io_clr) begin // @[mem2wb.scala 92:34]
      WriteRegW <= 5'h0;
    end else if (io_en) begin // @[mem2wb.scala 92:56]
      WriteRegW <= io_WriteRegM;
    end
    if (reset) begin // @[mem2wb.scala 57:34]
      csrWriteW <= 1'h0; // @[mem2wb.scala 57:34]
    end else if (io_clr) begin // @[mem2wb.scala 95:34]
      csrWriteW <= 1'h0;
    end else if (io_en) begin // @[mem2wb.scala 95:56]
      csrWriteW <= io_csrWriteM;
    end
    if (reset) begin // @[mem2wb.scala 58:38]
      WritecsrAddrW <= 12'h0; // @[mem2wb.scala 58:38]
    end else if (io_clr) begin // @[mem2wb.scala 96:34]
      WritecsrAddrW <= 12'h0;
    end else if (io_en) begin // @[mem2wb.scala 96:56]
      WritecsrAddrW <= io_WritecsrAddrM;
    end
    if (reset) begin // @[mem2wb.scala 60:28]
      PCW <= 64'h0; // @[mem2wb.scala 60:28]
    end else if (io_clr) begin // @[mem2wb.scala 98:34]
      PCW <= 64'h0;
    end else if (io_en) begin // @[mem2wb.scala 98:56]
      PCW <= io_PCM;
    end
    if (reset) begin // @[mem2wb.scala 62:39]
      ExceptionTypeW <= 31'h0; // @[mem2wb.scala 62:39]
    end else if (io_clr) begin // @[mem2wb.scala 100:34]
      ExceptionTypeW <= 31'h0;
    end else if (io_en) begin // @[mem2wb.scala 100:56]
      ExceptionTypeW <= io_ExceptionTypeM;
    end
    if (reset) begin // @[mem2wb.scala 64:43]
      BranchJump_JrW_Reg <= 1'h0; // @[mem2wb.scala 64:43]
    end else if (io_clr) begin // @[mem2wb.scala 101:49]
      BranchJump_JrW_Reg <= 1'h0;
    end else if (io_en) begin // @[mem2wb.scala 101:71]
      BranchJump_JrW_Reg <= io_BranchJump_JrM;
    end
    if (reset) begin // @[mem2wb.scala 69:40]
      CsrWritedataReg <= 64'h0; // @[mem2wb.scala 69:40]
    end else if (io_clr) begin // @[mem2wb.scala 107:34]
      CsrWritedataReg <= 64'h0;
    end else if (io_en) begin // @[mem2wb.scala 107:56]
      CsrWritedataReg <= io_CsrWritedataM;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWriteW = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ResultW = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  WriteRegW = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  csrWriteW = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  WritecsrAddrW = _RAND_4[11:0];
  _RAND_5 = {2{`RANDOM}};
  PCW = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  ExceptionTypeW = _RAND_6[30:0];
  _RAND_7 = {1{`RANDOM}};
  BranchJump_JrW_Reg = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  CsrWritedataReg = _RAND_8[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_addr_cal(
  input  [31:0] io_d_vaddr,
  output [31:0] io_d_paddr,
  output        io_d_cached
);
  assign io_d_paddr = io_d_vaddr; // @[addr_cal.scala 24:16]
  assign io_d_cached = io_d_vaddr[31:29] == 3'h4; // @[macros.scala 487:55]
endmodule
module ysyx_22040886_csa(
  input  [131:0] io_data_0,
  input  [131:0] io_data_1,
  input  [131:0] io_data_2,
  output [131:0] io_result_0,
  output [131:0] io_result_1
);
  wire [131:0] _io_result_0_T = io_data_0 ^ io_data_1; // @[hard_cal.scala 187:32]
  wire [131:0] _io_result_1_T = io_data_0 & io_data_1; // @[hard_cal.scala 188:37]
  wire [131:0] _io_result_1_T_1 = io_data_1 & io_data_2; // @[hard_cal.scala 188:65]
  wire [131:0] _io_result_1_T_2 = _io_result_1_T | _io_result_1_T_1; // @[hard_cal.scala 188:51]
  wire [131:0] _io_result_1_T_3 = io_data_2 & io_data_0; // @[hard_cal.scala 188:93]
  wire [131:0] _io_result_1_T_4 = _io_result_1_T_2 | _io_result_1_T_3; // @[hard_cal.scala 188:79]
  wire [132:0] _io_result_1_T_5 = {_io_result_1_T_4,1'h0}; // @[Cat.scala 31:58]
  assign io_result_0 = _io_result_0_T ^ io_data_2; // @[hard_cal.scala 187:45]
  assign io_result_1 = _io_result_1_T_5[131:0]; // @[hard_cal.scala 188:18]
endmodule
module ysyx_22040886_wallace_adder(
  input          clock,
  input          reset,
  input  [131:0] io_data_in_0,
  input  [131:0] io_data_in_1,
  input  [131:0] io_data_in_2,
  input  [131:0] io_data_in_3,
  input  [131:0] io_data_in_4,
  input  [131:0] io_data_in_5,
  input  [131:0] io_data_in_6,
  input  [131:0] io_data_in_7,
  input  [131:0] io_data_in_8,
  input  [131:0] io_data_in_9,
  input  [131:0] io_data_in_10,
  input  [131:0] io_data_in_11,
  input  [131:0] io_data_in_12,
  input  [131:0] io_data_in_13,
  input  [131:0] io_data_in_14,
  input  [131:0] io_data_in_15,
  input  [131:0] io_data_in_16,
  input  [131:0] io_data_in_17,
  input  [131:0] io_data_in_18,
  input  [131:0] io_data_in_19,
  input  [131:0] io_data_in_20,
  input  [131:0] io_data_in_21,
  input  [131:0] io_data_in_22,
  input  [131:0] io_data_in_23,
  input  [131:0] io_data_in_24,
  input  [131:0] io_data_in_25,
  input  [131:0] io_data_in_26,
  input  [131:0] io_data_in_27,
  input  [131:0] io_data_in_28,
  input  [131:0] io_data_in_29,
  input  [131:0] io_data_in_30,
  input  [131:0] io_data_in_31,
  input  [131:0] io_data_in_32,
  output [131:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
  reg [159:0] _RAND_6;
  reg [159:0] _RAND_7;
  reg [159:0] _RAND_8;
  reg [159:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [159:0] _RAND_11;
  reg [159:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [159:0] _RAND_14;
  reg [159:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [159:0] _RAND_17;
  reg [159:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [159:0] _RAND_20;
  reg [159:0] _RAND_21;
  reg [159:0] _RAND_22;
  reg [159:0] _RAND_23;
  reg [159:0] _RAND_24;
  reg [159:0] _RAND_25;
  reg [159:0] _RAND_26;
  reg [159:0] _RAND_27;
  reg [159:0] _RAND_28;
  reg [159:0] _RAND_29;
  reg [159:0] _RAND_30;
  reg [159:0] _RAND_31;
  reg [159:0] _RAND_32;
  reg [159:0] _RAND_33;
  reg [159:0] _RAND_34;
  reg [159:0] _RAND_35;
  reg [159:0] _RAND_36;
  reg [159:0] _RAND_37;
  reg [159:0] _RAND_38;
  reg [159:0] _RAND_39;
  reg [159:0] _RAND_40;
  reg [159:0] _RAND_41;
  reg [159:0] _RAND_42;
  reg [159:0] _RAND_43;
  reg [159:0] _RAND_44;
  reg [159:0] _RAND_45;
  reg [159:0] _RAND_46;
  reg [159:0] _RAND_47;
  reg [159:0] _RAND_48;
  reg [159:0] _RAND_49;
  reg [159:0] _RAND_50;
  reg [159:0] _RAND_51;
  reg [159:0] _RAND_52;
  reg [159:0] _RAND_53;
  reg [159:0] _RAND_54;
  reg [159:0] _RAND_55;
  reg [159:0] _RAND_56;
  reg [159:0] _RAND_57;
  reg [159:0] _RAND_58;
  reg [159:0] _RAND_59;
  reg [159:0] _RAND_60;
  reg [159:0] _RAND_61;
  reg [159:0] _RAND_62;
  reg [159:0] _RAND_63;
  reg [159:0] _RAND_64;
  reg [159:0] _RAND_65;
  reg [159:0] _RAND_66;
  reg [159:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [131:0] csa_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_1_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_1_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_1_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_1_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_1_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_2_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_2_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_2_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_2_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_2_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_3_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_3_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_3_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_3_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_3_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_4_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_4_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_4_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_4_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_4_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_5_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_5_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_5_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_5_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_5_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_6_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_6_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_6_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_6_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_6_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_7_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_7_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_7_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_7_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_7_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_8_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_8_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_8_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_8_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_8_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_9_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_9_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_9_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_9_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_9_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_10_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_10_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_10_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_10_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_10_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_11_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_11_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_11_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_11_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_11_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_12_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_12_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_12_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_12_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_12_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_13_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_13_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_13_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_13_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_13_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_14_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_14_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_14_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_14_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_14_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_15_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_15_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_15_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_15_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_15_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_16_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_16_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_16_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_16_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_16_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_17_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_17_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_17_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_17_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_17_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_18_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_18_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_18_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_18_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_18_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_19_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_19_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_19_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_19_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_19_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_20_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_20_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_20_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_20_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_20_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_21_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_21_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_21_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_21_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_21_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_22_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_22_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_22_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_22_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_22_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_23_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_23_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_23_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_23_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_23_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_24_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_24_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_24_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_24_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_24_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_25_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_25_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_25_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_25_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_25_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_26_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_26_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_26_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_26_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_26_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_27_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_27_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_27_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_27_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_27_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_28_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_28_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_28_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_28_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_28_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_29_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_29_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_29_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_29_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_29_io_result_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_30_io_data_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_30_io_data_1; // @[hard_cal.scala 209:61]
  wire [131:0] csa_30_io_data_2; // @[hard_cal.scala 209:61]
  wire [131:0] csa_30_io_result_0; // @[hard_cal.scala 209:61]
  wire [131:0] csa_30_io_result_1; // @[hard_cal.scala 209:61]
  reg [131:0] vec_data_out_data_reg__0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__4; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__5; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__6; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__7; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__8; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__9; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__10; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__11; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__12; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__13; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__14; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__15; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__16; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__17; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__18; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__19; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__20; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg__21; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_4; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_5; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_6; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_7; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_8; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_9; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_10; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_11; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_12; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_13; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_1_14; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_4; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_5; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_6; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_7; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_8; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_2_9; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_4; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_5; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_3_6; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_4_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_4_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_4_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_4_3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_4_4; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_5_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_5_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_5_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_5_3; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_6_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_6_1; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_out_data_reg_6_2; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_0; // @[hard_cal.scala 225:39]
  reg [131:0] vec_data_1; // @[hard_cal.scala 225:39]
  wire [131:0] vec_data_csa_adder__0_result_0 = csa_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__0_result_1 = csa_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__1_result_0 = csa_1_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__1_result_1 = csa_1_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__2_result_0 = csa_2_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__2_result_1 = csa_2_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__3_result_0 = csa_3_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__3_result_1 = csa_3_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__4_result_0 = csa_4_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__4_result_1 = csa_4_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__5_result_0 = csa_5_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__5_result_1 = csa_5_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__6_result_0 = csa_6_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__6_result_1 = csa_6_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__7_result_0 = csa_7_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__7_result_1 = csa_7_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__8_result_0 = csa_8_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__8_result_1 = csa_8_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__9_result_0 = csa_9_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__9_result_1 = csa_9_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__10_result_0 = csa_10_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder__10_result_1 = csa_10_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_0_result_0 = csa_11_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_0_result_1 = csa_11_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_1_result_0 = csa_12_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_1_result_1 = csa_12_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_2_result_0 = csa_13_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_2_result_1 = csa_13_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_3_result_0 = csa_14_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_3_result_1 = csa_14_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_4_result_0 = csa_15_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_4_result_1 = csa_15_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_5_result_0 = csa_16_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_5_result_1 = csa_16_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_6_result_0 = csa_17_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_1_6_result_1 = csa_17_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_0_result_0 = csa_18_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_0_result_1 = csa_18_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_1_result_0 = csa_19_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_1_result_1 = csa_19_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_2_result_0 = csa_20_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_2_result_1 = csa_20_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_3_result_0 = csa_21_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_3_result_1 = csa_21_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_4_result_0 = csa_22_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_2_4_result_1 = csa_22_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_0_result_0 = csa_23_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_0_result_1 = csa_23_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_1_result_0 = csa_24_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_1_result_1 = csa_24_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_2_result_0 = csa_25_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_3_2_result_1 = csa_25_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_4_0_result_0 = csa_26_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_4_0_result_1 = csa_26_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_4_1_result_0 = csa_27_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_4_1_result_1 = csa_27_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_5_0_result_0 = csa_28_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_5_0_result_1 = csa_28_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_6_0_result_0 = csa_29_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_6_0_result_1 = csa_29_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_7_0_result_0 = csa_30_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [131:0] vec_data_csa_adder_7_0_result_1 = csa_30_io_result_1; // @[hard_cal.scala 209:{36,36}]
  ysyx_22040886_csa csa ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_io_data_0),
    .io_data_1(csa_io_data_1),
    .io_data_2(csa_io_data_2),
    .io_result_0(csa_io_result_0),
    .io_result_1(csa_io_result_1)
  );
  ysyx_22040886_csa csa_1 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_1_io_data_0),
    .io_data_1(csa_1_io_data_1),
    .io_data_2(csa_1_io_data_2),
    .io_result_0(csa_1_io_result_0),
    .io_result_1(csa_1_io_result_1)
  );
  ysyx_22040886_csa csa_2 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_2_io_data_0),
    .io_data_1(csa_2_io_data_1),
    .io_data_2(csa_2_io_data_2),
    .io_result_0(csa_2_io_result_0),
    .io_result_1(csa_2_io_result_1)
  );
  ysyx_22040886_csa csa_3 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_3_io_data_0),
    .io_data_1(csa_3_io_data_1),
    .io_data_2(csa_3_io_data_2),
    .io_result_0(csa_3_io_result_0),
    .io_result_1(csa_3_io_result_1)
  );
  ysyx_22040886_csa csa_4 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_4_io_data_0),
    .io_data_1(csa_4_io_data_1),
    .io_data_2(csa_4_io_data_2),
    .io_result_0(csa_4_io_result_0),
    .io_result_1(csa_4_io_result_1)
  );
  ysyx_22040886_csa csa_5 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_5_io_data_0),
    .io_data_1(csa_5_io_data_1),
    .io_data_2(csa_5_io_data_2),
    .io_result_0(csa_5_io_result_0),
    .io_result_1(csa_5_io_result_1)
  );
  ysyx_22040886_csa csa_6 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_6_io_data_0),
    .io_data_1(csa_6_io_data_1),
    .io_data_2(csa_6_io_data_2),
    .io_result_0(csa_6_io_result_0),
    .io_result_1(csa_6_io_result_1)
  );
  ysyx_22040886_csa csa_7 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_7_io_data_0),
    .io_data_1(csa_7_io_data_1),
    .io_data_2(csa_7_io_data_2),
    .io_result_0(csa_7_io_result_0),
    .io_result_1(csa_7_io_result_1)
  );
  ysyx_22040886_csa csa_8 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_8_io_data_0),
    .io_data_1(csa_8_io_data_1),
    .io_data_2(csa_8_io_data_2),
    .io_result_0(csa_8_io_result_0),
    .io_result_1(csa_8_io_result_1)
  );
  ysyx_22040886_csa csa_9 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_9_io_data_0),
    .io_data_1(csa_9_io_data_1),
    .io_data_2(csa_9_io_data_2),
    .io_result_0(csa_9_io_result_0),
    .io_result_1(csa_9_io_result_1)
  );
  ysyx_22040886_csa csa_10 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_10_io_data_0),
    .io_data_1(csa_10_io_data_1),
    .io_data_2(csa_10_io_data_2),
    .io_result_0(csa_10_io_result_0),
    .io_result_1(csa_10_io_result_1)
  );
  ysyx_22040886_csa csa_11 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_11_io_data_0),
    .io_data_1(csa_11_io_data_1),
    .io_data_2(csa_11_io_data_2),
    .io_result_0(csa_11_io_result_0),
    .io_result_1(csa_11_io_result_1)
  );
  ysyx_22040886_csa csa_12 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_12_io_data_0),
    .io_data_1(csa_12_io_data_1),
    .io_data_2(csa_12_io_data_2),
    .io_result_0(csa_12_io_result_0),
    .io_result_1(csa_12_io_result_1)
  );
  ysyx_22040886_csa csa_13 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_13_io_data_0),
    .io_data_1(csa_13_io_data_1),
    .io_data_2(csa_13_io_data_2),
    .io_result_0(csa_13_io_result_0),
    .io_result_1(csa_13_io_result_1)
  );
  ysyx_22040886_csa csa_14 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_14_io_data_0),
    .io_data_1(csa_14_io_data_1),
    .io_data_2(csa_14_io_data_2),
    .io_result_0(csa_14_io_result_0),
    .io_result_1(csa_14_io_result_1)
  );
  ysyx_22040886_csa csa_15 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_15_io_data_0),
    .io_data_1(csa_15_io_data_1),
    .io_data_2(csa_15_io_data_2),
    .io_result_0(csa_15_io_result_0),
    .io_result_1(csa_15_io_result_1)
  );
  ysyx_22040886_csa csa_16 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_16_io_data_0),
    .io_data_1(csa_16_io_data_1),
    .io_data_2(csa_16_io_data_2),
    .io_result_0(csa_16_io_result_0),
    .io_result_1(csa_16_io_result_1)
  );
  ysyx_22040886_csa csa_17 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_17_io_data_0),
    .io_data_1(csa_17_io_data_1),
    .io_data_2(csa_17_io_data_2),
    .io_result_0(csa_17_io_result_0),
    .io_result_1(csa_17_io_result_1)
  );
  ysyx_22040886_csa csa_18 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_18_io_data_0),
    .io_data_1(csa_18_io_data_1),
    .io_data_2(csa_18_io_data_2),
    .io_result_0(csa_18_io_result_0),
    .io_result_1(csa_18_io_result_1)
  );
  ysyx_22040886_csa csa_19 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_19_io_data_0),
    .io_data_1(csa_19_io_data_1),
    .io_data_2(csa_19_io_data_2),
    .io_result_0(csa_19_io_result_0),
    .io_result_1(csa_19_io_result_1)
  );
  ysyx_22040886_csa csa_20 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_20_io_data_0),
    .io_data_1(csa_20_io_data_1),
    .io_data_2(csa_20_io_data_2),
    .io_result_0(csa_20_io_result_0),
    .io_result_1(csa_20_io_result_1)
  );
  ysyx_22040886_csa csa_21 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_21_io_data_0),
    .io_data_1(csa_21_io_data_1),
    .io_data_2(csa_21_io_data_2),
    .io_result_0(csa_21_io_result_0),
    .io_result_1(csa_21_io_result_1)
  );
  ysyx_22040886_csa csa_22 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_22_io_data_0),
    .io_data_1(csa_22_io_data_1),
    .io_data_2(csa_22_io_data_2),
    .io_result_0(csa_22_io_result_0),
    .io_result_1(csa_22_io_result_1)
  );
  ysyx_22040886_csa csa_23 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_23_io_data_0),
    .io_data_1(csa_23_io_data_1),
    .io_data_2(csa_23_io_data_2),
    .io_result_0(csa_23_io_result_0),
    .io_result_1(csa_23_io_result_1)
  );
  ysyx_22040886_csa csa_24 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_24_io_data_0),
    .io_data_1(csa_24_io_data_1),
    .io_data_2(csa_24_io_data_2),
    .io_result_0(csa_24_io_result_0),
    .io_result_1(csa_24_io_result_1)
  );
  ysyx_22040886_csa csa_25 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_25_io_data_0),
    .io_data_1(csa_25_io_data_1),
    .io_data_2(csa_25_io_data_2),
    .io_result_0(csa_25_io_result_0),
    .io_result_1(csa_25_io_result_1)
  );
  ysyx_22040886_csa csa_26 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_26_io_data_0),
    .io_data_1(csa_26_io_data_1),
    .io_data_2(csa_26_io_data_2),
    .io_result_0(csa_26_io_result_0),
    .io_result_1(csa_26_io_result_1)
  );
  ysyx_22040886_csa csa_27 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_27_io_data_0),
    .io_data_1(csa_27_io_data_1),
    .io_data_2(csa_27_io_data_2),
    .io_result_0(csa_27_io_result_0),
    .io_result_1(csa_27_io_result_1)
  );
  ysyx_22040886_csa csa_28 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_28_io_data_0),
    .io_data_1(csa_28_io_data_1),
    .io_data_2(csa_28_io_data_2),
    .io_result_0(csa_28_io_result_0),
    .io_result_1(csa_28_io_result_1)
  );
  ysyx_22040886_csa csa_29 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_29_io_data_0),
    .io_data_1(csa_29_io_data_1),
    .io_data_2(csa_29_io_data_2),
    .io_result_0(csa_29_io_result_0),
    .io_result_1(csa_29_io_result_1)
  );
  ysyx_22040886_csa csa_30 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_30_io_data_0),
    .io_data_1(csa_30_io_data_1),
    .io_data_2(csa_30_io_data_2),
    .io_result_0(csa_30_io_result_0),
    .io_result_1(csa_30_io_result_1)
  );
  assign io_result = vec_data_0 + vec_data_1; // @[hard_cal.scala 236:30]
  assign csa_io_data_0 = io_data_in_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_io_data_1 = io_data_in_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_io_data_2 = io_data_in_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_0 = io_data_in_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_1 = io_data_in_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_2 = io_data_in_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_0 = io_data_in_6; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_1 = io_data_in_7; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_2 = io_data_in_8; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_0 = io_data_in_9; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_1 = io_data_in_10; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_2 = io_data_in_11; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_0 = io_data_in_12; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_1 = io_data_in_13; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_2 = io_data_in_14; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_0 = io_data_in_15; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_1 = io_data_in_16; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_2 = io_data_in_17; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_0 = io_data_in_18; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_1 = io_data_in_19; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_2 = io_data_in_20; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_0 = io_data_in_21; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_1 = io_data_in_22; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_2 = io_data_in_23; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_0 = io_data_in_24; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_1 = io_data_in_25; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_2 = io_data_in_26; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_0 = io_data_in_27; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_1 = io_data_in_28; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_2 = io_data_in_29; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_0 = io_data_in_30; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_1 = io_data_in_31; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_2 = io_data_in_32; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_0 = vec_data_out_data_reg__0; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_1 = vec_data_out_data_reg__1; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_2 = vec_data_out_data_reg__2; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_0 = vec_data_out_data_reg__3; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_1 = vec_data_out_data_reg__4; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_2 = vec_data_out_data_reg__5; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_0 = vec_data_out_data_reg__6; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_1 = vec_data_out_data_reg__7; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_2 = vec_data_out_data_reg__8; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_0 = vec_data_out_data_reg__9; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_1 = vec_data_out_data_reg__10; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_2 = vec_data_out_data_reg__11; // @[hard_cal.scala 209:36 213:58]
  assign csa_15_io_data_0 = vec_data_out_data_reg__12; // @[hard_cal.scala 209:36 213:58]
  assign csa_15_io_data_1 = vec_data_out_data_reg__13; // @[hard_cal.scala 209:36 213:58]
  assign csa_15_io_data_2 = vec_data_out_data_reg__14; // @[hard_cal.scala 209:36 213:58]
  assign csa_16_io_data_0 = vec_data_out_data_reg__15; // @[hard_cal.scala 209:36 213:58]
  assign csa_16_io_data_1 = vec_data_out_data_reg__16; // @[hard_cal.scala 209:36 213:58]
  assign csa_16_io_data_2 = vec_data_out_data_reg__17; // @[hard_cal.scala 209:36 213:58]
  assign csa_17_io_data_0 = vec_data_out_data_reg__18; // @[hard_cal.scala 209:36 213:58]
  assign csa_17_io_data_1 = vec_data_out_data_reg__19; // @[hard_cal.scala 209:36 213:58]
  assign csa_17_io_data_2 = vec_data_out_data_reg__20; // @[hard_cal.scala 209:36 213:58]
  assign csa_18_io_data_0 = vec_data_out_data_reg_1_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_18_io_data_1 = vec_data_out_data_reg_1_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_18_io_data_2 = vec_data_out_data_reg_1_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_19_io_data_0 = vec_data_out_data_reg_1_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_19_io_data_1 = vec_data_out_data_reg_1_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_19_io_data_2 = vec_data_out_data_reg_1_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_20_io_data_0 = vec_data_out_data_reg_1_6; // @[hard_cal.scala 209:36 213:58]
  assign csa_20_io_data_1 = vec_data_out_data_reg_1_7; // @[hard_cal.scala 209:36 213:58]
  assign csa_20_io_data_2 = vec_data_out_data_reg_1_8; // @[hard_cal.scala 209:36 213:58]
  assign csa_21_io_data_0 = vec_data_out_data_reg_1_9; // @[hard_cal.scala 209:36 213:58]
  assign csa_21_io_data_1 = vec_data_out_data_reg_1_10; // @[hard_cal.scala 209:36 213:58]
  assign csa_21_io_data_2 = vec_data_out_data_reg_1_11; // @[hard_cal.scala 209:36 213:58]
  assign csa_22_io_data_0 = vec_data_out_data_reg_1_12; // @[hard_cal.scala 209:36 213:58]
  assign csa_22_io_data_1 = vec_data_out_data_reg_1_13; // @[hard_cal.scala 209:36 213:58]
  assign csa_22_io_data_2 = vec_data_out_data_reg_1_14; // @[hard_cal.scala 209:36 213:58]
  assign csa_23_io_data_0 = vec_data_out_data_reg_2_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_23_io_data_1 = vec_data_out_data_reg_2_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_23_io_data_2 = vec_data_out_data_reg_2_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_24_io_data_0 = vec_data_out_data_reg_2_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_24_io_data_1 = vec_data_out_data_reg_2_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_24_io_data_2 = vec_data_out_data_reg_2_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_25_io_data_0 = vec_data_out_data_reg_2_6; // @[hard_cal.scala 209:36 213:58]
  assign csa_25_io_data_1 = vec_data_out_data_reg_2_7; // @[hard_cal.scala 209:36 213:58]
  assign csa_25_io_data_2 = vec_data_out_data_reg_2_8; // @[hard_cal.scala 209:36 213:58]
  assign csa_26_io_data_0 = vec_data_out_data_reg_3_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_26_io_data_1 = vec_data_out_data_reg_3_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_26_io_data_2 = vec_data_out_data_reg_3_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_27_io_data_0 = vec_data_out_data_reg_3_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_27_io_data_1 = vec_data_out_data_reg_3_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_27_io_data_2 = vec_data_out_data_reg_3_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_28_io_data_0 = vec_data_out_data_reg_4_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_28_io_data_1 = vec_data_out_data_reg_4_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_28_io_data_2 = vec_data_out_data_reg_4_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_29_io_data_0 = vec_data_out_data_reg_5_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_29_io_data_1 = vec_data_out_data_reg_5_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_29_io_data_2 = vec_data_out_data_reg_5_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_30_io_data_0 = vec_data_out_data_reg_6_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_30_io_data_1 = vec_data_out_data_reg_6_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_30_io_data_2 = vec_data_out_data_reg_6_2; // @[hard_cal.scala 209:36 213:58]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__0 <= vec_data_csa_adder__0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__1 <= vec_data_csa_adder__0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__2 <= vec_data_csa_adder__1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__3 <= vec_data_csa_adder__1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__4 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__4 <= vec_data_csa_adder__2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__5 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__5 <= vec_data_csa_adder__2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__6 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__6 <= vec_data_csa_adder__3_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__7 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__7 <= vec_data_csa_adder__3_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__8 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__8 <= vec_data_csa_adder__4_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__9 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__9 <= vec_data_csa_adder__4_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__10 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__10 <= vec_data_csa_adder__5_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__11 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__11 <= vec_data_csa_adder__5_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__12 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__12 <= vec_data_csa_adder__6_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__13 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__13 <= vec_data_csa_adder__6_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__14 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__14 <= vec_data_csa_adder__7_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__15 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__15 <= vec_data_csa_adder__7_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__16 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__16 <= vec_data_csa_adder__8_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__17 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__17 <= vec_data_csa_adder__8_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__18 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__18 <= vec_data_csa_adder__9_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__19 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__19 <= vec_data_csa_adder__9_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__20 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__20 <= vec_data_csa_adder__10_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__21 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__21 <= vec_data_csa_adder__10_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_0 <= vec_data_csa_adder_1_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_1 <= vec_data_csa_adder_1_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_2 <= vec_data_csa_adder_1_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_3 <= vec_data_csa_adder_1_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_4 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_4 <= vec_data_csa_adder_1_2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_5 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_5 <= vec_data_csa_adder_1_2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_6 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_6 <= vec_data_csa_adder_1_3_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_7 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_7 <= vec_data_csa_adder_1_3_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_8 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_8 <= vec_data_csa_adder_1_4_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_9 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_9 <= vec_data_csa_adder_1_4_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_10 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_10 <= vec_data_csa_adder_1_5_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_11 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_11 <= vec_data_csa_adder_1_5_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_12 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_12 <= vec_data_csa_adder_1_6_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_13 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_13 <= vec_data_csa_adder_1_6_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_14 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_14 <= vec_data_out_data_reg__21; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_0 <= vec_data_csa_adder_2_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_1 <= vec_data_csa_adder_2_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_2 <= vec_data_csa_adder_2_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_3 <= vec_data_csa_adder_2_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_4 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_4 <= vec_data_csa_adder_2_2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_5 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_5 <= vec_data_csa_adder_2_2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_6 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_6 <= vec_data_csa_adder_2_3_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_7 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_7 <= vec_data_csa_adder_2_3_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_8 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_8 <= vec_data_csa_adder_2_4_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_9 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_9 <= vec_data_csa_adder_2_4_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_0 <= vec_data_csa_adder_3_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_1 <= vec_data_csa_adder_3_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_2 <= vec_data_csa_adder_3_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_3 <= vec_data_csa_adder_3_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_4 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_4 <= vec_data_csa_adder_3_2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_5 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_5 <= vec_data_csa_adder_3_2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_6 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_6 <= vec_data_out_data_reg_2_9; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_0 <= vec_data_csa_adder_4_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_1 <= vec_data_csa_adder_4_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_2 <= vec_data_csa_adder_4_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_3 <= vec_data_csa_adder_4_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_4 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_4 <= vec_data_out_data_reg_3_6; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_5_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_5_0 <= vec_data_csa_adder_5_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_5_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_5_1 <= vec_data_csa_adder_5_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_5_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_5_2 <= vec_data_out_data_reg_4_3; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_5_3 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_5_3 <= vec_data_out_data_reg_4_4; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_6_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_6_0 <= vec_data_csa_adder_6_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_6_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_6_1 <= vec_data_csa_adder_6_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_6_2 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_6_2 <= vec_data_out_data_reg_5_3; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_0 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_0 <= vec_data_csa_adder_7_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_1 <= 132'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_1 <= vec_data_csa_adder_7_0_result_1; // @[hard_cal.scala 226:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  vec_data_out_data_reg__0 = _RAND_0[131:0];
  _RAND_1 = {5{`RANDOM}};
  vec_data_out_data_reg__1 = _RAND_1[131:0];
  _RAND_2 = {5{`RANDOM}};
  vec_data_out_data_reg__2 = _RAND_2[131:0];
  _RAND_3 = {5{`RANDOM}};
  vec_data_out_data_reg__3 = _RAND_3[131:0];
  _RAND_4 = {5{`RANDOM}};
  vec_data_out_data_reg__4 = _RAND_4[131:0];
  _RAND_5 = {5{`RANDOM}};
  vec_data_out_data_reg__5 = _RAND_5[131:0];
  _RAND_6 = {5{`RANDOM}};
  vec_data_out_data_reg__6 = _RAND_6[131:0];
  _RAND_7 = {5{`RANDOM}};
  vec_data_out_data_reg__7 = _RAND_7[131:0];
  _RAND_8 = {5{`RANDOM}};
  vec_data_out_data_reg__8 = _RAND_8[131:0];
  _RAND_9 = {5{`RANDOM}};
  vec_data_out_data_reg__9 = _RAND_9[131:0];
  _RAND_10 = {5{`RANDOM}};
  vec_data_out_data_reg__10 = _RAND_10[131:0];
  _RAND_11 = {5{`RANDOM}};
  vec_data_out_data_reg__11 = _RAND_11[131:0];
  _RAND_12 = {5{`RANDOM}};
  vec_data_out_data_reg__12 = _RAND_12[131:0];
  _RAND_13 = {5{`RANDOM}};
  vec_data_out_data_reg__13 = _RAND_13[131:0];
  _RAND_14 = {5{`RANDOM}};
  vec_data_out_data_reg__14 = _RAND_14[131:0];
  _RAND_15 = {5{`RANDOM}};
  vec_data_out_data_reg__15 = _RAND_15[131:0];
  _RAND_16 = {5{`RANDOM}};
  vec_data_out_data_reg__16 = _RAND_16[131:0];
  _RAND_17 = {5{`RANDOM}};
  vec_data_out_data_reg__17 = _RAND_17[131:0];
  _RAND_18 = {5{`RANDOM}};
  vec_data_out_data_reg__18 = _RAND_18[131:0];
  _RAND_19 = {5{`RANDOM}};
  vec_data_out_data_reg__19 = _RAND_19[131:0];
  _RAND_20 = {5{`RANDOM}};
  vec_data_out_data_reg__20 = _RAND_20[131:0];
  _RAND_21 = {5{`RANDOM}};
  vec_data_out_data_reg__21 = _RAND_21[131:0];
  _RAND_22 = {5{`RANDOM}};
  vec_data_out_data_reg_1_0 = _RAND_22[131:0];
  _RAND_23 = {5{`RANDOM}};
  vec_data_out_data_reg_1_1 = _RAND_23[131:0];
  _RAND_24 = {5{`RANDOM}};
  vec_data_out_data_reg_1_2 = _RAND_24[131:0];
  _RAND_25 = {5{`RANDOM}};
  vec_data_out_data_reg_1_3 = _RAND_25[131:0];
  _RAND_26 = {5{`RANDOM}};
  vec_data_out_data_reg_1_4 = _RAND_26[131:0];
  _RAND_27 = {5{`RANDOM}};
  vec_data_out_data_reg_1_5 = _RAND_27[131:0];
  _RAND_28 = {5{`RANDOM}};
  vec_data_out_data_reg_1_6 = _RAND_28[131:0];
  _RAND_29 = {5{`RANDOM}};
  vec_data_out_data_reg_1_7 = _RAND_29[131:0];
  _RAND_30 = {5{`RANDOM}};
  vec_data_out_data_reg_1_8 = _RAND_30[131:0];
  _RAND_31 = {5{`RANDOM}};
  vec_data_out_data_reg_1_9 = _RAND_31[131:0];
  _RAND_32 = {5{`RANDOM}};
  vec_data_out_data_reg_1_10 = _RAND_32[131:0];
  _RAND_33 = {5{`RANDOM}};
  vec_data_out_data_reg_1_11 = _RAND_33[131:0];
  _RAND_34 = {5{`RANDOM}};
  vec_data_out_data_reg_1_12 = _RAND_34[131:0];
  _RAND_35 = {5{`RANDOM}};
  vec_data_out_data_reg_1_13 = _RAND_35[131:0];
  _RAND_36 = {5{`RANDOM}};
  vec_data_out_data_reg_1_14 = _RAND_36[131:0];
  _RAND_37 = {5{`RANDOM}};
  vec_data_out_data_reg_2_0 = _RAND_37[131:0];
  _RAND_38 = {5{`RANDOM}};
  vec_data_out_data_reg_2_1 = _RAND_38[131:0];
  _RAND_39 = {5{`RANDOM}};
  vec_data_out_data_reg_2_2 = _RAND_39[131:0];
  _RAND_40 = {5{`RANDOM}};
  vec_data_out_data_reg_2_3 = _RAND_40[131:0];
  _RAND_41 = {5{`RANDOM}};
  vec_data_out_data_reg_2_4 = _RAND_41[131:0];
  _RAND_42 = {5{`RANDOM}};
  vec_data_out_data_reg_2_5 = _RAND_42[131:0];
  _RAND_43 = {5{`RANDOM}};
  vec_data_out_data_reg_2_6 = _RAND_43[131:0];
  _RAND_44 = {5{`RANDOM}};
  vec_data_out_data_reg_2_7 = _RAND_44[131:0];
  _RAND_45 = {5{`RANDOM}};
  vec_data_out_data_reg_2_8 = _RAND_45[131:0];
  _RAND_46 = {5{`RANDOM}};
  vec_data_out_data_reg_2_9 = _RAND_46[131:0];
  _RAND_47 = {5{`RANDOM}};
  vec_data_out_data_reg_3_0 = _RAND_47[131:0];
  _RAND_48 = {5{`RANDOM}};
  vec_data_out_data_reg_3_1 = _RAND_48[131:0];
  _RAND_49 = {5{`RANDOM}};
  vec_data_out_data_reg_3_2 = _RAND_49[131:0];
  _RAND_50 = {5{`RANDOM}};
  vec_data_out_data_reg_3_3 = _RAND_50[131:0];
  _RAND_51 = {5{`RANDOM}};
  vec_data_out_data_reg_3_4 = _RAND_51[131:0];
  _RAND_52 = {5{`RANDOM}};
  vec_data_out_data_reg_3_5 = _RAND_52[131:0];
  _RAND_53 = {5{`RANDOM}};
  vec_data_out_data_reg_3_6 = _RAND_53[131:0];
  _RAND_54 = {5{`RANDOM}};
  vec_data_out_data_reg_4_0 = _RAND_54[131:0];
  _RAND_55 = {5{`RANDOM}};
  vec_data_out_data_reg_4_1 = _RAND_55[131:0];
  _RAND_56 = {5{`RANDOM}};
  vec_data_out_data_reg_4_2 = _RAND_56[131:0];
  _RAND_57 = {5{`RANDOM}};
  vec_data_out_data_reg_4_3 = _RAND_57[131:0];
  _RAND_58 = {5{`RANDOM}};
  vec_data_out_data_reg_4_4 = _RAND_58[131:0];
  _RAND_59 = {5{`RANDOM}};
  vec_data_out_data_reg_5_0 = _RAND_59[131:0];
  _RAND_60 = {5{`RANDOM}};
  vec_data_out_data_reg_5_1 = _RAND_60[131:0];
  _RAND_61 = {5{`RANDOM}};
  vec_data_out_data_reg_5_2 = _RAND_61[131:0];
  _RAND_62 = {5{`RANDOM}};
  vec_data_out_data_reg_5_3 = _RAND_62[131:0];
  _RAND_63 = {5{`RANDOM}};
  vec_data_out_data_reg_6_0 = _RAND_63[131:0];
  _RAND_64 = {5{`RANDOM}};
  vec_data_out_data_reg_6_1 = _RAND_64[131:0];
  _RAND_65 = {5{`RANDOM}};
  vec_data_out_data_reg_6_2 = _RAND_65[131:0];
  _RAND_66 = {5{`RANDOM}};
  vec_data_0 = _RAND_66[131:0];
  _RAND_67 = {5{`RANDOM}};
  vec_data_1 = _RAND_67[131:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_mul_hard(
  input         clock,
  input         reset,
  output [65:0] io_result_0,
  output [65:0] io_result_1,
  input  [65:0] io_data_0,
  input  [65:0] io_data_1,
  input         io_input_valid,
  output        io_Output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  cal_module_clock; // @[hard_cal.scala 300:28]
  wire  cal_module_reset; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_0; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_1; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_2; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_3; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_4; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_5; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_6; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_7; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_8; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_9; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_10; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_11; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_12; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_13; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_14; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_15; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_16; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_17; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_18; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_19; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_20; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_21; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_22; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_23; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_24; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_25; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_26; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_27; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_28; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_29; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_30; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_31; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_data_in_32; // @[hard_cal.scala 300:28]
  wire [131:0] cal_module_io_result; // @[hard_cal.scala 300:28]
  reg [131:0] regs_0; // @[hard_cal.scala 259:23]
  reg [131:0] regs_1; // @[hard_cal.scala 259:23]
  reg [6:0] counter; // @[hard_cal.scala 261:26]
  reg  cal_start; // @[hard_cal.scala 262:28]
  wire [6:0] _counter_T_1 = counter + 7'h1; // @[hard_cal.scala 264:39]
  wire  input_ready_to_be = ~cal_start; // @[hard_cal.scala 311:26]
  wire  _signed_T = io_input_valid & input_ready_to_be; // @[hard_cal.scala 265:35]
  reg [131:0] result_reg; // @[hard_cal.scala 266:29]
  reg [131:0] x_fu; // @[hard_cal.scala 269:23]
  wire [2:0] look_up_data = {regs_1[1],regs_1[0],1'h0}; // @[Cat.scala 31:58]
  wire [132:0] _booth_data_0_T = {regs_0, 1'h0}; // @[hard_cal.scala 284:38]
  wire [132:0] _booth_data_0_T_1 = {x_fu, 1'h0}; // @[hard_cal.scala 285:31]
  wire [131:0] _booth_data_0_T_3 = 3'h1 == look_up_data ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_0_T_5 = 3'h2 == look_up_data ? regs_0 : _booth_data_0_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_7 = 3'h3 == look_up_data ? _booth_data_0_T : {{1'd0}, _booth_data_0_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_9 = 3'h4 == look_up_data ? _booth_data_0_T_1 : _booth_data_0_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_11 = 3'h5 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_13 = 3'h6 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_15 = 3'h7 == look_up_data ? 133'h0 : _booth_data_0_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_0_T_17 = {1'h0,_booth_data_0_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_0_T_18 = {{1'd0}, _booth_data_0_T_17}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_1 = {regs_1[3],regs_1[2],regs_1[1]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_1_T_3 = 3'h1 == look_up_data_1 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_1_T_5 = 3'h2 == look_up_data_1 ? regs_0 : _booth_data_1_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_7 = 3'h3 == look_up_data_1 ? _booth_data_0_T : {{1'd0}, _booth_data_1_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_9 = 3'h4 == look_up_data_1 ? _booth_data_0_T_1 : _booth_data_1_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_11 = 3'h5 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_13 = 3'h6 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_15 = 3'h7 == look_up_data_1 ? 133'h0 : _booth_data_1_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_1_T_17 = {1'h0,_booth_data_1_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [68:0] _GEN_0 = {_booth_data_1_T_17, 2'h0}; // @[hard_cal.scala 290:19]
  wire [69:0] _booth_data_1_T_18 = {{1'd0}, _GEN_0}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_2 = {regs_1[5],regs_1[4],regs_1[3]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_2_T_3 = 3'h1 == look_up_data_2 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_2_T_5 = 3'h2 == look_up_data_2 ? regs_0 : _booth_data_2_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_7 = 3'h3 == look_up_data_2 ? _booth_data_0_T : {{1'd0}, _booth_data_2_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_9 = 3'h4 == look_up_data_2 ? _booth_data_0_T_1 : _booth_data_2_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_11 = 3'h5 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_13 = 3'h6 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_15 = 3'h7 == look_up_data_2 ? 133'h0 : _booth_data_2_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_2_T_17 = {1'h0,_booth_data_2_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [70:0] _GEN_1 = {_booth_data_2_T_17, 4'h0}; // @[hard_cal.scala 290:19]
  wire [73:0] _booth_data_2_T_18 = {{3'd0}, _GEN_1}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_3 = {regs_1[7],regs_1[6],regs_1[5]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_3_T_3 = 3'h1 == look_up_data_3 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_3_T_5 = 3'h2 == look_up_data_3 ? regs_0 : _booth_data_3_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_7 = 3'h3 == look_up_data_3 ? _booth_data_0_T : {{1'd0}, _booth_data_3_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_9 = 3'h4 == look_up_data_3 ? _booth_data_0_T_1 : _booth_data_3_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_11 = 3'h5 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_13 = 3'h6 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_15 = 3'h7 == look_up_data_3 ? 133'h0 : _booth_data_3_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_3_T_17 = {1'h0,_booth_data_3_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [72:0] _GEN_2 = {_booth_data_3_T_17, 6'h0}; // @[hard_cal.scala 290:19]
  wire [73:0] _booth_data_3_T_18 = {{1'd0}, _GEN_2}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_4 = {regs_1[9],regs_1[8],regs_1[7]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_4_T_3 = 3'h1 == look_up_data_4 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_4_T_5 = 3'h2 == look_up_data_4 ? regs_0 : _booth_data_4_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_7 = 3'h3 == look_up_data_4 ? _booth_data_0_T : {{1'd0}, _booth_data_4_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_9 = 3'h4 == look_up_data_4 ? _booth_data_0_T_1 : _booth_data_4_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_11 = 3'h5 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_13 = 3'h6 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_15 = 3'h7 == look_up_data_4 ? 133'h0 : _booth_data_4_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_4_T_17 = {1'h0,_booth_data_4_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [74:0] _GEN_3 = {_booth_data_4_T_17, 8'h0}; // @[hard_cal.scala 290:19]
  wire [81:0] _booth_data_4_T_18 = {{7'd0}, _GEN_3}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_5 = {regs_1[11],regs_1[10],regs_1[9]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_5_T_3 = 3'h1 == look_up_data_5 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_5_T_5 = 3'h2 == look_up_data_5 ? regs_0 : _booth_data_5_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_7 = 3'h3 == look_up_data_5 ? _booth_data_0_T : {{1'd0}, _booth_data_5_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_9 = 3'h4 == look_up_data_5 ? _booth_data_0_T_1 : _booth_data_5_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_11 = 3'h5 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_13 = 3'h6 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_15 = 3'h7 == look_up_data_5 ? 133'h0 : _booth_data_5_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_5_T_17 = {1'h0,_booth_data_5_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [76:0] _GEN_4 = {_booth_data_5_T_17, 10'h0}; // @[hard_cal.scala 290:19]
  wire [81:0] _booth_data_5_T_18 = {{5'd0}, _GEN_4}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_6 = {regs_1[13],regs_1[12],regs_1[11]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_6_T_3 = 3'h1 == look_up_data_6 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_6_T_5 = 3'h2 == look_up_data_6 ? regs_0 : _booth_data_6_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_7 = 3'h3 == look_up_data_6 ? _booth_data_0_T : {{1'd0}, _booth_data_6_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_9 = 3'h4 == look_up_data_6 ? _booth_data_0_T_1 : _booth_data_6_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_11 = 3'h5 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_13 = 3'h6 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_15 = 3'h7 == look_up_data_6 ? 133'h0 : _booth_data_6_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_6_T_17 = {1'h0,_booth_data_6_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [78:0] _GEN_5 = {_booth_data_6_T_17, 12'h0}; // @[hard_cal.scala 290:19]
  wire [81:0] _booth_data_6_T_18 = {{3'd0}, _GEN_5}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_7 = {regs_1[15],regs_1[14],regs_1[13]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_7_T_3 = 3'h1 == look_up_data_7 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_7_T_5 = 3'h2 == look_up_data_7 ? regs_0 : _booth_data_7_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_7 = 3'h3 == look_up_data_7 ? _booth_data_0_T : {{1'd0}, _booth_data_7_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_9 = 3'h4 == look_up_data_7 ? _booth_data_0_T_1 : _booth_data_7_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_11 = 3'h5 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_13 = 3'h6 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_15 = 3'h7 == look_up_data_7 ? 133'h0 : _booth_data_7_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_7_T_17 = {1'h0,_booth_data_7_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [80:0] _GEN_6 = {_booth_data_7_T_17, 14'h0}; // @[hard_cal.scala 290:19]
  wire [81:0] _booth_data_7_T_18 = {{1'd0}, _GEN_6}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_8 = {regs_1[17],regs_1[16],regs_1[15]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_8_T_3 = 3'h1 == look_up_data_8 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_8_T_5 = 3'h2 == look_up_data_8 ? regs_0 : _booth_data_8_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_7 = 3'h3 == look_up_data_8 ? _booth_data_0_T : {{1'd0}, _booth_data_8_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_9 = 3'h4 == look_up_data_8 ? _booth_data_0_T_1 : _booth_data_8_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_11 = 3'h5 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_13 = 3'h6 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_15 = 3'h7 == look_up_data_8 ? 133'h0 : _booth_data_8_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_8_T_17 = {1'h0,_booth_data_8_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [82:0] _GEN_7 = {_booth_data_8_T_17, 16'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_8_T_18 = {{15'd0}, _GEN_7}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_9 = {regs_1[19],regs_1[18],regs_1[17]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_9_T_3 = 3'h1 == look_up_data_9 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_9_T_5 = 3'h2 == look_up_data_9 ? regs_0 : _booth_data_9_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_7 = 3'h3 == look_up_data_9 ? _booth_data_0_T : {{1'd0}, _booth_data_9_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_9 = 3'h4 == look_up_data_9 ? _booth_data_0_T_1 : _booth_data_9_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_11 = 3'h5 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_13 = 3'h6 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_15 = 3'h7 == look_up_data_9 ? 133'h0 : _booth_data_9_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_9_T_17 = {1'h0,_booth_data_9_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [84:0] _GEN_8 = {_booth_data_9_T_17, 18'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_9_T_18 = {{13'd0}, _GEN_8}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_10 = {regs_1[21],regs_1[20],regs_1[19]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_10_T_3 = 3'h1 == look_up_data_10 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_10_T_5 = 3'h2 == look_up_data_10 ? regs_0 : _booth_data_10_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_7 = 3'h3 == look_up_data_10 ? _booth_data_0_T : {{1'd0}, _booth_data_10_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_9 = 3'h4 == look_up_data_10 ? _booth_data_0_T_1 : _booth_data_10_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_11 = 3'h5 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_13 = 3'h6 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_15 = 3'h7 == look_up_data_10 ? 133'h0 : _booth_data_10_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_10_T_17 = {1'h0,_booth_data_10_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [86:0] _GEN_9 = {_booth_data_10_T_17, 20'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_10_T_18 = {{11'd0}, _GEN_9}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_11 = {regs_1[23],regs_1[22],regs_1[21]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_11_T_3 = 3'h1 == look_up_data_11 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_11_T_5 = 3'h2 == look_up_data_11 ? regs_0 : _booth_data_11_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_7 = 3'h3 == look_up_data_11 ? _booth_data_0_T : {{1'd0}, _booth_data_11_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_9 = 3'h4 == look_up_data_11 ? _booth_data_0_T_1 : _booth_data_11_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_11 = 3'h5 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_13 = 3'h6 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_15 = 3'h7 == look_up_data_11 ? 133'h0 : _booth_data_11_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_11_T_17 = {1'h0,_booth_data_11_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [88:0] _GEN_10 = {_booth_data_11_T_17, 22'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_11_T_18 = {{9'd0}, _GEN_10}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_12 = {regs_1[25],regs_1[24],regs_1[23]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_12_T_3 = 3'h1 == look_up_data_12 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_12_T_5 = 3'h2 == look_up_data_12 ? regs_0 : _booth_data_12_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_7 = 3'h3 == look_up_data_12 ? _booth_data_0_T : {{1'd0}, _booth_data_12_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_9 = 3'h4 == look_up_data_12 ? _booth_data_0_T_1 : _booth_data_12_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_11 = 3'h5 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_13 = 3'h6 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_15 = 3'h7 == look_up_data_12 ? 133'h0 : _booth_data_12_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_12_T_17 = {1'h0,_booth_data_12_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [90:0] _GEN_11 = {_booth_data_12_T_17, 24'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_12_T_18 = {{7'd0}, _GEN_11}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_13 = {regs_1[27],regs_1[26],regs_1[25]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_13_T_3 = 3'h1 == look_up_data_13 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_13_T_5 = 3'h2 == look_up_data_13 ? regs_0 : _booth_data_13_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_7 = 3'h3 == look_up_data_13 ? _booth_data_0_T : {{1'd0}, _booth_data_13_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_9 = 3'h4 == look_up_data_13 ? _booth_data_0_T_1 : _booth_data_13_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_11 = 3'h5 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_13 = 3'h6 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_15 = 3'h7 == look_up_data_13 ? 133'h0 : _booth_data_13_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_13_T_17 = {1'h0,_booth_data_13_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [92:0] _GEN_12 = {_booth_data_13_T_17, 26'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_13_T_18 = {{5'd0}, _GEN_12}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_14 = {regs_1[29],regs_1[28],regs_1[27]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_14_T_3 = 3'h1 == look_up_data_14 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_14_T_5 = 3'h2 == look_up_data_14 ? regs_0 : _booth_data_14_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_7 = 3'h3 == look_up_data_14 ? _booth_data_0_T : {{1'd0}, _booth_data_14_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_9 = 3'h4 == look_up_data_14 ? _booth_data_0_T_1 : _booth_data_14_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_11 = 3'h5 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_13 = 3'h6 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_15 = 3'h7 == look_up_data_14 ? 133'h0 : _booth_data_14_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_14_T_17 = {1'h0,_booth_data_14_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [94:0] _GEN_13 = {_booth_data_14_T_17, 28'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_14_T_18 = {{3'd0}, _GEN_13}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_15 = {regs_1[31],regs_1[30],regs_1[29]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_15_T_3 = 3'h1 == look_up_data_15 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_15_T_5 = 3'h2 == look_up_data_15 ? regs_0 : _booth_data_15_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_7 = 3'h3 == look_up_data_15 ? _booth_data_0_T : {{1'd0}, _booth_data_15_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_9 = 3'h4 == look_up_data_15 ? _booth_data_0_T_1 : _booth_data_15_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_11 = 3'h5 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_13 = 3'h6 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_15 = 3'h7 == look_up_data_15 ? 133'h0 : _booth_data_15_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_15_T_17 = {1'h0,_booth_data_15_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [96:0] _GEN_14 = {_booth_data_15_T_17, 30'h0}; // @[hard_cal.scala 290:19]
  wire [97:0] _booth_data_15_T_18 = {{1'd0}, _GEN_14}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_16 = {regs_1[33],regs_1[32],regs_1[31]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_16_T_3 = 3'h1 == look_up_data_16 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_16_T_5 = 3'h2 == look_up_data_16 ? regs_0 : _booth_data_16_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_7 = 3'h3 == look_up_data_16 ? _booth_data_0_T : {{1'd0}, _booth_data_16_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_9 = 3'h4 == look_up_data_16 ? _booth_data_0_T_1 : _booth_data_16_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_11 = 3'h5 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_13 = 3'h6 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_15 = 3'h7 == look_up_data_16 ? 133'h0 : _booth_data_16_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_16_T_17 = {1'h0,_booth_data_16_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [98:0] _GEN_15 = {_booth_data_16_T_17, 32'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_16_T_18 = {{31'd0}, _GEN_15}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_17 = {regs_1[35],regs_1[34],regs_1[33]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_17_T_3 = 3'h1 == look_up_data_17 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_17_T_5 = 3'h2 == look_up_data_17 ? regs_0 : _booth_data_17_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_7 = 3'h3 == look_up_data_17 ? _booth_data_0_T : {{1'd0}, _booth_data_17_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_9 = 3'h4 == look_up_data_17 ? _booth_data_0_T_1 : _booth_data_17_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_11 = 3'h5 == look_up_data_17 ? {{1'd0}, x_fu} : _booth_data_17_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_13 = 3'h6 == look_up_data_17 ? {{1'd0}, x_fu} : _booth_data_17_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_15 = 3'h7 == look_up_data_17 ? 133'h0 : _booth_data_17_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_17_T_17 = {1'h0,_booth_data_17_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [100:0] _GEN_16 = {_booth_data_17_T_17, 34'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_17_T_18 = {{29'd0}, _GEN_16}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_18 = {regs_1[37],regs_1[36],regs_1[35]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_18_T_3 = 3'h1 == look_up_data_18 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_18_T_5 = 3'h2 == look_up_data_18 ? regs_0 : _booth_data_18_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_7 = 3'h3 == look_up_data_18 ? _booth_data_0_T : {{1'd0}, _booth_data_18_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_9 = 3'h4 == look_up_data_18 ? _booth_data_0_T_1 : _booth_data_18_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_11 = 3'h5 == look_up_data_18 ? {{1'd0}, x_fu} : _booth_data_18_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_13 = 3'h6 == look_up_data_18 ? {{1'd0}, x_fu} : _booth_data_18_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_15 = 3'h7 == look_up_data_18 ? 133'h0 : _booth_data_18_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_18_T_17 = {1'h0,_booth_data_18_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [102:0] _GEN_17 = {_booth_data_18_T_17, 36'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_18_T_18 = {{27'd0}, _GEN_17}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_19 = {regs_1[39],regs_1[38],regs_1[37]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_19_T_3 = 3'h1 == look_up_data_19 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_19_T_5 = 3'h2 == look_up_data_19 ? regs_0 : _booth_data_19_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_7 = 3'h3 == look_up_data_19 ? _booth_data_0_T : {{1'd0}, _booth_data_19_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_9 = 3'h4 == look_up_data_19 ? _booth_data_0_T_1 : _booth_data_19_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_11 = 3'h5 == look_up_data_19 ? {{1'd0}, x_fu} : _booth_data_19_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_13 = 3'h6 == look_up_data_19 ? {{1'd0}, x_fu} : _booth_data_19_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_15 = 3'h7 == look_up_data_19 ? 133'h0 : _booth_data_19_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_19_T_17 = {1'h0,_booth_data_19_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [104:0] _GEN_18 = {_booth_data_19_T_17, 38'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_19_T_18 = {{25'd0}, _GEN_18}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_20 = {regs_1[41],regs_1[40],regs_1[39]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_20_T_3 = 3'h1 == look_up_data_20 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_20_T_5 = 3'h2 == look_up_data_20 ? regs_0 : _booth_data_20_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_7 = 3'h3 == look_up_data_20 ? _booth_data_0_T : {{1'd0}, _booth_data_20_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_9 = 3'h4 == look_up_data_20 ? _booth_data_0_T_1 : _booth_data_20_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_11 = 3'h5 == look_up_data_20 ? {{1'd0}, x_fu} : _booth_data_20_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_13 = 3'h6 == look_up_data_20 ? {{1'd0}, x_fu} : _booth_data_20_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_15 = 3'h7 == look_up_data_20 ? 133'h0 : _booth_data_20_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_20_T_17 = {1'h0,_booth_data_20_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [106:0] _GEN_19 = {_booth_data_20_T_17, 40'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_20_T_18 = {{23'd0}, _GEN_19}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_21 = {regs_1[43],regs_1[42],regs_1[41]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_21_T_3 = 3'h1 == look_up_data_21 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_21_T_5 = 3'h2 == look_up_data_21 ? regs_0 : _booth_data_21_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_7 = 3'h3 == look_up_data_21 ? _booth_data_0_T : {{1'd0}, _booth_data_21_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_9 = 3'h4 == look_up_data_21 ? _booth_data_0_T_1 : _booth_data_21_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_11 = 3'h5 == look_up_data_21 ? {{1'd0}, x_fu} : _booth_data_21_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_13 = 3'h6 == look_up_data_21 ? {{1'd0}, x_fu} : _booth_data_21_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_15 = 3'h7 == look_up_data_21 ? 133'h0 : _booth_data_21_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_21_T_17 = {1'h0,_booth_data_21_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [108:0] _GEN_20 = {_booth_data_21_T_17, 42'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_21_T_18 = {{21'd0}, _GEN_20}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_22 = {regs_1[45],regs_1[44],regs_1[43]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_22_T_3 = 3'h1 == look_up_data_22 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_22_T_5 = 3'h2 == look_up_data_22 ? regs_0 : _booth_data_22_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_7 = 3'h3 == look_up_data_22 ? _booth_data_0_T : {{1'd0}, _booth_data_22_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_9 = 3'h4 == look_up_data_22 ? _booth_data_0_T_1 : _booth_data_22_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_11 = 3'h5 == look_up_data_22 ? {{1'd0}, x_fu} : _booth_data_22_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_13 = 3'h6 == look_up_data_22 ? {{1'd0}, x_fu} : _booth_data_22_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_15 = 3'h7 == look_up_data_22 ? 133'h0 : _booth_data_22_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_22_T_17 = {1'h0,_booth_data_22_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [110:0] _GEN_21 = {_booth_data_22_T_17, 44'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_22_T_18 = {{19'd0}, _GEN_21}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_23 = {regs_1[47],regs_1[46],regs_1[45]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_23_T_3 = 3'h1 == look_up_data_23 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_23_T_5 = 3'h2 == look_up_data_23 ? regs_0 : _booth_data_23_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_7 = 3'h3 == look_up_data_23 ? _booth_data_0_T : {{1'd0}, _booth_data_23_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_9 = 3'h4 == look_up_data_23 ? _booth_data_0_T_1 : _booth_data_23_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_11 = 3'h5 == look_up_data_23 ? {{1'd0}, x_fu} : _booth_data_23_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_13 = 3'h6 == look_up_data_23 ? {{1'd0}, x_fu} : _booth_data_23_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_15 = 3'h7 == look_up_data_23 ? 133'h0 : _booth_data_23_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_23_T_17 = {1'h0,_booth_data_23_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [112:0] _GEN_22 = {_booth_data_23_T_17, 46'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_23_T_18 = {{17'd0}, _GEN_22}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_24 = {regs_1[49],regs_1[48],regs_1[47]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_24_T_3 = 3'h1 == look_up_data_24 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_24_T_5 = 3'h2 == look_up_data_24 ? regs_0 : _booth_data_24_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_7 = 3'h3 == look_up_data_24 ? _booth_data_0_T : {{1'd0}, _booth_data_24_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_9 = 3'h4 == look_up_data_24 ? _booth_data_0_T_1 : _booth_data_24_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_11 = 3'h5 == look_up_data_24 ? {{1'd0}, x_fu} : _booth_data_24_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_13 = 3'h6 == look_up_data_24 ? {{1'd0}, x_fu} : _booth_data_24_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_15 = 3'h7 == look_up_data_24 ? 133'h0 : _booth_data_24_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_24_T_17 = {1'h0,_booth_data_24_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [114:0] _GEN_23 = {_booth_data_24_T_17, 48'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_24_T_18 = {{15'd0}, _GEN_23}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_25 = {regs_1[51],regs_1[50],regs_1[49]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_25_T_3 = 3'h1 == look_up_data_25 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_25_T_5 = 3'h2 == look_up_data_25 ? regs_0 : _booth_data_25_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_7 = 3'h3 == look_up_data_25 ? _booth_data_0_T : {{1'd0}, _booth_data_25_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_9 = 3'h4 == look_up_data_25 ? _booth_data_0_T_1 : _booth_data_25_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_11 = 3'h5 == look_up_data_25 ? {{1'd0}, x_fu} : _booth_data_25_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_13 = 3'h6 == look_up_data_25 ? {{1'd0}, x_fu} : _booth_data_25_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_15 = 3'h7 == look_up_data_25 ? 133'h0 : _booth_data_25_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_25_T_17 = {1'h0,_booth_data_25_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [116:0] _GEN_24 = {_booth_data_25_T_17, 50'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_25_T_18 = {{13'd0}, _GEN_24}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_26 = {regs_1[53],regs_1[52],regs_1[51]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_26_T_3 = 3'h1 == look_up_data_26 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_26_T_5 = 3'h2 == look_up_data_26 ? regs_0 : _booth_data_26_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_7 = 3'h3 == look_up_data_26 ? _booth_data_0_T : {{1'd0}, _booth_data_26_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_9 = 3'h4 == look_up_data_26 ? _booth_data_0_T_1 : _booth_data_26_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_11 = 3'h5 == look_up_data_26 ? {{1'd0}, x_fu} : _booth_data_26_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_13 = 3'h6 == look_up_data_26 ? {{1'd0}, x_fu} : _booth_data_26_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_15 = 3'h7 == look_up_data_26 ? 133'h0 : _booth_data_26_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_26_T_17 = {1'h0,_booth_data_26_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [118:0] _GEN_25 = {_booth_data_26_T_17, 52'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_26_T_18 = {{11'd0}, _GEN_25}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_27 = {regs_1[55],regs_1[54],regs_1[53]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_27_T_3 = 3'h1 == look_up_data_27 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_27_T_5 = 3'h2 == look_up_data_27 ? regs_0 : _booth_data_27_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_7 = 3'h3 == look_up_data_27 ? _booth_data_0_T : {{1'd0}, _booth_data_27_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_9 = 3'h4 == look_up_data_27 ? _booth_data_0_T_1 : _booth_data_27_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_11 = 3'h5 == look_up_data_27 ? {{1'd0}, x_fu} : _booth_data_27_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_13 = 3'h6 == look_up_data_27 ? {{1'd0}, x_fu} : _booth_data_27_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_15 = 3'h7 == look_up_data_27 ? 133'h0 : _booth_data_27_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_27_T_17 = {1'h0,_booth_data_27_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [120:0] _GEN_26 = {_booth_data_27_T_17, 54'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_27_T_18 = {{9'd0}, _GEN_26}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_28 = {regs_1[57],regs_1[56],regs_1[55]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_28_T_3 = 3'h1 == look_up_data_28 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_28_T_5 = 3'h2 == look_up_data_28 ? regs_0 : _booth_data_28_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_7 = 3'h3 == look_up_data_28 ? _booth_data_0_T : {{1'd0}, _booth_data_28_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_9 = 3'h4 == look_up_data_28 ? _booth_data_0_T_1 : _booth_data_28_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_11 = 3'h5 == look_up_data_28 ? {{1'd0}, x_fu} : _booth_data_28_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_13 = 3'h6 == look_up_data_28 ? {{1'd0}, x_fu} : _booth_data_28_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_15 = 3'h7 == look_up_data_28 ? 133'h0 : _booth_data_28_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_28_T_17 = {1'h0,_booth_data_28_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [122:0] _GEN_27 = {_booth_data_28_T_17, 56'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_28_T_18 = {{7'd0}, _GEN_27}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_29 = {regs_1[59],regs_1[58],regs_1[57]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_29_T_3 = 3'h1 == look_up_data_29 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_29_T_5 = 3'h2 == look_up_data_29 ? regs_0 : _booth_data_29_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_7 = 3'h3 == look_up_data_29 ? _booth_data_0_T : {{1'd0}, _booth_data_29_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_9 = 3'h4 == look_up_data_29 ? _booth_data_0_T_1 : _booth_data_29_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_11 = 3'h5 == look_up_data_29 ? {{1'd0}, x_fu} : _booth_data_29_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_13 = 3'h6 == look_up_data_29 ? {{1'd0}, x_fu} : _booth_data_29_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_15 = 3'h7 == look_up_data_29 ? 133'h0 : _booth_data_29_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_29_T_17 = {1'h0,_booth_data_29_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [124:0] _GEN_28 = {_booth_data_29_T_17, 58'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_29_T_18 = {{5'd0}, _GEN_28}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_30 = {regs_1[61],regs_1[60],regs_1[59]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_30_T_3 = 3'h1 == look_up_data_30 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_30_T_5 = 3'h2 == look_up_data_30 ? regs_0 : _booth_data_30_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_7 = 3'h3 == look_up_data_30 ? _booth_data_0_T : {{1'd0}, _booth_data_30_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_9 = 3'h4 == look_up_data_30 ? _booth_data_0_T_1 : _booth_data_30_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_11 = 3'h5 == look_up_data_30 ? {{1'd0}, x_fu} : _booth_data_30_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_13 = 3'h6 == look_up_data_30 ? {{1'd0}, x_fu} : _booth_data_30_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_15 = 3'h7 == look_up_data_30 ? 133'h0 : _booth_data_30_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_30_T_17 = {1'h0,_booth_data_30_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [126:0] _GEN_29 = {_booth_data_30_T_17, 60'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_30_T_18 = {{3'd0}, _GEN_29}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_31 = {regs_1[63],regs_1[62],regs_1[61]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_31_T_3 = 3'h1 == look_up_data_31 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_31_T_5 = 3'h2 == look_up_data_31 ? regs_0 : _booth_data_31_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_7 = 3'h3 == look_up_data_31 ? _booth_data_0_T : {{1'd0}, _booth_data_31_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_9 = 3'h4 == look_up_data_31 ? _booth_data_0_T_1 : _booth_data_31_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_11 = 3'h5 == look_up_data_31 ? {{1'd0}, x_fu} : _booth_data_31_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_13 = 3'h6 == look_up_data_31 ? {{1'd0}, x_fu} : _booth_data_31_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_15 = 3'h7 == look_up_data_31 ? 133'h0 : _booth_data_31_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_31_T_17 = {1'h0,_booth_data_31_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [128:0] _GEN_30 = {_booth_data_31_T_17, 62'h0}; // @[hard_cal.scala 290:19]
  wire [129:0] _booth_data_31_T_18 = {{1'd0}, _GEN_30}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_32 = {regs_1[65],regs_1[64],regs_1[63]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_32_T_3 = 3'h1 == look_up_data_32 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_32_T_5 = 3'h2 == look_up_data_32 ? regs_0 : _booth_data_32_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_7 = 3'h3 == look_up_data_32 ? _booth_data_0_T : {{1'd0}, _booth_data_32_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_9 = 3'h4 == look_up_data_32 ? _booth_data_0_T_1 : _booth_data_32_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_11 = 3'h5 == look_up_data_32 ? {{1'd0}, x_fu} : _booth_data_32_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_13 = 3'h6 == look_up_data_32 ? {{1'd0}, x_fu} : _booth_data_32_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_15 = 3'h7 == look_up_data_32 ? 133'h0 : _booth_data_32_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_32_T_17 = {1'h0,_booth_data_32_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [130:0] _GEN_31 = {_booth_data_32_T_17, 64'h0}; // @[hard_cal.scala 290:19]
  wire [193:0] _booth_data_32_T_18 = {{63'd0}, _GEN_31}; // @[hard_cal.scala 290:19]
  wire [65:0] _x_fu_T_1 = ~io_data_0; // @[hard_cal.scala 295:56]
  wire [65:0] _x_fu_T_3 = _x_fu_T_1 + 66'h1; // @[hard_cal.scala 295:70]
  wire [3:0] _cal_start_T_2 = 4'h9 - 4'h1; // @[hard_cal.scala 302:115]
  wire [6:0] _GEN_32 = {{3'd0}, _cal_start_T_2}; // @[hard_cal.scala 302:81]
  wire  _cal_start_T_4 = counter == _GEN_32 ? 1'h0 : cal_start; // @[hard_cal.scala 302:72]
  ysyx_22040886_wallace_adder cal_module ( // @[hard_cal.scala 300:28]
    .clock(cal_module_clock),
    .reset(cal_module_reset),
    .io_data_in_0(cal_module_io_data_in_0),
    .io_data_in_1(cal_module_io_data_in_1),
    .io_data_in_2(cal_module_io_data_in_2),
    .io_data_in_3(cal_module_io_data_in_3),
    .io_data_in_4(cal_module_io_data_in_4),
    .io_data_in_5(cal_module_io_data_in_5),
    .io_data_in_6(cal_module_io_data_in_6),
    .io_data_in_7(cal_module_io_data_in_7),
    .io_data_in_8(cal_module_io_data_in_8),
    .io_data_in_9(cal_module_io_data_in_9),
    .io_data_in_10(cal_module_io_data_in_10),
    .io_data_in_11(cal_module_io_data_in_11),
    .io_data_in_12(cal_module_io_data_in_12),
    .io_data_in_13(cal_module_io_data_in_13),
    .io_data_in_14(cal_module_io_data_in_14),
    .io_data_in_15(cal_module_io_data_in_15),
    .io_data_in_16(cal_module_io_data_in_16),
    .io_data_in_17(cal_module_io_data_in_17),
    .io_data_in_18(cal_module_io_data_in_18),
    .io_data_in_19(cal_module_io_data_in_19),
    .io_data_in_20(cal_module_io_data_in_20),
    .io_data_in_21(cal_module_io_data_in_21),
    .io_data_in_22(cal_module_io_data_in_22),
    .io_data_in_23(cal_module_io_data_in_23),
    .io_data_in_24(cal_module_io_data_in_24),
    .io_data_in_25(cal_module_io_data_in_25),
    .io_data_in_26(cal_module_io_data_in_26),
    .io_data_in_27(cal_module_io_data_in_27),
    .io_data_in_28(cal_module_io_data_in_28),
    .io_data_in_29(cal_module_io_data_in_29),
    .io_data_in_30(cal_module_io_data_in_30),
    .io_data_in_31(cal_module_io_data_in_31),
    .io_data_in_32(cal_module_io_data_in_32),
    .io_result(cal_module_io_result)
  );
  assign io_result_0 = cal_start ? cal_module_io_result[65:0] : result_reg[65:0]; // @[hard_cal.scala 308:24]
  assign io_result_1 = cal_start ? cal_module_io_result[131:66] : result_reg[131:66]; // @[hard_cal.scala 309:24]
  assign io_Output_valid = counter == _GEN_32; // @[hard_cal.scala 310:34]
  assign cal_module_clock = clock;
  assign cal_module_reset = reset;
  assign cal_module_io_data_in_0 = {{64'd0}, _booth_data_0_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_1 = {{62'd0}, _booth_data_1_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_2 = {{58'd0}, _booth_data_2_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_3 = {{58'd0}, _booth_data_3_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_4 = {{50'd0}, _booth_data_4_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_5 = {{50'd0}, _booth_data_5_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_6 = {{50'd0}, _booth_data_6_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_7 = {{50'd0}, _booth_data_7_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_8 = {{34'd0}, _booth_data_8_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_9 = {{34'd0}, _booth_data_9_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_10 = {{34'd0}, _booth_data_10_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_11 = {{34'd0}, _booth_data_11_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_12 = {{34'd0}, _booth_data_12_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_13 = {{34'd0}, _booth_data_13_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_14 = {{34'd0}, _booth_data_14_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_15 = {{34'd0}, _booth_data_15_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_16 = {{2'd0}, _booth_data_16_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_17 = {{2'd0}, _booth_data_17_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_18 = {{2'd0}, _booth_data_18_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_19 = {{2'd0}, _booth_data_19_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_20 = {{2'd0}, _booth_data_20_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_21 = {{2'd0}, _booth_data_21_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_22 = {{2'd0}, _booth_data_22_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_23 = {{2'd0}, _booth_data_23_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_24 = {{2'd0}, _booth_data_24_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_25 = {{2'd0}, _booth_data_25_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_26 = {{2'd0}, _booth_data_26_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_27 = {{2'd0}, _booth_data_27_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_28 = {{2'd0}, _booth_data_28_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_29 = {{2'd0}, _booth_data_29_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_30 = {{2'd0}, _booth_data_30_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_31 = {{2'd0}, _booth_data_31_T_18}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_32 = _booth_data_32_T_18[131:0]; // @[hard_cal.scala 268:26 280:27]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 259:23]
      regs_0 <= 132'h0; // @[hard_cal.scala 259:23]
    end else if (_signed_T) begin // @[hard_cal.scala 294:19]
      regs_0 <= {{66'd0}, io_data_0};
    end
    if (reset) begin // @[hard_cal.scala 259:23]
      regs_1 <= 132'h0; // @[hard_cal.scala 259:23]
    end else if (_signed_T) begin // @[hard_cal.scala 296:19]
      regs_1 <= {{66'd0}, io_data_1};
    end
    if (reset) begin // @[hard_cal.scala 261:26]
      counter <= 7'h0; // @[hard_cal.scala 261:26]
    end else if (cal_start) begin // @[hard_cal.scala 264:19]
      counter <= _counter_T_1;
    end else begin
      counter <= 7'h0;
    end
    if (reset) begin // @[hard_cal.scala 262:28]
      cal_start <= 1'h0; // @[hard_cal.scala 262:28]
    end else begin
      cal_start <= _signed_T | _cal_start_T_4; // @[hard_cal.scala 302:15]
    end
    if (reset) begin // @[hard_cal.scala 266:29]
      result_reg <= 132'h0; // @[hard_cal.scala 266:29]
    end else if (cal_start) begin // @[hard_cal.scala 307:22]
      result_reg <= cal_module_io_result;
    end
    if (reset) begin // @[hard_cal.scala 269:23]
      x_fu <= 132'h0; // @[hard_cal.scala 269:23]
    end else if (_signed_T) begin // @[hard_cal.scala 295:18]
      x_fu <= {{66'd0}, _x_fu_T_3};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  regs_0 = _RAND_0[131:0];
  _RAND_1 = {5{`RANDOM}};
  regs_1 = _RAND_1[131:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {5{`RANDOM}};
  result_reg = _RAND_4[131:0];
  _RAND_5 = {5{`RANDOM}};
  x_fu = _RAND_5[131:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_csa_31(
  input  [67:0] io_data_0,
  input  [67:0] io_data_1,
  input  [67:0] io_data_2,
  output [67:0] io_result_0,
  output [67:0] io_result_1
);
  wire [67:0] _io_result_0_T = io_data_0 ^ io_data_1; // @[hard_cal.scala 187:32]
  wire [67:0] _io_result_1_T = io_data_0 & io_data_1; // @[hard_cal.scala 188:37]
  wire [67:0] _io_result_1_T_1 = io_data_1 & io_data_2; // @[hard_cal.scala 188:65]
  wire [67:0] _io_result_1_T_2 = _io_result_1_T | _io_result_1_T_1; // @[hard_cal.scala 188:51]
  wire [67:0] _io_result_1_T_3 = io_data_2 & io_data_0; // @[hard_cal.scala 188:93]
  wire [67:0] _io_result_1_T_4 = _io_result_1_T_2 | _io_result_1_T_3; // @[hard_cal.scala 188:79]
  wire [68:0] _io_result_1_T_5 = {_io_result_1_T_4,1'h0}; // @[Cat.scala 31:58]
  assign io_result_0 = _io_result_0_T ^ io_data_2; // @[hard_cal.scala 187:45]
  assign io_result_1 = _io_result_1_T_5[67:0]; // @[hard_cal.scala 188:18]
endmodule
module ysyx_22040886_wallace_adder_1(
  input         clock,
  input         reset,
  input  [67:0] io_data_in_0,
  input  [67:0] io_data_in_1,
  input  [67:0] io_data_in_2,
  input  [67:0] io_data_in_3,
  input  [67:0] io_data_in_4,
  input  [67:0] io_data_in_5,
  input  [67:0] io_data_in_6,
  input  [67:0] io_data_in_7,
  input  [67:0] io_data_in_8,
  input  [67:0] io_data_in_9,
  input  [67:0] io_data_in_10,
  input  [67:0] io_data_in_11,
  input  [67:0] io_data_in_12,
  input  [67:0] io_data_in_13,
  input  [67:0] io_data_in_14,
  input  [67:0] io_data_in_15,
  input  [67:0] io_data_in_16,
  output [67:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [95:0] _RAND_20;
  reg [95:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [95:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  wire [67:0] csa_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_1_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_1_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_1_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_1_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_1_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_2_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_2_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_2_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_2_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_2_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_3_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_3_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_3_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_3_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_3_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_4_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_4_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_4_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_4_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_4_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_5_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_5_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_5_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_5_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_5_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_6_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_6_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_6_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_6_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_6_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_7_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_7_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_7_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_7_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_7_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_8_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_8_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_8_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_8_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_8_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_9_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_9_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_9_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_9_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_9_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_10_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_10_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_10_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_10_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_10_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_11_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_11_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_11_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_11_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_11_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_12_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_12_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_12_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_12_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_12_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_13_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_13_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_13_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_13_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_13_io_result_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_14_io_data_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_14_io_data_1; // @[hard_cal.scala 209:61]
  wire [67:0] csa_14_io_data_2; // @[hard_cal.scala 209:61]
  wire [67:0] csa_14_io_result_0; // @[hard_cal.scala 209:61]
  wire [67:0] csa_14_io_result_1; // @[hard_cal.scala 209:61]
  reg [67:0] vec_data_out_data_reg__0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__1; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__2; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__3; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__4; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__5; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__6; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__7; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__8; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__9; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__10; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg__11; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_1; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_2; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_3; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_4; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_5; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_6; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_1_7; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_1; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_2; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_3; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_4; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_2_5; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_3_0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_3_1; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_3_2; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_3_3; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_4_0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_4_1; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_out_data_reg_4_2; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_0; // @[hard_cal.scala 225:39]
  reg [67:0] vec_data_1; // @[hard_cal.scala 225:39]
  wire [67:0] vec_data_csa_adder__0_result_0 = csa_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__0_result_1 = csa_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__1_result_0 = csa_1_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__1_result_1 = csa_1_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__2_result_0 = csa_2_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__2_result_1 = csa_2_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__3_result_0 = csa_3_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__3_result_1 = csa_3_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__4_result_0 = csa_4_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder__4_result_1 = csa_4_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_0_result_0 = csa_5_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_0_result_1 = csa_5_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_1_result_0 = csa_6_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_1_result_1 = csa_6_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_2_result_0 = csa_7_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_2_result_1 = csa_7_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_3_result_0 = csa_8_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_1_3_result_1 = csa_8_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_2_0_result_0 = csa_9_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_2_0_result_1 = csa_9_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_2_1_result_0 = csa_10_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_2_1_result_1 = csa_10_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_3_0_result_0 = csa_11_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_3_0_result_1 = csa_11_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_3_1_result_0 = csa_12_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_3_1_result_1 = csa_12_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_4_0_result_0 = csa_13_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_4_0_result_1 = csa_13_io_result_1; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_5_0_result_0 = csa_14_io_result_0; // @[hard_cal.scala 209:{36,36}]
  wire [67:0] vec_data_csa_adder_5_0_result_1 = csa_14_io_result_1; // @[hard_cal.scala 209:{36,36}]
  ysyx_22040886_csa_31 csa ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_io_data_0),
    .io_data_1(csa_io_data_1),
    .io_data_2(csa_io_data_2),
    .io_result_0(csa_io_result_0),
    .io_result_1(csa_io_result_1)
  );
  ysyx_22040886_csa_31 csa_1 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_1_io_data_0),
    .io_data_1(csa_1_io_data_1),
    .io_data_2(csa_1_io_data_2),
    .io_result_0(csa_1_io_result_0),
    .io_result_1(csa_1_io_result_1)
  );
  ysyx_22040886_csa_31 csa_2 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_2_io_data_0),
    .io_data_1(csa_2_io_data_1),
    .io_data_2(csa_2_io_data_2),
    .io_result_0(csa_2_io_result_0),
    .io_result_1(csa_2_io_result_1)
  );
  ysyx_22040886_csa_31 csa_3 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_3_io_data_0),
    .io_data_1(csa_3_io_data_1),
    .io_data_2(csa_3_io_data_2),
    .io_result_0(csa_3_io_result_0),
    .io_result_1(csa_3_io_result_1)
  );
  ysyx_22040886_csa_31 csa_4 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_4_io_data_0),
    .io_data_1(csa_4_io_data_1),
    .io_data_2(csa_4_io_data_2),
    .io_result_0(csa_4_io_result_0),
    .io_result_1(csa_4_io_result_1)
  );
  ysyx_22040886_csa_31 csa_5 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_5_io_data_0),
    .io_data_1(csa_5_io_data_1),
    .io_data_2(csa_5_io_data_2),
    .io_result_0(csa_5_io_result_0),
    .io_result_1(csa_5_io_result_1)
  );
  ysyx_22040886_csa_31 csa_6 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_6_io_data_0),
    .io_data_1(csa_6_io_data_1),
    .io_data_2(csa_6_io_data_2),
    .io_result_0(csa_6_io_result_0),
    .io_result_1(csa_6_io_result_1)
  );
  ysyx_22040886_csa_31 csa_7 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_7_io_data_0),
    .io_data_1(csa_7_io_data_1),
    .io_data_2(csa_7_io_data_2),
    .io_result_0(csa_7_io_result_0),
    .io_result_1(csa_7_io_result_1)
  );
  ysyx_22040886_csa_31 csa_8 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_8_io_data_0),
    .io_data_1(csa_8_io_data_1),
    .io_data_2(csa_8_io_data_2),
    .io_result_0(csa_8_io_result_0),
    .io_result_1(csa_8_io_result_1)
  );
  ysyx_22040886_csa_31 csa_9 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_9_io_data_0),
    .io_data_1(csa_9_io_data_1),
    .io_data_2(csa_9_io_data_2),
    .io_result_0(csa_9_io_result_0),
    .io_result_1(csa_9_io_result_1)
  );
  ysyx_22040886_csa_31 csa_10 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_10_io_data_0),
    .io_data_1(csa_10_io_data_1),
    .io_data_2(csa_10_io_data_2),
    .io_result_0(csa_10_io_result_0),
    .io_result_1(csa_10_io_result_1)
  );
  ysyx_22040886_csa_31 csa_11 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_11_io_data_0),
    .io_data_1(csa_11_io_data_1),
    .io_data_2(csa_11_io_data_2),
    .io_result_0(csa_11_io_result_0),
    .io_result_1(csa_11_io_result_1)
  );
  ysyx_22040886_csa_31 csa_12 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_12_io_data_0),
    .io_data_1(csa_12_io_data_1),
    .io_data_2(csa_12_io_data_2),
    .io_result_0(csa_12_io_result_0),
    .io_result_1(csa_12_io_result_1)
  );
  ysyx_22040886_csa_31 csa_13 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_13_io_data_0),
    .io_data_1(csa_13_io_data_1),
    .io_data_2(csa_13_io_data_2),
    .io_result_0(csa_13_io_result_0),
    .io_result_1(csa_13_io_result_1)
  );
  ysyx_22040886_csa_31 csa_14 ( // @[hard_cal.scala 209:61]
    .io_data_0(csa_14_io_data_0),
    .io_data_1(csa_14_io_data_1),
    .io_data_2(csa_14_io_data_2),
    .io_result_0(csa_14_io_result_0),
    .io_result_1(csa_14_io_result_1)
  );
  assign io_result = vec_data_0 + vec_data_1; // @[hard_cal.scala 236:30]
  assign csa_io_data_0 = io_data_in_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_io_data_1 = io_data_in_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_io_data_2 = io_data_in_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_0 = io_data_in_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_1 = io_data_in_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_1_io_data_2 = io_data_in_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_0 = io_data_in_6; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_1 = io_data_in_7; // @[hard_cal.scala 209:36 213:58]
  assign csa_2_io_data_2 = io_data_in_8; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_0 = io_data_in_9; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_1 = io_data_in_10; // @[hard_cal.scala 209:36 213:58]
  assign csa_3_io_data_2 = io_data_in_11; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_0 = io_data_in_12; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_1 = io_data_in_13; // @[hard_cal.scala 209:36 213:58]
  assign csa_4_io_data_2 = io_data_in_14; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_0 = vec_data_out_data_reg__0; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_1 = vec_data_out_data_reg__1; // @[hard_cal.scala 209:36 213:58]
  assign csa_5_io_data_2 = vec_data_out_data_reg__2; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_0 = vec_data_out_data_reg__3; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_1 = vec_data_out_data_reg__4; // @[hard_cal.scala 209:36 213:58]
  assign csa_6_io_data_2 = vec_data_out_data_reg__5; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_0 = vec_data_out_data_reg__6; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_1 = vec_data_out_data_reg__7; // @[hard_cal.scala 209:36 213:58]
  assign csa_7_io_data_2 = vec_data_out_data_reg__8; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_0 = vec_data_out_data_reg__9; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_1 = vec_data_out_data_reg__10; // @[hard_cal.scala 209:36 213:58]
  assign csa_8_io_data_2 = vec_data_out_data_reg__11; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_0 = vec_data_out_data_reg_1_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_1 = vec_data_out_data_reg_1_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_9_io_data_2 = vec_data_out_data_reg_1_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_0 = vec_data_out_data_reg_1_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_1 = vec_data_out_data_reg_1_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_10_io_data_2 = vec_data_out_data_reg_1_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_0 = vec_data_out_data_reg_2_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_1 = vec_data_out_data_reg_2_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_11_io_data_2 = vec_data_out_data_reg_2_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_0 = vec_data_out_data_reg_2_3; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_1 = vec_data_out_data_reg_2_4; // @[hard_cal.scala 209:36 213:58]
  assign csa_12_io_data_2 = vec_data_out_data_reg_2_5; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_0 = vec_data_out_data_reg_3_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_1 = vec_data_out_data_reg_3_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_13_io_data_2 = vec_data_out_data_reg_3_2; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_0 = vec_data_out_data_reg_4_0; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_1 = vec_data_out_data_reg_4_1; // @[hard_cal.scala 209:36 213:58]
  assign csa_14_io_data_2 = vec_data_out_data_reg_4_2; // @[hard_cal.scala 209:36 213:58]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__0 <= vec_data_csa_adder__0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__1 <= vec_data_csa_adder__0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__2 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__2 <= vec_data_csa_adder__1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__3 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__3 <= vec_data_csa_adder__1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__4 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__4 <= vec_data_csa_adder__2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__5 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__5 <= vec_data_csa_adder__2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__6 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__6 <= vec_data_csa_adder__3_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__7 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__7 <= vec_data_csa_adder__3_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__8 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__8 <= vec_data_csa_adder__4_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__9 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__9 <= vec_data_csa_adder__4_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__10 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__10 <= io_data_in_15; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg__11 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg__11 <= io_data_in_16; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_0 <= vec_data_csa_adder_1_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_1 <= vec_data_csa_adder_1_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_2 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_2 <= vec_data_csa_adder_1_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_3 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_3 <= vec_data_csa_adder_1_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_4 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_4 <= vec_data_csa_adder_1_2_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_5 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_5 <= vec_data_csa_adder_1_2_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_6 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_6 <= vec_data_csa_adder_1_3_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_1_7 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_1_7 <= vec_data_csa_adder_1_3_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_0 <= vec_data_csa_adder_2_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_1 <= vec_data_csa_adder_2_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_2 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_2 <= vec_data_csa_adder_2_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_3 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_3 <= vec_data_csa_adder_2_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_4 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_4 <= vec_data_out_data_reg_1_6; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_2_5 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_2_5 <= vec_data_out_data_reg_1_7; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_0 <= vec_data_csa_adder_3_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_1 <= vec_data_csa_adder_3_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_2 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_2 <= vec_data_csa_adder_3_1_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_3_3 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_3_3 <= vec_data_csa_adder_3_1_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_0 <= vec_data_csa_adder_4_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_1 <= vec_data_csa_adder_4_0_result_1; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_out_data_reg_4_2 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_out_data_reg_4_2 <= vec_data_out_data_reg_3_3; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_0 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_0 <= vec_data_csa_adder_5_0_result_0; // @[hard_cal.scala 226:26]
    end
    if (reset) begin // @[hard_cal.scala 225:39]
      vec_data_1 <= 68'h0; // @[hard_cal.scala 225:39]
    end else begin
      vec_data_1 <= vec_data_csa_adder_5_0_result_1; // @[hard_cal.scala 226:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  vec_data_out_data_reg__0 = _RAND_0[67:0];
  _RAND_1 = {3{`RANDOM}};
  vec_data_out_data_reg__1 = _RAND_1[67:0];
  _RAND_2 = {3{`RANDOM}};
  vec_data_out_data_reg__2 = _RAND_2[67:0];
  _RAND_3 = {3{`RANDOM}};
  vec_data_out_data_reg__3 = _RAND_3[67:0];
  _RAND_4 = {3{`RANDOM}};
  vec_data_out_data_reg__4 = _RAND_4[67:0];
  _RAND_5 = {3{`RANDOM}};
  vec_data_out_data_reg__5 = _RAND_5[67:0];
  _RAND_6 = {3{`RANDOM}};
  vec_data_out_data_reg__6 = _RAND_6[67:0];
  _RAND_7 = {3{`RANDOM}};
  vec_data_out_data_reg__7 = _RAND_7[67:0];
  _RAND_8 = {3{`RANDOM}};
  vec_data_out_data_reg__8 = _RAND_8[67:0];
  _RAND_9 = {3{`RANDOM}};
  vec_data_out_data_reg__9 = _RAND_9[67:0];
  _RAND_10 = {3{`RANDOM}};
  vec_data_out_data_reg__10 = _RAND_10[67:0];
  _RAND_11 = {3{`RANDOM}};
  vec_data_out_data_reg__11 = _RAND_11[67:0];
  _RAND_12 = {3{`RANDOM}};
  vec_data_out_data_reg_1_0 = _RAND_12[67:0];
  _RAND_13 = {3{`RANDOM}};
  vec_data_out_data_reg_1_1 = _RAND_13[67:0];
  _RAND_14 = {3{`RANDOM}};
  vec_data_out_data_reg_1_2 = _RAND_14[67:0];
  _RAND_15 = {3{`RANDOM}};
  vec_data_out_data_reg_1_3 = _RAND_15[67:0];
  _RAND_16 = {3{`RANDOM}};
  vec_data_out_data_reg_1_4 = _RAND_16[67:0];
  _RAND_17 = {3{`RANDOM}};
  vec_data_out_data_reg_1_5 = _RAND_17[67:0];
  _RAND_18 = {3{`RANDOM}};
  vec_data_out_data_reg_1_6 = _RAND_18[67:0];
  _RAND_19 = {3{`RANDOM}};
  vec_data_out_data_reg_1_7 = _RAND_19[67:0];
  _RAND_20 = {3{`RANDOM}};
  vec_data_out_data_reg_2_0 = _RAND_20[67:0];
  _RAND_21 = {3{`RANDOM}};
  vec_data_out_data_reg_2_1 = _RAND_21[67:0];
  _RAND_22 = {3{`RANDOM}};
  vec_data_out_data_reg_2_2 = _RAND_22[67:0];
  _RAND_23 = {3{`RANDOM}};
  vec_data_out_data_reg_2_3 = _RAND_23[67:0];
  _RAND_24 = {3{`RANDOM}};
  vec_data_out_data_reg_2_4 = _RAND_24[67:0];
  _RAND_25 = {3{`RANDOM}};
  vec_data_out_data_reg_2_5 = _RAND_25[67:0];
  _RAND_26 = {3{`RANDOM}};
  vec_data_out_data_reg_3_0 = _RAND_26[67:0];
  _RAND_27 = {3{`RANDOM}};
  vec_data_out_data_reg_3_1 = _RAND_27[67:0];
  _RAND_28 = {3{`RANDOM}};
  vec_data_out_data_reg_3_2 = _RAND_28[67:0];
  _RAND_29 = {3{`RANDOM}};
  vec_data_out_data_reg_3_3 = _RAND_29[67:0];
  _RAND_30 = {3{`RANDOM}};
  vec_data_out_data_reg_4_0 = _RAND_30[67:0];
  _RAND_31 = {3{`RANDOM}};
  vec_data_out_data_reg_4_1 = _RAND_31[67:0];
  _RAND_32 = {3{`RANDOM}};
  vec_data_out_data_reg_4_2 = _RAND_32[67:0];
  _RAND_33 = {3{`RANDOM}};
  vec_data_0 = _RAND_33[67:0];
  _RAND_34 = {3{`RANDOM}};
  vec_data_1 = _RAND_34[67:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_mul_hard_1(
  input         clock,
  input         reset,
  output [33:0] io_result_0,
  input  [33:0] io_data_0,
  input  [33:0] io_data_1,
  input         io_input_valid,
  output        io_Output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  cal_module_clock; // @[hard_cal.scala 300:28]
  wire  cal_module_reset; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_0; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_1; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_2; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_3; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_4; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_5; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_6; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_7; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_8; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_9; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_10; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_11; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_12; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_13; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_14; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_15; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_data_in_16; // @[hard_cal.scala 300:28]
  wire [67:0] cal_module_io_result; // @[hard_cal.scala 300:28]
  reg [67:0] regs_0; // @[hard_cal.scala 259:23]
  reg [67:0] regs_1; // @[hard_cal.scala 259:23]
  reg [5:0] counter; // @[hard_cal.scala 261:26]
  reg  cal_start; // @[hard_cal.scala 262:28]
  wire [5:0] _counter_T_1 = counter + 6'h1; // @[hard_cal.scala 264:39]
  wire  input_ready_to_be = ~cal_start; // @[hard_cal.scala 311:26]
  wire  _signed_T = io_input_valid & input_ready_to_be; // @[hard_cal.scala 265:35]
  reg [67:0] result_reg; // @[hard_cal.scala 266:29]
  reg [67:0] x_fu; // @[hard_cal.scala 269:23]
  wire [2:0] look_up_data = {regs_1[1],regs_1[0],1'h0}; // @[Cat.scala 31:58]
  wire [68:0] _booth_data_0_T = {regs_0, 1'h0}; // @[hard_cal.scala 284:38]
  wire [68:0] _booth_data_0_T_1 = {x_fu, 1'h0}; // @[hard_cal.scala 285:31]
  wire [67:0] _booth_data_0_T_3 = 3'h1 == look_up_data ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_0_T_5 = 3'h2 == look_up_data ? regs_0 : _booth_data_0_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_7 = 3'h3 == look_up_data ? _booth_data_0_T : {{1'd0}, _booth_data_0_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_9 = 3'h4 == look_up_data ? _booth_data_0_T_1 : _booth_data_0_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_11 = 3'h5 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_13 = 3'h6 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_15 = 3'h7 == look_up_data ? 69'h0 : _booth_data_0_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_0_lo_lo = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    _booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_0_lo = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15
    [33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],booth_data_0_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_0_T_46 = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    _booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    booth_data_0_lo_lo,booth_data_0_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_0_T_48 = {_booth_data_0_T_46,_booth_data_0_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [64:0] _booth_data_0_T_49 = {{1'd0}, _booth_data_0_T_48}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_1 = {regs_1[3],regs_1[2],regs_1[1]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_1_T_3 = 3'h1 == look_up_data_1 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_1_T_5 = 3'h2 == look_up_data_1 ? regs_0 : _booth_data_1_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_7 = 3'h3 == look_up_data_1 ? _booth_data_0_T : {{1'd0}, _booth_data_1_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_9 = 3'h4 == look_up_data_1 ? _booth_data_0_T_1 : _booth_data_1_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_11 = 3'h5 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_13 = 3'h6 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_15 = 3'h7 == look_up_data_1 ? 69'h0 : _booth_data_1_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_1_lo_lo = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    _booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_1_lo = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15
    [33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],booth_data_1_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_1_T_46 = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    _booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    booth_data_1_lo_lo,booth_data_1_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_1_T_48 = {_booth_data_1_T_46,_booth_data_1_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [65:0] _GEN_0 = {_booth_data_1_T_48, 2'h0}; // @[hard_cal.scala 290:19]
  wire [66:0] _booth_data_1_T_49 = {{1'd0}, _GEN_0}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_2 = {regs_1[5],regs_1[4],regs_1[3]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_2_T_3 = 3'h1 == look_up_data_2 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_2_T_5 = 3'h2 == look_up_data_2 ? regs_0 : _booth_data_2_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_7 = 3'h3 == look_up_data_2 ? _booth_data_0_T : {{1'd0}, _booth_data_2_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_9 = 3'h4 == look_up_data_2 ? _booth_data_0_T_1 : _booth_data_2_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_11 = 3'h5 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_13 = 3'h6 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_15 = 3'h7 == look_up_data_2 ? 69'h0 : _booth_data_2_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_2_lo_lo = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    _booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_2_lo = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15
    [33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],booth_data_2_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_2_T_46 = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    _booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    booth_data_2_lo_lo,booth_data_2_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_2_T_48 = {_booth_data_2_T_46,_booth_data_2_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [67:0] _GEN_1 = {_booth_data_2_T_48, 4'h0}; // @[hard_cal.scala 290:19]
  wire [70:0] _booth_data_2_T_49 = {{3'd0}, _GEN_1}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_3 = {regs_1[7],regs_1[6],regs_1[5]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_3_T_3 = 3'h1 == look_up_data_3 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_3_T_5 = 3'h2 == look_up_data_3 ? regs_0 : _booth_data_3_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_7 = 3'h3 == look_up_data_3 ? _booth_data_0_T : {{1'd0}, _booth_data_3_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_9 = 3'h4 == look_up_data_3 ? _booth_data_0_T_1 : _booth_data_3_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_11 = 3'h5 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_13 = 3'h6 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_15 = 3'h7 == look_up_data_3 ? 69'h0 : _booth_data_3_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_3_lo_lo = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    _booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_3_lo = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15
    [33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],booth_data_3_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_3_T_46 = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    _booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    booth_data_3_lo_lo,booth_data_3_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_3_T_48 = {_booth_data_3_T_46,_booth_data_3_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [69:0] _GEN_2 = {_booth_data_3_T_48, 6'h0}; // @[hard_cal.scala 290:19]
  wire [70:0] _booth_data_3_T_49 = {{1'd0}, _GEN_2}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_4 = {regs_1[9],regs_1[8],regs_1[7]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_4_T_3 = 3'h1 == look_up_data_4 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_4_T_5 = 3'h2 == look_up_data_4 ? regs_0 : _booth_data_4_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_7 = 3'h3 == look_up_data_4 ? _booth_data_0_T : {{1'd0}, _booth_data_4_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_9 = 3'h4 == look_up_data_4 ? _booth_data_0_T_1 : _booth_data_4_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_11 = 3'h5 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_13 = 3'h6 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_15 = 3'h7 == look_up_data_4 ? 69'h0 : _booth_data_4_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_4_lo_lo = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    _booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_4_lo = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15
    [33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],booth_data_4_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_4_T_46 = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    _booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    booth_data_4_lo_lo,booth_data_4_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_4_T_48 = {_booth_data_4_T_46,_booth_data_4_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [71:0] _GEN_3 = {_booth_data_4_T_48, 8'h0}; // @[hard_cal.scala 290:19]
  wire [78:0] _booth_data_4_T_49 = {{7'd0}, _GEN_3}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_5 = {regs_1[11],regs_1[10],regs_1[9]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_5_T_3 = 3'h1 == look_up_data_5 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_5_T_5 = 3'h2 == look_up_data_5 ? regs_0 : _booth_data_5_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_7 = 3'h3 == look_up_data_5 ? _booth_data_0_T : {{1'd0}, _booth_data_5_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_9 = 3'h4 == look_up_data_5 ? _booth_data_0_T_1 : _booth_data_5_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_11 = 3'h5 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_13 = 3'h6 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_15 = 3'h7 == look_up_data_5 ? 69'h0 : _booth_data_5_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_5_lo_lo = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    _booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_5_lo = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15
    [33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],booth_data_5_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_5_T_46 = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    _booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    booth_data_5_lo_lo,booth_data_5_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_5_T_48 = {_booth_data_5_T_46,_booth_data_5_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [73:0] _GEN_4 = {_booth_data_5_T_48, 10'h0}; // @[hard_cal.scala 290:19]
  wire [78:0] _booth_data_5_T_49 = {{5'd0}, _GEN_4}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_6 = {regs_1[13],regs_1[12],regs_1[11]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_6_T_3 = 3'h1 == look_up_data_6 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_6_T_5 = 3'h2 == look_up_data_6 ? regs_0 : _booth_data_6_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_7 = 3'h3 == look_up_data_6 ? _booth_data_0_T : {{1'd0}, _booth_data_6_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_9 = 3'h4 == look_up_data_6 ? _booth_data_0_T_1 : _booth_data_6_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_11 = 3'h5 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_13 = 3'h6 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_15 = 3'h7 == look_up_data_6 ? 69'h0 : _booth_data_6_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_6_lo_lo = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    _booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_6_lo = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15
    [33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],booth_data_6_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_6_T_46 = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    _booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    booth_data_6_lo_lo,booth_data_6_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_6_T_48 = {_booth_data_6_T_46,_booth_data_6_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [75:0] _GEN_5 = {_booth_data_6_T_48, 12'h0}; // @[hard_cal.scala 290:19]
  wire [78:0] _booth_data_6_T_49 = {{3'd0}, _GEN_5}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_7 = {regs_1[15],regs_1[14],regs_1[13]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_7_T_3 = 3'h1 == look_up_data_7 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_7_T_5 = 3'h2 == look_up_data_7 ? regs_0 : _booth_data_7_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_7 = 3'h3 == look_up_data_7 ? _booth_data_0_T : {{1'd0}, _booth_data_7_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_9 = 3'h4 == look_up_data_7 ? _booth_data_0_T_1 : _booth_data_7_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_11 = 3'h5 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_13 = 3'h6 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_15 = 3'h7 == look_up_data_7 ? 69'h0 : _booth_data_7_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_7_lo_lo = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    _booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_7_lo = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15
    [33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],booth_data_7_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_7_T_46 = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    _booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    booth_data_7_lo_lo,booth_data_7_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_7_T_48 = {_booth_data_7_T_46,_booth_data_7_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [77:0] _GEN_6 = {_booth_data_7_T_48, 14'h0}; // @[hard_cal.scala 290:19]
  wire [78:0] _booth_data_7_T_49 = {{1'd0}, _GEN_6}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_8 = {regs_1[17],regs_1[16],regs_1[15]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_8_T_3 = 3'h1 == look_up_data_8 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_8_T_5 = 3'h2 == look_up_data_8 ? regs_0 : _booth_data_8_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_7 = 3'h3 == look_up_data_8 ? _booth_data_0_T : {{1'd0}, _booth_data_8_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_9 = 3'h4 == look_up_data_8 ? _booth_data_0_T_1 : _booth_data_8_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_11 = 3'h5 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_13 = 3'h6 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_15 = 3'h7 == look_up_data_8 ? 69'h0 : _booth_data_8_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_8_lo_lo = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    _booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_8_lo = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15
    [33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],booth_data_8_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_8_T_46 = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    _booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    booth_data_8_lo_lo,booth_data_8_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_8_T_48 = {_booth_data_8_T_46,_booth_data_8_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [79:0] _GEN_7 = {_booth_data_8_T_48, 16'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_8_T_49 = {{15'd0}, _GEN_7}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_9 = {regs_1[19],regs_1[18],regs_1[17]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_9_T_3 = 3'h1 == look_up_data_9 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_9_T_5 = 3'h2 == look_up_data_9 ? regs_0 : _booth_data_9_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_7 = 3'h3 == look_up_data_9 ? _booth_data_0_T : {{1'd0}, _booth_data_9_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_9 = 3'h4 == look_up_data_9 ? _booth_data_0_T_1 : _booth_data_9_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_11 = 3'h5 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_13 = 3'h6 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_15 = 3'h7 == look_up_data_9 ? 69'h0 : _booth_data_9_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_9_lo_lo = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    _booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_9_lo = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15
    [33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],booth_data_9_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_9_T_46 = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    _booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    booth_data_9_lo_lo,booth_data_9_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_9_T_48 = {_booth_data_9_T_46,_booth_data_9_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [81:0] _GEN_8 = {_booth_data_9_T_48, 18'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_9_T_49 = {{13'd0}, _GEN_8}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_10 = {regs_1[21],regs_1[20],regs_1[19]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_10_T_3 = 3'h1 == look_up_data_10 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_10_T_5 = 3'h2 == look_up_data_10 ? regs_0 : _booth_data_10_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_7 = 3'h3 == look_up_data_10 ? _booth_data_0_T : {{1'd0}, _booth_data_10_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_9 = 3'h4 == look_up_data_10 ? _booth_data_0_T_1 : _booth_data_10_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_11 = 3'h5 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_13 = 3'h6 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_15 = 3'h7 == look_up_data_10 ? 69'h0 : _booth_data_10_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_10_lo_lo = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_10_lo = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[
    33],booth_data_10_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_10_T_46 = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[
    33],booth_data_10_lo_lo,booth_data_10_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_10_T_48 = {_booth_data_10_T_46,_booth_data_10_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [83:0] _GEN_9 = {_booth_data_10_T_48, 20'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_10_T_49 = {{11'd0}, _GEN_9}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_11 = {regs_1[23],regs_1[22],regs_1[21]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_11_T_3 = 3'h1 == look_up_data_11 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_11_T_5 = 3'h2 == look_up_data_11 ? regs_0 : _booth_data_11_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_7 = 3'h3 == look_up_data_11 ? _booth_data_0_T : {{1'd0}, _booth_data_11_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_9 = 3'h4 == look_up_data_11 ? _booth_data_0_T_1 : _booth_data_11_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_11 = 3'h5 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_13 = 3'h6 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_15 = 3'h7 == look_up_data_11 ? 69'h0 : _booth_data_11_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_11_lo_lo = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_11_lo = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[
    33],booth_data_11_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_11_T_46 = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[
    33],booth_data_11_lo_lo,booth_data_11_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_11_T_48 = {_booth_data_11_T_46,_booth_data_11_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [85:0] _GEN_10 = {_booth_data_11_T_48, 22'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_11_T_49 = {{9'd0}, _GEN_10}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_12 = {regs_1[25],regs_1[24],regs_1[23]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_12_T_3 = 3'h1 == look_up_data_12 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_12_T_5 = 3'h2 == look_up_data_12 ? regs_0 : _booth_data_12_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_7 = 3'h3 == look_up_data_12 ? _booth_data_0_T : {{1'd0}, _booth_data_12_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_9 = 3'h4 == look_up_data_12 ? _booth_data_0_T_1 : _booth_data_12_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_11 = 3'h5 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_13 = 3'h6 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_15 = 3'h7 == look_up_data_12 ? 69'h0 : _booth_data_12_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_12_lo_lo = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_12_lo = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[
    33],booth_data_12_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_12_T_46 = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[
    33],booth_data_12_lo_lo,booth_data_12_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_12_T_48 = {_booth_data_12_T_46,_booth_data_12_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [87:0] _GEN_11 = {_booth_data_12_T_48, 24'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_12_T_49 = {{7'd0}, _GEN_11}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_13 = {regs_1[27],regs_1[26],regs_1[25]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_13_T_3 = 3'h1 == look_up_data_13 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_13_T_5 = 3'h2 == look_up_data_13 ? regs_0 : _booth_data_13_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_7 = 3'h3 == look_up_data_13 ? _booth_data_0_T : {{1'd0}, _booth_data_13_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_9 = 3'h4 == look_up_data_13 ? _booth_data_0_T_1 : _booth_data_13_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_11 = 3'h5 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_13 = 3'h6 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_15 = 3'h7 == look_up_data_13 ? 69'h0 : _booth_data_13_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_13_lo_lo = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_13_lo = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[
    33],booth_data_13_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_13_T_46 = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[
    33],booth_data_13_lo_lo,booth_data_13_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_13_T_48 = {_booth_data_13_T_46,_booth_data_13_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [89:0] _GEN_12 = {_booth_data_13_T_48, 26'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_13_T_49 = {{5'd0}, _GEN_12}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_14 = {regs_1[29],regs_1[28],regs_1[27]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_14_T_3 = 3'h1 == look_up_data_14 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_14_T_5 = 3'h2 == look_up_data_14 ? regs_0 : _booth_data_14_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_7 = 3'h3 == look_up_data_14 ? _booth_data_0_T : {{1'd0}, _booth_data_14_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_9 = 3'h4 == look_up_data_14 ? _booth_data_0_T_1 : _booth_data_14_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_11 = 3'h5 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_13 = 3'h6 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_15 = 3'h7 == look_up_data_14 ? 69'h0 : _booth_data_14_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_14_lo_lo = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_14_lo = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[
    33],booth_data_14_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_14_T_46 = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[
    33],booth_data_14_lo_lo,booth_data_14_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_14_T_48 = {_booth_data_14_T_46,_booth_data_14_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [91:0] _GEN_13 = {_booth_data_14_T_48, 28'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_14_T_49 = {{3'd0}, _GEN_13}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_15 = {regs_1[31],regs_1[30],regs_1[29]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_15_T_3 = 3'h1 == look_up_data_15 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_15_T_5 = 3'h2 == look_up_data_15 ? regs_0 : _booth_data_15_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_7 = 3'h3 == look_up_data_15 ? _booth_data_0_T : {{1'd0}, _booth_data_15_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_9 = 3'h4 == look_up_data_15 ? _booth_data_0_T_1 : _booth_data_15_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_11 = 3'h5 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_13 = 3'h6 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_15 = 3'h7 == look_up_data_15 ? 69'h0 : _booth_data_15_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_15_lo_lo = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_15_lo = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[
    33],booth_data_15_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_15_T_46 = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[
    33],booth_data_15_lo_lo,booth_data_15_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_15_T_48 = {_booth_data_15_T_46,_booth_data_15_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [93:0] _GEN_14 = {_booth_data_15_T_48, 30'h0}; // @[hard_cal.scala 290:19]
  wire [94:0] _booth_data_15_T_49 = {{1'd0}, _GEN_14}; // @[hard_cal.scala 290:19]
  wire [2:0] look_up_data_16 = {regs_1[33],regs_1[32],regs_1[31]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_16_T_3 = 3'h1 == look_up_data_16 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_16_T_5 = 3'h2 == look_up_data_16 ? regs_0 : _booth_data_16_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_7 = 3'h3 == look_up_data_16 ? _booth_data_0_T : {{1'd0}, _booth_data_16_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_9 = 3'h4 == look_up_data_16 ? _booth_data_0_T_1 : _booth_data_16_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_11 = 3'h5 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_13 = 3'h6 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_15 = 3'h7 == look_up_data_16 ? 69'h0 : _booth_data_16_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_16_lo_lo = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_16_lo = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[
    33],booth_data_16_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_16_T_46 = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[
    33],booth_data_16_lo_lo,booth_data_16_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_16_T_48 = {_booth_data_16_T_46,_booth_data_16_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [95:0] _GEN_15 = {_booth_data_16_T_48, 32'h0}; // @[hard_cal.scala 290:19]
  wire [126:0] _booth_data_16_T_49 = {{31'd0}, _GEN_15}; // @[hard_cal.scala 290:19]
  wire [33:0] _x_fu_T_1 = ~io_data_0; // @[hard_cal.scala 295:56]
  wire [33:0] _x_fu_T_3 = _x_fu_T_1 + 34'h1; // @[hard_cal.scala 295:70]
  wire [2:0] _cal_start_T_2 = 3'h7 - 3'h1; // @[hard_cal.scala 302:115]
  wire [5:0] _GEN_16 = {{3'd0}, _cal_start_T_2}; // @[hard_cal.scala 302:81]
  wire  _cal_start_T_4 = counter == _GEN_16 ? 1'h0 : cal_start; // @[hard_cal.scala 302:72]
  ysyx_22040886_wallace_adder_1 cal_module ( // @[hard_cal.scala 300:28]
    .clock(cal_module_clock),
    .reset(cal_module_reset),
    .io_data_in_0(cal_module_io_data_in_0),
    .io_data_in_1(cal_module_io_data_in_1),
    .io_data_in_2(cal_module_io_data_in_2),
    .io_data_in_3(cal_module_io_data_in_3),
    .io_data_in_4(cal_module_io_data_in_4),
    .io_data_in_5(cal_module_io_data_in_5),
    .io_data_in_6(cal_module_io_data_in_6),
    .io_data_in_7(cal_module_io_data_in_7),
    .io_data_in_8(cal_module_io_data_in_8),
    .io_data_in_9(cal_module_io_data_in_9),
    .io_data_in_10(cal_module_io_data_in_10),
    .io_data_in_11(cal_module_io_data_in_11),
    .io_data_in_12(cal_module_io_data_in_12),
    .io_data_in_13(cal_module_io_data_in_13),
    .io_data_in_14(cal_module_io_data_in_14),
    .io_data_in_15(cal_module_io_data_in_15),
    .io_data_in_16(cal_module_io_data_in_16),
    .io_result(cal_module_io_result)
  );
  assign io_result_0 = cal_start ? cal_module_io_result[33:0] : result_reg[33:0]; // @[hard_cal.scala 308:24]
  assign io_Output_valid = counter == _GEN_16; // @[hard_cal.scala 310:34]
  assign cal_module_clock = clock;
  assign cal_module_reset = reset;
  assign cal_module_io_data_in_0 = {{3'd0}, _booth_data_0_T_49}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_1 = {{1'd0}, _booth_data_1_T_49}; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_2 = _booth_data_2_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_3 = _booth_data_3_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_4 = _booth_data_4_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_5 = _booth_data_5_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_6 = _booth_data_6_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_7 = _booth_data_7_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_8 = _booth_data_8_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_9 = _booth_data_9_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_10 = _booth_data_10_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_11 = _booth_data_11_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_12 = _booth_data_12_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_13 = _booth_data_13_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_14 = _booth_data_14_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_15 = _booth_data_15_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  assign cal_module_io_data_in_16 = _booth_data_16_T_49[67:0]; // @[hard_cal.scala 268:26 280:27]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 259:23]
      regs_0 <= 68'h0; // @[hard_cal.scala 259:23]
    end else if (_signed_T) begin // @[hard_cal.scala 294:19]
      regs_0 <= {{34'd0}, io_data_0};
    end
    if (reset) begin // @[hard_cal.scala 259:23]
      regs_1 <= 68'h0; // @[hard_cal.scala 259:23]
    end else if (_signed_T) begin // @[hard_cal.scala 296:19]
      regs_1 <= {{34'd0}, io_data_1};
    end
    if (reset) begin // @[hard_cal.scala 261:26]
      counter <= 6'h0; // @[hard_cal.scala 261:26]
    end else if (cal_start) begin // @[hard_cal.scala 264:19]
      counter <= _counter_T_1;
    end else begin
      counter <= 6'h0;
    end
    if (reset) begin // @[hard_cal.scala 262:28]
      cal_start <= 1'h0; // @[hard_cal.scala 262:28]
    end else begin
      cal_start <= _signed_T | _cal_start_T_4; // @[hard_cal.scala 302:15]
    end
    if (reset) begin // @[hard_cal.scala 266:29]
      result_reg <= 68'h0; // @[hard_cal.scala 266:29]
    end else if (cal_start) begin // @[hard_cal.scala 307:22]
      result_reg <= cal_module_io_result;
    end
    if (reset) begin // @[hard_cal.scala 269:23]
      x_fu <= 68'h0; // @[hard_cal.scala 269:23]
    end else if (_signed_T) begin // @[hard_cal.scala 295:18]
      x_fu <= {{34'd0}, _x_fu_T_3};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  regs_0 = _RAND_0[67:0];
  _RAND_1 = {3{`RANDOM}};
  regs_1 = _RAND_1[67:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {3{`RANDOM}};
  result_reg = _RAND_4[67:0];
  _RAND_5 = {3{`RANDOM}};
  x_fu = _RAND_5[67:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_div_simple(
  input         clock,
  input         reset,
  output [63:0] io_result_0,
  output [63:0] io_result_1,
  input  [63:0] io_data_0,
  input  [63:0] io_data_1,
  input         io_input_valid,
  output        io_Output_valid,
  input         io_signed
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] regs_0; // @[hard_cal.scala 65:23]
  reg [127:0] regs_1; // @[hard_cal.scala 65:23]
  reg [6:0] counter; // @[hard_cal.scala 67:26]
  reg  cal_start; // @[hard_cal.scala 68:28]
  wire  input_ready_to_be = ~cal_start; // @[hard_cal.scala 108:26]
  wire  _cal_start_T = io_input_valid & input_ready_to_be; // @[hard_cal.scala 69:37]
  wire  _cal_start_T_2 = counter == 7'h40 ? 1'h0 : cal_start; // @[hard_cal.scala 69:72]
  wire [6:0] _counter_T_1 = counter + 7'h1; // @[hard_cal.scala 70:39]
  reg [63:0] result_reg; // @[hard_cal.scala 72:29]
  wire [63:0] _data_in_0_T_2 = ~io_data_0; // @[hard_cal.scala 76:59]
  wire [63:0] _data_in_0_T_4 = _data_in_0_T_2 + 64'h1; // @[hard_cal.scala 76:76]
  wire [63:0] data_in_0 = io_signed & io_data_0[63] ? _data_in_0_T_4 : io_data_0; // @[hard_cal.scala 76:17]
  wire [63:0] _data_in_1_T_2 = ~io_data_1; // @[hard_cal.scala 76:59]
  wire [63:0] _data_in_1_T_4 = _data_in_1_T_2 + 64'h1; // @[hard_cal.scala 76:76]
  wire [63:0] data_in_1 = io_signed & io_data_1[63] ? _data_in_1_T_4 : io_data_1; // @[hard_cal.scala 76:17]
  wire [1:0] _T_2 = {io_data_0[63],io_data_1[63]}; // @[Cat.scala 31:58]
  wire  _T_6_1 = 2'h1 == _T_2 ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _T_8_0 = 2'h0 == _T_2 ? 1'h0 : 2'h1 == _T_2 | 2'h2 == _T_2; // @[Mux.scala 81:58]
  wire  _T_8_1 = 2'h0 == _T_2 ? 1'h0 : _T_6_1; // @[Mux.scala 81:58]
  wire  result_sign_0 = io_signed & _T_8_0; // @[hard_cal.scala 79:23]
  wire  result_sign_1 = io_signed & _T_8_1; // @[hard_cal.scala 79:23]
  wire [64:0] _by_divide_num_T_1 = regs_0[127:63]; // @[hard_cal.scala 93:58]
  wire [64:0] _by_divide_num_T_4 = {1'h0,regs_1[63:0]}; // @[hard_cal.scala 93:103]
  wire [64:0] by_divide_num = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 93:65]
  wire  minus_answer = $signed(by_divide_num) >= 65'sh0; // @[hard_cal.scala 94:35]
  wire [64:0] _regs0_to_be_T = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 95:58]
  wire [63:0] _regs0_to_be_T_3 = minus_answer ? _regs0_to_be_T[63:0] : regs_0[126:63]; // @[hard_cal.scala 95:30]
  wire [127:0] regs0_to_be = {_regs0_to_be_T_3,regs_0[62:0],1'h0}; // @[Cat.scala 31:58]
  wire [64:0] _result_reg_T = {result_reg, 1'h0}; // @[hard_cal.scala 99:49]
  wire [63:0] _result_reg_T_2 = {_result_reg_T[63:1],minus_answer}; // @[Cat.scala 31:58]
  wire [63:0] _io_result_0_T = ~_result_reg_T_2; // @[hard_cal.scala 105:38]
  wire [63:0] _io_result_0_T_2 = _io_result_0_T + 64'h1; // @[hard_cal.scala 105:60]
  wire [63:0] _io_result_1_T = ~_regs0_to_be_T_3; // @[hard_cal.scala 105:38]
  wire [63:0] _io_result_1_T_2 = _io_result_1_T + 64'h1; // @[hard_cal.scala 105:60]
  wire [6:0] _io_Output_valid_T_1 = 7'h40 - 7'h1; // @[hard_cal.scala 107:45]
  assign io_result_0 = result_sign_0 ? _io_result_0_T_2 : _result_reg_T_2; // @[hard_cal.scala 105:17]
  assign io_result_1 = result_sign_1 ? _io_result_1_T_2 : _regs0_to_be_T_3; // @[hard_cal.scala 105:17]
  assign io_Output_valid = counter == _io_Output_valid_T_1; // @[hard_cal.scala 107:33]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 65:23]
      regs_0 <= 128'h0; // @[hard_cal.scala 65:23]
    end else if (_cal_start_T) begin // @[hard_cal.scala 96:19]
      regs_0 <= {{64'd0}, data_in_0};
    end else if (cal_start) begin // @[hard_cal.scala 96:70]
      regs_0 <= regs0_to_be;
    end
    if (reset) begin // @[hard_cal.scala 65:23]
      regs_1 <= 128'h0; // @[hard_cal.scala 65:23]
    end else if (_cal_start_T) begin // @[hard_cal.scala 98:19]
      regs_1 <= {{64'd0}, data_in_1};
    end
    if (reset) begin // @[hard_cal.scala 67:26]
      counter <= 7'h0; // @[hard_cal.scala 67:26]
    end else if (cal_start) begin // @[hard_cal.scala 70:19]
      counter <= _counter_T_1;
    end else begin
      counter <= 7'h0;
    end
    if (reset) begin // @[hard_cal.scala 68:28]
      cal_start <= 1'h0; // @[hard_cal.scala 68:28]
    end else begin
      cal_start <= io_input_valid & input_ready_to_be | _cal_start_T_2; // @[hard_cal.scala 69:15]
    end
    if (reset) begin // @[hard_cal.scala 72:29]
      result_reg <= 64'h0; // @[hard_cal.scala 72:29]
    end else if (cal_start) begin // @[hard_cal.scala 99:22]
      result_reg <= _result_reg_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  regs_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  regs_1 = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  result_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_div_simple_1(
  input         clock,
  input         reset,
  output [31:0] io_result_0,
  output [31:0] io_result_1,
  input  [31:0] io_data_0,
  input  [31:0] io_data_1,
  input         io_input_valid,
  output        io_Output_valid,
  input         io_signed
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[hard_cal.scala 65:23]
  reg [63:0] regs_1; // @[hard_cal.scala 65:23]
  reg [5:0] counter; // @[hard_cal.scala 67:26]
  reg  cal_start; // @[hard_cal.scala 68:28]
  wire  input_ready_to_be = ~cal_start; // @[hard_cal.scala 108:26]
  wire  _cal_start_T = io_input_valid & input_ready_to_be; // @[hard_cal.scala 69:37]
  wire  _cal_start_T_2 = counter == 6'h20 ? 1'h0 : cal_start; // @[hard_cal.scala 69:72]
  wire [5:0] _counter_T_1 = counter + 6'h1; // @[hard_cal.scala 70:39]
  reg [31:0] result_reg; // @[hard_cal.scala 72:29]
  wire [31:0] _data_in_0_T_2 = ~io_data_0; // @[hard_cal.scala 76:59]
  wire [31:0] _data_in_0_T_4 = _data_in_0_T_2 + 32'h1; // @[hard_cal.scala 76:76]
  wire [31:0] data_in_0 = io_signed & io_data_0[31] ? _data_in_0_T_4 : io_data_0; // @[hard_cal.scala 76:17]
  wire [31:0] _data_in_1_T_2 = ~io_data_1; // @[hard_cal.scala 76:59]
  wire [31:0] _data_in_1_T_4 = _data_in_1_T_2 + 32'h1; // @[hard_cal.scala 76:76]
  wire [31:0] data_in_1 = io_signed & io_data_1[31] ? _data_in_1_T_4 : io_data_1; // @[hard_cal.scala 76:17]
  wire [1:0] _T_2 = {io_data_0[31],io_data_1[31]}; // @[Cat.scala 31:58]
  wire  _T_6_1 = 2'h1 == _T_2 ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _T_8_0 = 2'h0 == _T_2 ? 1'h0 : 2'h1 == _T_2 | 2'h2 == _T_2; // @[Mux.scala 81:58]
  wire  _T_8_1 = 2'h0 == _T_2 ? 1'h0 : _T_6_1; // @[Mux.scala 81:58]
  wire  result_sign_0 = io_signed & _T_8_0; // @[hard_cal.scala 79:23]
  wire  result_sign_1 = io_signed & _T_8_1; // @[hard_cal.scala 79:23]
  wire [32:0] _by_divide_num_T_1 = regs_0[63:31]; // @[hard_cal.scala 93:58]
  wire [32:0] _by_divide_num_T_4 = {1'h0,regs_1[31:0]}; // @[hard_cal.scala 93:103]
  wire [32:0] by_divide_num = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 93:65]
  wire  minus_answer = $signed(by_divide_num) >= 33'sh0; // @[hard_cal.scala 94:35]
  wire [32:0] _regs0_to_be_T = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 95:58]
  wire [31:0] _regs0_to_be_T_3 = minus_answer ? _regs0_to_be_T[31:0] : regs_0[62:31]; // @[hard_cal.scala 95:30]
  wire [63:0] regs0_to_be = {_regs0_to_be_T_3,regs_0[30:0],1'h0}; // @[Cat.scala 31:58]
  wire [32:0] _result_reg_T = {result_reg, 1'h0}; // @[hard_cal.scala 99:49]
  wire [31:0] _result_reg_T_2 = {_result_reg_T[31:1],minus_answer}; // @[Cat.scala 31:58]
  wire [31:0] _io_result_0_T = ~_result_reg_T_2; // @[hard_cal.scala 105:38]
  wire [31:0] _io_result_0_T_2 = _io_result_0_T + 32'h1; // @[hard_cal.scala 105:60]
  wire [31:0] _io_result_1_T = ~_regs0_to_be_T_3; // @[hard_cal.scala 105:38]
  wire [31:0] _io_result_1_T_2 = _io_result_1_T + 32'h1; // @[hard_cal.scala 105:60]
  wire [5:0] _io_Output_valid_T_1 = 6'h20 - 6'h1; // @[hard_cal.scala 107:45]
  assign io_result_0 = result_sign_0 ? _io_result_0_T_2 : _result_reg_T_2; // @[hard_cal.scala 105:17]
  assign io_result_1 = result_sign_1 ? _io_result_1_T_2 : _regs0_to_be_T_3; // @[hard_cal.scala 105:17]
  assign io_Output_valid = counter == _io_Output_valid_T_1; // @[hard_cal.scala 107:33]
  always @(posedge clock) begin
    if (reset) begin // @[hard_cal.scala 65:23]
      regs_0 <= 64'h0; // @[hard_cal.scala 65:23]
    end else if (_cal_start_T) begin // @[hard_cal.scala 96:19]
      regs_0 <= {{32'd0}, data_in_0};
    end else if (cal_start) begin // @[hard_cal.scala 96:70]
      regs_0 <= regs0_to_be;
    end
    if (reset) begin // @[hard_cal.scala 65:23]
      regs_1 <= 64'h0; // @[hard_cal.scala 65:23]
    end else if (_cal_start_T) begin // @[hard_cal.scala 98:19]
      regs_1 <= {{32'd0}, data_in_1};
    end
    if (reset) begin // @[hard_cal.scala 67:26]
      counter <= 6'h0; // @[hard_cal.scala 67:26]
    end else if (cal_start) begin // @[hard_cal.scala 70:19]
      counter <= _counter_T_1;
    end else begin
      counter <= 6'h0;
    end
    if (reset) begin // @[hard_cal.scala 68:28]
      cal_start <= 1'h0; // @[hard_cal.scala 68:28]
    end else begin
      cal_start <= io_input_valid & input_ready_to_be | _cal_start_T_2; // @[hard_cal.scala 69:15]
    end
    if (reset) begin // @[hard_cal.scala 72:29]
      result_reg <= 32'h0; // @[hard_cal.scala 72:29]
    end else if (cal_start) begin // @[hard_cal.scala 99:22]
      result_reg <= _result_reg_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  result_reg = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_muldiv(
  input         clock,
  input         reset,
  input         io_en,
  input  [23:0] io_ctrl,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_data_out,
  output        io_pending
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  mul_hard_clock; // @[muldiv.scala 356:32]
  wire  mul_hard_reset; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_result_0; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_result_1; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_data_0; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_data_1; // @[muldiv.scala 356:32]
  wire  mul_hard_io_input_valid; // @[muldiv.scala 356:32]
  wire  mul_hard_io_Output_valid; // @[muldiv.scala 356:32]
  wire  mul_hard_1_clock; // @[muldiv.scala 357:39]
  wire  mul_hard_1_reset; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_result_0; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_data_0; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_data_1; // @[muldiv.scala 357:39]
  wire  mul_hard_1_io_input_valid; // @[muldiv.scala 357:39]
  wire  mul_hard_1_io_Output_valid; // @[muldiv.scala 357:39]
  wire  div_simple_clock; // @[muldiv.scala 385:32]
  wire  div_simple_reset; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_result_0; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_result_1; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_data_0; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_data_1; // @[muldiv.scala 385:32]
  wire  div_simple_io_input_valid; // @[muldiv.scala 385:32]
  wire  div_simple_io_Output_valid; // @[muldiv.scala 385:32]
  wire  div_simple_io_signed; // @[muldiv.scala 385:32]
  wire  div_simple_1_clock; // @[muldiv.scala 386:39]
  wire  div_simple_1_reset; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_result_0; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_result_1; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_data_0; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_data_1; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_input_valid; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_Output_valid; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_signed; // @[muldiv.scala 386:39]
  wire [23:0] _cal_mul_T_1 = {{9'd0}, io_ctrl[23:9]}; // @[muldiv.scala 300:48]
  wire [23:0] _cal_mul_T_3 = {{12'd0}, io_ctrl[23:12]}; // @[muldiv.scala 300:71]
  wire [23:0] _cal_mul_T_6 = {{10'd0}, io_ctrl[23:10]}; // @[muldiv.scala 301:20]
  wire  _cal_mul_T_8 = _cal_mul_T_1[0] | _cal_mul_T_3[0] | _cal_mul_T_6[0]; // @[muldiv.scala 300:87]
  wire [23:0] _cal_mul_T_9 = {{11'd0}, io_ctrl[23:11]}; // @[muldiv.scala 301:46]
  wire  _cal_mul_T_11 = _cal_mul_T_8 | _cal_mul_T_9[0]; // @[muldiv.scala 301:36]
  wire  cal_mul = io_en & _cal_mul_T_11; // @[muldiv.scala 300:34]
  wire [23:0] _cal_div_T_1 = {{1'd0}, io_ctrl[23:1]}; // @[muldiv.scala 302:48]
  wire [23:0] _cal_div_T_6 = {{3'd0}, io_ctrl[23:3]}; // @[muldiv.scala 303:21]
  wire  _cal_div_T_8 = _cal_div_T_1[0] | io_ctrl[0] | _cal_div_T_6[0]; // @[muldiv.scala 302:85]
  wire [23:0] _cal_div_T_9 = {{2'd0}, io_ctrl[23:2]}; // @[muldiv.scala 303:45]
  wire  _cal_div_T_11 = _cal_div_T_8 | _cal_div_T_9[0]; // @[muldiv.scala 303:35]
  wire  cal_div = io_en & _cal_div_T_11; // @[muldiv.scala 302:34]
  wire [23:0] _cal_divw_T_1 = {{4'd0}, io_ctrl[23:4]}; // @[muldiv.scala 304:44]
  wire [23:0] _cal_divw_T_3 = {{5'd0}, io_ctrl[23:5]}; // @[muldiv.scala 304:69]
  wire [23:0] _cal_divw_T_6 = {{6'd0}, io_ctrl[23:6]}; // @[muldiv.scala 304:99]
  wire [23:0] _cal_divw_T_9 = {{7'd0}, io_ctrl[23:7]}; // @[muldiv.scala 304:125]
  wire  cal_divw = io_en & (_cal_divw_T_1[0] | _cal_divw_T_3[0] | _cal_divw_T_6[0] | _cal_divw_T_9[0]); // @[muldiv.scala 304:33]
  wire [23:0] _cal_mulw_T_1 = {{8'd0}, io_ctrl[23:8]}; // @[muldiv.scala 305:45]
  wire  cal_mulw = io_en & _cal_mulw_T_1[0]; // @[muldiv.scala 305:33]
  reg [3:0] work_state; // @[muldiv.scala 308:30]
  reg [23:0] ctrl_data; // @[muldiv.scala 315:28]
  wire  _work_state_T = work_state == 4'h0; // @[muldiv.scala 317:34]
  wire  _work_state_T_1 = cal_mul & work_state == 4'h0; // @[muldiv.scala 317:20]
  wire  _work_state_T_3 = cal_mulw & _work_state_T; // @[muldiv.scala 318:20]
  wire  _work_state_T_5 = cal_div & _work_state_T; // @[muldiv.scala 319:20]
  wire  _work_state_T_7 = cal_divw & _work_state_T; // @[muldiv.scala 320:20]
  wire  _work_state_T_8 = work_state == 4'h1; // @[muldiv.scala 321:37]
  wire  _work_state_T_9 = work_state == 4'h2; // @[muldiv.scala 321:69]
  wire  _cal_end_mul_T_1 = _work_state_T_8 & mul_hard_io_Output_valid; // @[muldiv.scala 368:43]
  wire  _cal_end_mul_T_3 = _work_state_T_9 & mul_hard_1_io_Output_valid; // @[muldiv.scala 369:44]
  wire  cal_end_mul = _cal_end_mul_T_1 | _cal_end_mul_T_3; // @[Mux.scala 101:16]
  wire  _work_state_T_11 = cal_end_mul & (work_state == 4'h1 | work_state == 4'h2); // @[muldiv.scala 321:22]
  wire  _work_state_T_12 = work_state == 4'h3; // @[muldiv.scala 322:38]
  wire  _work_state_T_13 = work_state == 4'h5; // @[muldiv.scala 322:70]
  wire  _cal_end_div_T_1 = _work_state_T_12 & div_simple_io_Output_valid; // @[muldiv.scala 397:43]
  wire  _cal_end_div_T_3 = _work_state_T_13 & div_simple_1_io_Output_valid; // @[muldiv.scala 398:44]
  wire  cal_end_div = _cal_end_div_T_1 | _cal_end_div_T_3; // @[Mux.scala 101:16]
  wire  _work_state_T_15 = cal_end_div & (work_state == 4'h3 | work_state == 4'h5); // @[muldiv.scala 322:23]
  wire  _work_state_T_16 = work_state == 4'h4; // @[muldiv.scala 323:21]
  wire [3:0] _work_state_T_17 = _work_state_T_16 ? 4'h0 : work_state; // @[Mux.scala 101:16]
  wire [3:0] _work_state_T_18 = _work_state_T_15 ? 4'h4 : _work_state_T_17; // @[Mux.scala 101:16]
  wire [3:0] _work_state_T_19 = _work_state_T_11 ? 4'h4 : _work_state_T_18; // @[Mux.scala 101:16]
  wire [3:0] _work_state_T_20 = _work_state_T_7 ? 4'h5 : _work_state_T_19; // @[Mux.scala 101:16]
  wire  cal_signed = _cal_mul_T_1[0] | _cal_mul_T_6[0] | _cal_mulw_T_1[0] | _cal_mul_T_3[0]; // @[muldiv.scala 358:95]
  wire [65:0] _T_3 = {2'h3,io_in1}; // @[Cat.scala 31:58]
  wire [65:0] _T_5 = {2'h0,io_in1}; // @[Cat.scala 31:58]
  wire [65:0] _T_6 = io_in1[63] ? _T_3 : _T_5; // @[macros.scala 436:8]
  wire [64:0] _T_8 = {1'h0,io_in1}; // @[Cat.scala 31:58]
  wire [65:0] _T_13 = {2'h3,io_in2}; // @[Cat.scala 31:58]
  wire [65:0] _T_15 = {2'h0,io_in2}; // @[Cat.scala 31:58]
  wire [65:0] _T_16 = io_in2[63] ? _T_13 : _T_15; // @[macros.scala 436:8]
  wire [64:0] _T_18 = {1'h0,io_in2}; // @[Cat.scala 31:58]
  wire [33:0] _T_24 = {2'h3,io_in1[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_26 = {2'h0,io_in1[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_27 = io_in1[31] ? _T_24 : _T_26; // @[macros.scala 436:8]
  wire [32:0] _T_30 = {1'h0,io_in1[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_36 = {2'h3,io_in2[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_38 = {2'h0,io_in2[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_39 = io_in2[31] ? _T_36 : _T_38; // @[macros.scala 436:8]
  wire [32:0] _T_42 = {1'h0,io_in2[31:0]}; // @[Cat.scala 31:58]
  wire [131:0] final_result = {mul_hard_io_result_1,mul_hard_io_result_0}; // @[Cat.scala 31:58]
  reg [63:0] mul_cal_reg; // @[muldiv.scala 372:34]
  wire [23:0] _access_mul_result_T = {{9'd0}, ctrl_data[23:9]}; // @[muldiv.scala 374:30]
  wire [23:0] _access_mul_result_T_3 = {{10'd0}, ctrl_data[23:10]}; // @[muldiv.scala 375:30]
  wire [23:0] _access_mul_result_T_6 = {{11'd0}, ctrl_data[23:11]}; // @[muldiv.scala 376:30]
  wire [23:0] _access_mul_result_T_9 = {{12'd0}, ctrl_data[23:12]}; // @[muldiv.scala 377:30]
  wire [23:0] _access_mul_result_T_12 = {{8'd0}, ctrl_data[23:8]}; // @[muldiv.scala 378:30]
  wire [7:0] access_mul_result_lo_lo = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31]
    ,mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_mul_result_lo = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],access_mul_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_mul_result_T_47 = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31
    ],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],access_mul_result_lo_lo,access_mul_result_lo}; // @[Cat.scala 31:58]
  wire [63:0] _access_mul_result_T_49 = {_access_mul_result_T_47,mul_hard_1_io_result_0[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _access_mul_result_T_50 = _access_mul_result_T[0] ? final_result[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_51 = _access_mul_result_T_3[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_52 = _access_mul_result_T_6[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_53 = _access_mul_result_T_9[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_54 = _access_mul_result_T_12[0] ? _access_mul_result_T_49 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_55 = _access_mul_result_T_50 | _access_mul_result_T_51; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_56 = _access_mul_result_T_55 | _access_mul_result_T_52; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_57 = _access_mul_result_T_56 | _access_mul_result_T_53; // @[Mux.scala 27:73]
  wire [63:0] access_mul_result = _access_mul_result_T_57 | _access_mul_result_T_54; // @[Mux.scala 27:73]
  wire [63:0] cal_mul_result = cal_end_mul ? access_mul_result : mul_cal_reg; // @[muldiv.scala 380:30]
  reg [63:0] div_cal_reg; // @[muldiv.scala 400:34]
  wire [23:0] _access_div_result_T = {{1'd0}, ctrl_data[23:1]}; // @[muldiv.scala 402:30]
  wire [23:0] _access_div_result_T_4 = {{3'd0}, ctrl_data[23:3]}; // @[muldiv.scala 404:30]
  wire [23:0] _access_div_result_T_6 = {{2'd0}, ctrl_data[23:2]}; // @[muldiv.scala 405:30]
  wire [23:0] _access_div_result_T_8 = {{4'd0}, ctrl_data[23:4]}; // @[muldiv.scala 406:30]
  wire [7:0] access_div_result_lo_lo = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_div_result_lo = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0
    [31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0
    [31],div_simple_1_io_result_0[31],access_div_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_42 = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],access_div_result_lo_lo,access_div_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_43 = div_simple_1_io_result_0; // @[macros.scala 440:65]
  wire [63:0] _access_div_result_T_44 = {_access_div_result_T_42,_access_div_result_T_43}; // @[Cat.scala 31:58]
  wire [23:0] _access_div_result_T_45 = {{5'd0}, ctrl_data[23:5]}; // @[muldiv.scala 407:30]
  wire [23:0] _access_div_result_T_82 = {{6'd0}, ctrl_data[23:6]}; // @[muldiv.scala 408:30]
  wire [7:0] access_div_result_lo_lo_2 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_div_result_lo_2 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],access_div_result_lo_lo_2}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_116 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],access_div_result_lo_lo_2,access_div_result_lo_2}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_117 = div_simple_1_io_result_1; // @[macros.scala 440:65]
  wire [63:0] _access_div_result_T_118 = {_access_div_result_T_116,_access_div_result_T_117}; // @[Cat.scala 31:58]
  wire [23:0] _access_div_result_T_119 = {{7'd0}, ctrl_data[23:7]}; // @[muldiv.scala 409:30]
  wire [63:0] _access_div_result_T_156 = _access_div_result_T[0] ? div_simple_io_result_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_157 = ctrl_data[0] ? div_simple_io_result_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_158 = _access_div_result_T_4[0] ? div_simple_io_result_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_159 = _access_div_result_T_6[0] ? div_simple_io_result_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_160 = _access_div_result_T_8[0] ? _access_div_result_T_44 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_161 = _access_div_result_T_45[0] ? _access_div_result_T_44 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_162 = _access_div_result_T_82[0] ? _access_div_result_T_118 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_163 = _access_div_result_T_119[0] ? _access_div_result_T_118 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_164 = _access_div_result_T_156 | _access_div_result_T_157; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_165 = _access_div_result_T_164 | _access_div_result_T_158; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_166 = _access_div_result_T_165 | _access_div_result_T_159; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_167 = _access_div_result_T_166 | _access_div_result_T_160; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_168 = _access_div_result_T_167 | _access_div_result_T_161; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_169 = _access_div_result_T_168 | _access_div_result_T_162; // @[Mux.scala 27:73]
  wire [63:0] access_div_result = _access_div_result_T_169 | _access_div_result_T_163; // @[Mux.scala 27:73]
  wire [63:0] cal_div_result = cal_end_div ? access_div_result : div_cal_reg; // @[muldiv.scala 411:30]
  wire [63:0] _io_data_out_T_26 = _cal_div_T_1[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_27 = io_ctrl[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_28 = _cal_divw_T_1[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_29 = _cal_divw_T_3[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_30 = _cal_div_T_6[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_31 = _cal_div_T_9[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_32 = _cal_divw_T_6[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_33 = _cal_divw_T_9[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_34 = _cal_mul_T_1[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_35 = _cal_mulw_T_1[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_36 = _cal_mul_T_6[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_37 = _cal_mul_T_9[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_38 = _cal_mul_T_3[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_39 = _io_data_out_T_26 | _io_data_out_T_27; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_40 = _io_data_out_T_39 | _io_data_out_T_28; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_41 = _io_data_out_T_40 | _io_data_out_T_29; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_42 = _io_data_out_T_41 | _io_data_out_T_30; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_43 = _io_data_out_T_42 | _io_data_out_T_31; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_44 = _io_data_out_T_43 | _io_data_out_T_32; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_45 = _io_data_out_T_44 | _io_data_out_T_33; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_46 = _io_data_out_T_45 | _io_data_out_T_34; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_47 = _io_data_out_T_46 | _io_data_out_T_35; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_48 = _io_data_out_T_47 | _io_data_out_T_36; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_49 = _io_data_out_T_48 | _io_data_out_T_37; // @[Mux.scala 27:73]
  ysyx_22040886_mul_hard mul_hard ( // @[muldiv.scala 356:32]
    .clock(mul_hard_clock),
    .reset(mul_hard_reset),
    .io_result_0(mul_hard_io_result_0),
    .io_result_1(mul_hard_io_result_1),
    .io_data_0(mul_hard_io_data_0),
    .io_data_1(mul_hard_io_data_1),
    .io_input_valid(mul_hard_io_input_valid),
    .io_Output_valid(mul_hard_io_Output_valid)
  );
  ysyx_22040886_mul_hard_1 mul_hard_1 ( // @[muldiv.scala 357:39]
    .clock(mul_hard_1_clock),
    .reset(mul_hard_1_reset),
    .io_result_0(mul_hard_1_io_result_0),
    .io_data_0(mul_hard_1_io_data_0),
    .io_data_1(mul_hard_1_io_data_1),
    .io_input_valid(mul_hard_1_io_input_valid),
    .io_Output_valid(mul_hard_1_io_Output_valid)
  );
  ysyx_22040886_div_simple div_simple ( // @[muldiv.scala 385:32]
    .clock(div_simple_clock),
    .reset(div_simple_reset),
    .io_result_0(div_simple_io_result_0),
    .io_result_1(div_simple_io_result_1),
    .io_data_0(div_simple_io_data_0),
    .io_data_1(div_simple_io_data_1),
    .io_input_valid(div_simple_io_input_valid),
    .io_Output_valid(div_simple_io_Output_valid),
    .io_signed(div_simple_io_signed)
  );
  ysyx_22040886_div_simple_1 div_simple_1 ( // @[muldiv.scala 386:39]
    .clock(div_simple_1_clock),
    .reset(div_simple_1_reset),
    .io_result_0(div_simple_1_io_result_0),
    .io_result_1(div_simple_1_io_result_1),
    .io_data_0(div_simple_1_io_data_0),
    .io_data_1(div_simple_1_io_data_1),
    .io_input_valid(div_simple_1_io_input_valid),
    .io_Output_valid(div_simple_1_io_Output_valid),
    .io_signed(div_simple_1_io_signed)
  );
  assign io_data_out = _io_data_out_T_49 | _io_data_out_T_38; // @[Mux.scala 27:73]
  assign io_pending = work_state != 4'h0 & work_state != 4'h4 | _work_state_T & (cal_mul | cal_mulw | cal_div | cal_divw
    ); // @[muldiv.scala 455:79]
  assign mul_hard_clock = clock;
  assign mul_hard_reset = reset;
  assign mul_hard_io_data_0 = cal_signed ? _T_6 : {{1'd0}, _T_8}; // @[muldiv.scala 361:34]
  assign mul_hard_io_data_1 = cal_signed ? _T_16 : {{1'd0}, _T_18}; // @[muldiv.scala 362:34]
  assign mul_hard_io_input_valid = _work_state_T & cal_mul; // @[muldiv.scala 365:66]
  assign mul_hard_1_clock = clock;
  assign mul_hard_1_reset = reset;
  assign mul_hard_1_io_data_0 = cal_signed ? _T_27 : {{1'd0}, _T_30}; // @[muldiv.scala 363:41]
  assign mul_hard_1_io_data_1 = cal_signed ? _T_39 : {{1'd0}, _T_42}; // @[muldiv.scala 364:41]
  assign mul_hard_1_io_input_valid = _work_state_T & cal_mulw; // @[muldiv.scala 366:72]
  assign div_simple_clock = clock;
  assign div_simple_reset = reset;
  assign div_simple_io_data_0 = io_in1; // @[muldiv.scala 390:28]
  assign div_simple_io_data_1 = io_in2; // @[muldiv.scala 391:28]
  assign div_simple_io_input_valid = _work_state_T & cal_div; // @[muldiv.scala 394:66]
  assign div_simple_io_signed = _cal_div_T_1[0] | _cal_divw_T_1[0] | _cal_div_T_6[0] | _cal_divw_T_6[0]; // @[muldiv.scala 387:96]
  assign div_simple_1_clock = clock;
  assign div_simple_1_reset = reset;
  assign div_simple_1_io_data_0 = io_in1[31:0]; // @[muldiv.scala 392:35]
  assign div_simple_1_io_data_1 = io_in2[31:0]; // @[muldiv.scala 393:35]
  assign div_simple_1_io_input_valid = _work_state_T & cal_divw; // @[muldiv.scala 395:72]
  assign div_simple_1_io_signed = _cal_div_T_1[0] | _cal_divw_T_1[0] | _cal_div_T_6[0] | _cal_divw_T_6[0]; // @[muldiv.scala 387:96]
  always @(posedge clock) begin
    if (reset) begin // @[muldiv.scala 308:30]
      work_state <= 4'h0; // @[muldiv.scala 308:30]
    end else if (_work_state_T_1) begin // @[Mux.scala 101:16]
      work_state <= 4'h1;
    end else if (_work_state_T_3) begin // @[Mux.scala 101:16]
      work_state <= 4'h2;
    end else if (_work_state_T_5) begin // @[Mux.scala 101:16]
      work_state <= 4'h3;
    end else begin
      work_state <= _work_state_T_20;
    end
    if (reset) begin // @[muldiv.scala 315:28]
      ctrl_data <= 24'h0; // @[muldiv.scala 315:28]
    end else if (_work_state_T) begin // @[muldiv.scala 325:22]
      ctrl_data <= io_ctrl;
    end
    if (reset) begin // @[muldiv.scala 372:34]
      mul_cal_reg <= 64'h0; // @[muldiv.scala 372:34]
    end else if (cal_end_mul) begin // @[muldiv.scala 380:30]
      mul_cal_reg <= access_mul_result;
    end
    if (reset) begin // @[muldiv.scala 400:34]
      div_cal_reg <= 64'h0; // @[muldiv.scala 400:34]
    end else if (cal_end_div) begin // @[muldiv.scala 411:30]
      div_cal_reg <= access_div_result;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  work_state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  ctrl_data = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  mul_cal_reg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  div_cal_reg = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_regfile(
  input         clock,
  input         reset,
  input  [4:0]  io_A1,
  input  [4:0]  io_A2,
  input         io_WE3,
  input  [4:0]  io_A3,
  input  [63:0] io_WD3,
  output [63:0] io_RD1,
  output [63:0] io_RD2
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[regfile.scala 24:23]
  reg [63:0] regs_1; // @[regfile.scala 24:23]
  reg [63:0] regs_2; // @[regfile.scala 24:23]
  reg [63:0] regs_3; // @[regfile.scala 24:23]
  reg [63:0] regs_4; // @[regfile.scala 24:23]
  reg [63:0] regs_5; // @[regfile.scala 24:23]
  reg [63:0] regs_6; // @[regfile.scala 24:23]
  reg [63:0] regs_7; // @[regfile.scala 24:23]
  reg [63:0] regs_8; // @[regfile.scala 24:23]
  reg [63:0] regs_9; // @[regfile.scala 24:23]
  reg [63:0] regs_10; // @[regfile.scala 24:23]
  reg [63:0] regs_11; // @[regfile.scala 24:23]
  reg [63:0] regs_12; // @[regfile.scala 24:23]
  reg [63:0] regs_13; // @[regfile.scala 24:23]
  reg [63:0] regs_14; // @[regfile.scala 24:23]
  reg [63:0] regs_15; // @[regfile.scala 24:23]
  reg [63:0] regs_16; // @[regfile.scala 24:23]
  reg [63:0] regs_17; // @[regfile.scala 24:23]
  reg [63:0] regs_18; // @[regfile.scala 24:23]
  reg [63:0] regs_19; // @[regfile.scala 24:23]
  reg [63:0] regs_20; // @[regfile.scala 24:23]
  reg [63:0] regs_21; // @[regfile.scala 24:23]
  reg [63:0] regs_22; // @[regfile.scala 24:23]
  reg [63:0] regs_23; // @[regfile.scala 24:23]
  reg [63:0] regs_24; // @[regfile.scala 24:23]
  reg [63:0] regs_25; // @[regfile.scala 24:23]
  reg [63:0] regs_26; // @[regfile.scala 24:23]
  reg [63:0] regs_27; // @[regfile.scala 24:23]
  reg [63:0] regs_28; // @[regfile.scala 24:23]
  reg [63:0] regs_29; // @[regfile.scala 24:23]
  reg [63:0] regs_30; // @[regfile.scala 24:23]
  reg [63:0] regs_31; // @[regfile.scala 24:23]
  wire [63:0] _GEN_1 = 5'h1 == io_A3 ? regs_1 : regs_0; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_2 = 5'h2 == io_A3 ? regs_2 : _GEN_1; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_3 = 5'h3 == io_A3 ? regs_3 : _GEN_2; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_4 = 5'h4 == io_A3 ? regs_4 : _GEN_3; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_5 = 5'h5 == io_A3 ? regs_5 : _GEN_4; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_6 = 5'h6 == io_A3 ? regs_6 : _GEN_5; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_7 = 5'h7 == io_A3 ? regs_7 : _GEN_6; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_8 = 5'h8 == io_A3 ? regs_8 : _GEN_7; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_9 = 5'h9 == io_A3 ? regs_9 : _GEN_8; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_10 = 5'ha == io_A3 ? regs_10 : _GEN_9; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_11 = 5'hb == io_A3 ? regs_11 : _GEN_10; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_12 = 5'hc == io_A3 ? regs_12 : _GEN_11; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_13 = 5'hd == io_A3 ? regs_13 : _GEN_12; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_14 = 5'he == io_A3 ? regs_14 : _GEN_13; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_15 = 5'hf == io_A3 ? regs_15 : _GEN_14; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_16 = 5'h10 == io_A3 ? regs_16 : _GEN_15; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_17 = 5'h11 == io_A3 ? regs_17 : _GEN_16; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_18 = 5'h12 == io_A3 ? regs_18 : _GEN_17; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_19 = 5'h13 == io_A3 ? regs_19 : _GEN_18; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_20 = 5'h14 == io_A3 ? regs_20 : _GEN_19; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_21 = 5'h15 == io_A3 ? regs_21 : _GEN_20; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_22 = 5'h16 == io_A3 ? regs_22 : _GEN_21; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_23 = 5'h17 == io_A3 ? regs_23 : _GEN_22; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_24 = 5'h18 == io_A3 ? regs_24 : _GEN_23; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_25 = 5'h19 == io_A3 ? regs_25 : _GEN_24; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_26 = 5'h1a == io_A3 ? regs_26 : _GEN_25; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_27 = 5'h1b == io_A3 ? regs_27 : _GEN_26; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_28 = 5'h1c == io_A3 ? regs_28 : _GEN_27; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_29 = 5'h1d == io_A3 ? regs_29 : _GEN_28; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_30 = 5'h1e == io_A3 ? regs_30 : _GEN_29; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_65 = 5'h1 == io_A1 ? regs_1 : regs_0; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_66 = 5'h2 == io_A1 ? regs_2 : _GEN_65; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_67 = 5'h3 == io_A1 ? regs_3 : _GEN_66; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_68 = 5'h4 == io_A1 ? regs_4 : _GEN_67; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_69 = 5'h5 == io_A1 ? regs_5 : _GEN_68; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_70 = 5'h6 == io_A1 ? regs_6 : _GEN_69; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_71 = 5'h7 == io_A1 ? regs_7 : _GEN_70; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_72 = 5'h8 == io_A1 ? regs_8 : _GEN_71; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_73 = 5'h9 == io_A1 ? regs_9 : _GEN_72; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_74 = 5'ha == io_A1 ? regs_10 : _GEN_73; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_75 = 5'hb == io_A1 ? regs_11 : _GEN_74; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_76 = 5'hc == io_A1 ? regs_12 : _GEN_75; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_77 = 5'hd == io_A1 ? regs_13 : _GEN_76; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_78 = 5'he == io_A1 ? regs_14 : _GEN_77; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_79 = 5'hf == io_A1 ? regs_15 : _GEN_78; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_80 = 5'h10 == io_A1 ? regs_16 : _GEN_79; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_81 = 5'h11 == io_A1 ? regs_17 : _GEN_80; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_82 = 5'h12 == io_A1 ? regs_18 : _GEN_81; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_83 = 5'h13 == io_A1 ? regs_19 : _GEN_82; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_84 = 5'h14 == io_A1 ? regs_20 : _GEN_83; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_85 = 5'h15 == io_A1 ? regs_21 : _GEN_84; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_86 = 5'h16 == io_A1 ? regs_22 : _GEN_85; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_87 = 5'h17 == io_A1 ? regs_23 : _GEN_86; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_88 = 5'h18 == io_A1 ? regs_24 : _GEN_87; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_89 = 5'h19 == io_A1 ? regs_25 : _GEN_88; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_90 = 5'h1a == io_A1 ? regs_26 : _GEN_89; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_91 = 5'h1b == io_A1 ? regs_27 : _GEN_90; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_92 = 5'h1c == io_A1 ? regs_28 : _GEN_91; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_93 = 5'h1d == io_A1 ? regs_29 : _GEN_92; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_94 = 5'h1e == io_A1 ? regs_30 : _GEN_93; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_95 = 5'h1f == io_A1 ? regs_31 : _GEN_94; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_97 = 5'h1 == io_A2 ? regs_1 : regs_0; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_98 = 5'h2 == io_A2 ? regs_2 : _GEN_97; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_99 = 5'h3 == io_A2 ? regs_3 : _GEN_98; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_100 = 5'h4 == io_A2 ? regs_4 : _GEN_99; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_101 = 5'h5 == io_A2 ? regs_5 : _GEN_100; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_102 = 5'h6 == io_A2 ? regs_6 : _GEN_101; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_103 = 5'h7 == io_A2 ? regs_7 : _GEN_102; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_104 = 5'h8 == io_A2 ? regs_8 : _GEN_103; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_105 = 5'h9 == io_A2 ? regs_9 : _GEN_104; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_106 = 5'ha == io_A2 ? regs_10 : _GEN_105; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_107 = 5'hb == io_A2 ? regs_11 : _GEN_106; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_108 = 5'hc == io_A2 ? regs_12 : _GEN_107; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_109 = 5'hd == io_A2 ? regs_13 : _GEN_108; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_110 = 5'he == io_A2 ? regs_14 : _GEN_109; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_111 = 5'hf == io_A2 ? regs_15 : _GEN_110; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_112 = 5'h10 == io_A2 ? regs_16 : _GEN_111; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_113 = 5'h11 == io_A2 ? regs_17 : _GEN_112; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_114 = 5'h12 == io_A2 ? regs_18 : _GEN_113; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_115 = 5'h13 == io_A2 ? regs_19 : _GEN_114; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_116 = 5'h14 == io_A2 ? regs_20 : _GEN_115; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_117 = 5'h15 == io_A2 ? regs_21 : _GEN_116; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_118 = 5'h16 == io_A2 ? regs_22 : _GEN_117; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_119 = 5'h17 == io_A2 ? regs_23 : _GEN_118; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_120 = 5'h18 == io_A2 ? regs_24 : _GEN_119; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_121 = 5'h19 == io_A2 ? regs_25 : _GEN_120; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_122 = 5'h1a == io_A2 ? regs_26 : _GEN_121; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_123 = 5'h1b == io_A2 ? regs_27 : _GEN_122; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_124 = 5'h1c == io_A2 ? regs_28 : _GEN_123; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_125 = 5'h1d == io_A2 ? regs_29 : _GEN_124; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_126 = 5'h1e == io_A2 ? regs_30 : _GEN_125; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_127 = 5'h1f == io_A2 ? regs_31 : _GEN_126; // @[regfile.scala 32:{19,19}]
  assign io_RD1 = io_WE3 & io_A1 == io_A3 & io_A1 != 5'h0 ? io_WD3 : _GEN_95; // @[regfile.scala 31:19]
  assign io_RD2 = io_WE3 & io_A2 == io_A3 & io_A2 != 5'h0 ? io_WD3 : _GEN_127; // @[regfile.scala 32:19]
  always @(posedge clock) begin
    if (reset) begin // @[regfile.scala 24:23]
      regs_0 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h0 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_0 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_0 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_0 <= _GEN_30;
      end
    end else begin
      regs_0 <= 64'h0; // @[regfile.scala 25:13]
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_1 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_1 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_1 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_1 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_2 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h2 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_2 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_2 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_2 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_3 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h3 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_3 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_3 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_3 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_4 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h4 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_4 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_4 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_4 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_5 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h5 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_5 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_5 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_5 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_6 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h6 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_6 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_6 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_6 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_7 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h7 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_7 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_7 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_7 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_8 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h8 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_8 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_8 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_8 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_9 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h9 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_9 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_9 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_9 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_10 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'ha == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_10 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_10 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_10 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_11 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'hb == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_11 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_11 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_11 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_12 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'hc == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_12 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_12 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_12 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_13 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'hd == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_13 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_13 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_13 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_14 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'he == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_14 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_14 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_14 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_15 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'hf == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_15 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_15 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_15 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_16 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h10 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_16 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_16 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_16 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_17 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h11 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_17 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_17 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_17 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_18 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h12 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_18 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_18 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_18 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_19 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h13 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_19 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_19 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_19 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_20 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h14 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_20 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_20 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_20 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_21 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h15 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_21 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_21 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_21 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_22 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h16 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_22 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_22 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_22 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_23 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h17 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_23 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_23 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_23 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_24 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h18 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_24 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_24 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_24 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_25 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h19 == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_25 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_25 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_25 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_26 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1a == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_26 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_26 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_26 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_27 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1b == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_27 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_27 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_27 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_28 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1c == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_28 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_28 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_28 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_29 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1d == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_29 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_29 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_29 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_30 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1e == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_30 <= io_WD3;
      end else if (5'h1f == io_A3) begin // @[regfile.scala 26:23]
        regs_30 <= regs_31; // @[regfile.scala 26:23]
      end else begin
        regs_30 <= _GEN_30;
      end
    end
    if (reset) begin // @[regfile.scala 24:23]
      regs_31 <= 64'h0; // @[regfile.scala 24:23]
    end else if (5'h1f == io_A3) begin // @[regfile.scala 26:17]
      if (io_WE3 & io_A3 != 5'h0) begin // @[regfile.scala 26:23]
        regs_31 <= io_WD3;
      end else if (!(5'h1f == io_A3)) begin // @[regfile.scala 26:23]
        regs_31 <= _GEN_30;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_Look_up_table_read_first_with_bundle(
  input         clock,
  input         reset,
  input  [3:0]  io_ar_addr,
  input  [3:0]  io_aw_addr,
  input         io_write,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input  [31:0] io_in_pre_pc_target,
  input  [6:0]  io_in_pre_lookup_data,
  input  [3:0]  io_in_pre_hashcode,
  input  [1:0]  io_in_pre_pht,
  input  [6:0]  io_in_pre_bht,
  input         io_in_pre_decoder_branchD_flag,
  input         io_in_pre_decoder_jump,
  input  [5:0]  io_in_pre_decoder_branchdata,
  input         io_in_pre_decoder_jr,
  input         io_in_true_branch_state,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output [1:0]  io_out_exception_type,
  output [31:0] io_out_pre_pc_target,
  output [6:0]  io_out_pre_lookup_data,
  output [3:0]  io_out_pre_hashcode,
  output [1:0]  io_out_pre_pht,
  output [6:0]  io_out_pre_bht,
  output        io_out_pre_decoder_branchD_flag,
  output        io_out_pre_decoder_jump,
  output [5:0]  io_out_pre_decoder_branchdata,
  output        io_out_pre_decoder_jr,
  output        io_out_true_branch_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] btb_0_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_0_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_0_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_0_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_0_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_0_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_0_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_0_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_1_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_1_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_1_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_1_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_1_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_1_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_1_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_1_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_1_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_2_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_2_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_2_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_2_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_2_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_2_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_2_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_2_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_2_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_3_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_3_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_3_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_3_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_3_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_3_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_3_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_3_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_3_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_4_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_4_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_4_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_4_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_4_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_4_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_4_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_4_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_4_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_5_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_5_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_5_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_5_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_5_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_5_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_5_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_5_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_5_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_6_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_6_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_6_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_6_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_6_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_6_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_6_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_6_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_6_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_7_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_7_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_7_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_7_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_7_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_7_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_7_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_7_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_7_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_8_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_8_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_8_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_8_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_8_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_8_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_8_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_8_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_8_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_9_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_9_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_9_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_9_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_9_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_9_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_9_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_9_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_9_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_10_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_10_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_10_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_10_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_10_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_10_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_10_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_10_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_10_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_11_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_11_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_11_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_11_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_11_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_11_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_11_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_11_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_11_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_12_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_12_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_12_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_12_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_12_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_12_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_12_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_12_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_12_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_13_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_13_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_13_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_13_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_13_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_13_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_13_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_13_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_13_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_14_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_14_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_14_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_14_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_14_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_14_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_14_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_14_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_14_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_15_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_15_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_15_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_15_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_15_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_15_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_15_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_15_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_true_branch_state; // @[ports_lookup_table.scala 105:22]
  wire  _GEN_1 = 4'h1 == io_ar_addr ? btb_1_true_branch_state : btb_0_true_branch_state; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_2 = 4'h2 == io_ar_addr ? btb_2_true_branch_state : _GEN_1; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_3 = 4'h3 == io_ar_addr ? btb_3_true_branch_state : _GEN_2; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_4 = 4'h4 == io_ar_addr ? btb_4_true_branch_state : _GEN_3; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_5 = 4'h5 == io_ar_addr ? btb_5_true_branch_state : _GEN_4; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_6 = 4'h6 == io_ar_addr ? btb_6_true_branch_state : _GEN_5; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_7 = 4'h7 == io_ar_addr ? btb_7_true_branch_state : _GEN_6; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_8 = 4'h8 == io_ar_addr ? btb_8_true_branch_state : _GEN_7; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_9 = 4'h9 == io_ar_addr ? btb_9_true_branch_state : _GEN_8; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_10 = 4'ha == io_ar_addr ? btb_10_true_branch_state : _GEN_9; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_11 = 4'hb == io_ar_addr ? btb_11_true_branch_state : _GEN_10; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_12 = 4'hc == io_ar_addr ? btb_12_true_branch_state : _GEN_11; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_13 = 4'hd == io_ar_addr ? btb_13_true_branch_state : _GEN_12; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_14 = 4'he == io_ar_addr ? btb_14_true_branch_state : _GEN_13; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_17 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_jr : btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_18 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_jr : _GEN_17; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_19 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_jr : _GEN_18; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_20 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_jr : _GEN_19; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_21 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_jr : _GEN_20; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_22 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_jr : _GEN_21; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_23 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_jr : _GEN_22; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_24 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_jr : _GEN_23; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_25 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_jr : _GEN_24; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_26 = 4'ha == io_ar_addr ? btb_10_pre_decoder_jr : _GEN_25; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_27 = 4'hb == io_ar_addr ? btb_11_pre_decoder_jr : _GEN_26; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_28 = 4'hc == io_ar_addr ? btb_12_pre_decoder_jr : _GEN_27; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_29 = 4'hd == io_ar_addr ? btb_13_pre_decoder_jr : _GEN_28; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_30 = 4'he == io_ar_addr ? btb_14_pre_decoder_jr : _GEN_29; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_33 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_branchdata : btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_34 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_branchdata : _GEN_33; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_35 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_branchdata : _GEN_34; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_36 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_branchdata : _GEN_35; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_37 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_branchdata : _GEN_36; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_38 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_branchdata : _GEN_37; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_39 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_branchdata : _GEN_38; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_40 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_branchdata : _GEN_39; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_41 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_branchdata : _GEN_40; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_42 = 4'ha == io_ar_addr ? btb_10_pre_decoder_branchdata : _GEN_41; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_43 = 4'hb == io_ar_addr ? btb_11_pre_decoder_branchdata : _GEN_42; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_44 = 4'hc == io_ar_addr ? btb_12_pre_decoder_branchdata : _GEN_43; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_45 = 4'hd == io_ar_addr ? btb_13_pre_decoder_branchdata : _GEN_44; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_46 = 4'he == io_ar_addr ? btb_14_pre_decoder_branchdata : _GEN_45; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_49 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_jump : btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_50 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_jump : _GEN_49; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_51 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_jump : _GEN_50; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_52 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_jump : _GEN_51; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_53 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_jump : _GEN_52; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_54 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_jump : _GEN_53; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_55 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_jump : _GEN_54; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_56 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_jump : _GEN_55; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_57 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_jump : _GEN_56; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_58 = 4'ha == io_ar_addr ? btb_10_pre_decoder_jump : _GEN_57; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_59 = 4'hb == io_ar_addr ? btb_11_pre_decoder_jump : _GEN_58; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_60 = 4'hc == io_ar_addr ? btb_12_pre_decoder_jump : _GEN_59; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_61 = 4'hd == io_ar_addr ? btb_13_pre_decoder_jump : _GEN_60; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_62 = 4'he == io_ar_addr ? btb_14_pre_decoder_jump : _GEN_61; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_65 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_branchD_flag : btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_66 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_branchD_flag : _GEN_65; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_67 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_branchD_flag : _GEN_66; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_68 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_branchD_flag : _GEN_67; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_69 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_branchD_flag : _GEN_68; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_70 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_branchD_flag : _GEN_69; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_71 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_branchD_flag : _GEN_70; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_72 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_branchD_flag : _GEN_71; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_73 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_branchD_flag : _GEN_72; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_74 = 4'ha == io_ar_addr ? btb_10_pre_decoder_branchD_flag : _GEN_73; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_75 = 4'hb == io_ar_addr ? btb_11_pre_decoder_branchD_flag : _GEN_74; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_76 = 4'hc == io_ar_addr ? btb_12_pre_decoder_branchD_flag : _GEN_75; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_77 = 4'hd == io_ar_addr ? btb_13_pre_decoder_branchD_flag : _GEN_76; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_78 = 4'he == io_ar_addr ? btb_14_pre_decoder_branchD_flag : _GEN_77; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_81 = 4'h1 == io_ar_addr ? btb_1_pre_bht : btb_0_pre_bht; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_82 = 4'h2 == io_ar_addr ? btb_2_pre_bht : _GEN_81; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_83 = 4'h3 == io_ar_addr ? btb_3_pre_bht : _GEN_82; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_84 = 4'h4 == io_ar_addr ? btb_4_pre_bht : _GEN_83; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_85 = 4'h5 == io_ar_addr ? btb_5_pre_bht : _GEN_84; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_86 = 4'h6 == io_ar_addr ? btb_6_pre_bht : _GEN_85; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_87 = 4'h7 == io_ar_addr ? btb_7_pre_bht : _GEN_86; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_88 = 4'h8 == io_ar_addr ? btb_8_pre_bht : _GEN_87; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_89 = 4'h9 == io_ar_addr ? btb_9_pre_bht : _GEN_88; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_90 = 4'ha == io_ar_addr ? btb_10_pre_bht : _GEN_89; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_91 = 4'hb == io_ar_addr ? btb_11_pre_bht : _GEN_90; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_92 = 4'hc == io_ar_addr ? btb_12_pre_bht : _GEN_91; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_93 = 4'hd == io_ar_addr ? btb_13_pre_bht : _GEN_92; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_94 = 4'he == io_ar_addr ? btb_14_pre_bht : _GEN_93; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_97 = 4'h1 == io_ar_addr ? btb_1_pre_pht : btb_0_pre_pht; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_98 = 4'h2 == io_ar_addr ? btb_2_pre_pht : _GEN_97; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_99 = 4'h3 == io_ar_addr ? btb_3_pre_pht : _GEN_98; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_100 = 4'h4 == io_ar_addr ? btb_4_pre_pht : _GEN_99; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_101 = 4'h5 == io_ar_addr ? btb_5_pre_pht : _GEN_100; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_102 = 4'h6 == io_ar_addr ? btb_6_pre_pht : _GEN_101; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_103 = 4'h7 == io_ar_addr ? btb_7_pre_pht : _GEN_102; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_104 = 4'h8 == io_ar_addr ? btb_8_pre_pht : _GEN_103; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_105 = 4'h9 == io_ar_addr ? btb_9_pre_pht : _GEN_104; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_106 = 4'ha == io_ar_addr ? btb_10_pre_pht : _GEN_105; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_107 = 4'hb == io_ar_addr ? btb_11_pre_pht : _GEN_106; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_108 = 4'hc == io_ar_addr ? btb_12_pre_pht : _GEN_107; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_109 = 4'hd == io_ar_addr ? btb_13_pre_pht : _GEN_108; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_110 = 4'he == io_ar_addr ? btb_14_pre_pht : _GEN_109; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_113 = 4'h1 == io_ar_addr ? btb_1_pre_hashcode : btb_0_pre_hashcode; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_114 = 4'h2 == io_ar_addr ? btb_2_pre_hashcode : _GEN_113; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_115 = 4'h3 == io_ar_addr ? btb_3_pre_hashcode : _GEN_114; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_116 = 4'h4 == io_ar_addr ? btb_4_pre_hashcode : _GEN_115; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_117 = 4'h5 == io_ar_addr ? btb_5_pre_hashcode : _GEN_116; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_118 = 4'h6 == io_ar_addr ? btb_6_pre_hashcode : _GEN_117; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_119 = 4'h7 == io_ar_addr ? btb_7_pre_hashcode : _GEN_118; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_120 = 4'h8 == io_ar_addr ? btb_8_pre_hashcode : _GEN_119; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_121 = 4'h9 == io_ar_addr ? btb_9_pre_hashcode : _GEN_120; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_122 = 4'ha == io_ar_addr ? btb_10_pre_hashcode : _GEN_121; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_123 = 4'hb == io_ar_addr ? btb_11_pre_hashcode : _GEN_122; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_124 = 4'hc == io_ar_addr ? btb_12_pre_hashcode : _GEN_123; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_125 = 4'hd == io_ar_addr ? btb_13_pre_hashcode : _GEN_124; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_126 = 4'he == io_ar_addr ? btb_14_pre_hashcode : _GEN_125; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_129 = 4'h1 == io_ar_addr ? btb_1_pre_lookup_data : btb_0_pre_lookup_data; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_130 = 4'h2 == io_ar_addr ? btb_2_pre_lookup_data : _GEN_129; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_131 = 4'h3 == io_ar_addr ? btb_3_pre_lookup_data : _GEN_130; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_132 = 4'h4 == io_ar_addr ? btb_4_pre_lookup_data : _GEN_131; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_133 = 4'h5 == io_ar_addr ? btb_5_pre_lookup_data : _GEN_132; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_134 = 4'h6 == io_ar_addr ? btb_6_pre_lookup_data : _GEN_133; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_135 = 4'h7 == io_ar_addr ? btb_7_pre_lookup_data : _GEN_134; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_136 = 4'h8 == io_ar_addr ? btb_8_pre_lookup_data : _GEN_135; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_137 = 4'h9 == io_ar_addr ? btb_9_pre_lookup_data : _GEN_136; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_138 = 4'ha == io_ar_addr ? btb_10_pre_lookup_data : _GEN_137; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_139 = 4'hb == io_ar_addr ? btb_11_pre_lookup_data : _GEN_138; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_140 = 4'hc == io_ar_addr ? btb_12_pre_lookup_data : _GEN_139; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_141 = 4'hd == io_ar_addr ? btb_13_pre_lookup_data : _GEN_140; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_142 = 4'he == io_ar_addr ? btb_14_pre_lookup_data : _GEN_141; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_145 = 4'h1 == io_ar_addr ? btb_1_pre_pc_target : btb_0_pre_pc_target; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_146 = 4'h2 == io_ar_addr ? btb_2_pre_pc_target : _GEN_145; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_147 = 4'h3 == io_ar_addr ? btb_3_pre_pc_target : _GEN_146; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_148 = 4'h4 == io_ar_addr ? btb_4_pre_pc_target : _GEN_147; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_149 = 4'h5 == io_ar_addr ? btb_5_pre_pc_target : _GEN_148; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_150 = 4'h6 == io_ar_addr ? btb_6_pre_pc_target : _GEN_149; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_151 = 4'h7 == io_ar_addr ? btb_7_pre_pc_target : _GEN_150; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_152 = 4'h8 == io_ar_addr ? btb_8_pre_pc_target : _GEN_151; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_153 = 4'h9 == io_ar_addr ? btb_9_pre_pc_target : _GEN_152; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_154 = 4'ha == io_ar_addr ? btb_10_pre_pc_target : _GEN_153; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_155 = 4'hb == io_ar_addr ? btb_11_pre_pc_target : _GEN_154; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_156 = 4'hc == io_ar_addr ? btb_12_pre_pc_target : _GEN_155; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_157 = 4'hd == io_ar_addr ? btb_13_pre_pc_target : _GEN_156; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_158 = 4'he == io_ar_addr ? btb_14_pre_pc_target : _GEN_157; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_161 = 4'h1 == io_ar_addr ? btb_1_exception_type : btb_0_exception_type; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_162 = 4'h2 == io_ar_addr ? btb_2_exception_type : _GEN_161; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_163 = 4'h3 == io_ar_addr ? btb_3_exception_type : _GEN_162; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_164 = 4'h4 == io_ar_addr ? btb_4_exception_type : _GEN_163; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_165 = 4'h5 == io_ar_addr ? btb_5_exception_type : _GEN_164; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_166 = 4'h6 == io_ar_addr ? btb_6_exception_type : _GEN_165; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_167 = 4'h7 == io_ar_addr ? btb_7_exception_type : _GEN_166; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_168 = 4'h8 == io_ar_addr ? btb_8_exception_type : _GEN_167; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_169 = 4'h9 == io_ar_addr ? btb_9_exception_type : _GEN_168; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_170 = 4'ha == io_ar_addr ? btb_10_exception_type : _GEN_169; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_171 = 4'hb == io_ar_addr ? btb_11_exception_type : _GEN_170; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_172 = 4'hc == io_ar_addr ? btb_12_exception_type : _GEN_171; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_173 = 4'hd == io_ar_addr ? btb_13_exception_type : _GEN_172; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_174 = 4'he == io_ar_addr ? btb_14_exception_type : _GEN_173; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_177 = 4'h1 == io_ar_addr ? btb_1_inst : btb_0_inst; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_178 = 4'h2 == io_ar_addr ? btb_2_inst : _GEN_177; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_179 = 4'h3 == io_ar_addr ? btb_3_inst : _GEN_178; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_180 = 4'h4 == io_ar_addr ? btb_4_inst : _GEN_179; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_181 = 4'h5 == io_ar_addr ? btb_5_inst : _GEN_180; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_182 = 4'h6 == io_ar_addr ? btb_6_inst : _GEN_181; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_183 = 4'h7 == io_ar_addr ? btb_7_inst : _GEN_182; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_184 = 4'h8 == io_ar_addr ? btb_8_inst : _GEN_183; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_185 = 4'h9 == io_ar_addr ? btb_9_inst : _GEN_184; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_186 = 4'ha == io_ar_addr ? btb_10_inst : _GEN_185; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_187 = 4'hb == io_ar_addr ? btb_11_inst : _GEN_186; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_188 = 4'hc == io_ar_addr ? btb_12_inst : _GEN_187; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_189 = 4'hd == io_ar_addr ? btb_13_inst : _GEN_188; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_190 = 4'he == io_ar_addr ? btb_14_inst : _GEN_189; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_193 = 4'h1 == io_ar_addr ? btb_1_pc : btb_0_pc; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_194 = 4'h2 == io_ar_addr ? btb_2_pc : _GEN_193; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_195 = 4'h3 == io_ar_addr ? btb_3_pc : _GEN_194; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_196 = 4'h4 == io_ar_addr ? btb_4_pc : _GEN_195; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_197 = 4'h5 == io_ar_addr ? btb_5_pc : _GEN_196; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_198 = 4'h6 == io_ar_addr ? btb_6_pc : _GEN_197; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_199 = 4'h7 == io_ar_addr ? btb_7_pc : _GEN_198; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_200 = 4'h8 == io_ar_addr ? btb_8_pc : _GEN_199; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_201 = 4'h9 == io_ar_addr ? btb_9_pc : _GEN_200; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_202 = 4'ha == io_ar_addr ? btb_10_pc : _GEN_201; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_203 = 4'hb == io_ar_addr ? btb_11_pc : _GEN_202; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_204 = 4'hc == io_ar_addr ? btb_12_pc : _GEN_203; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_205 = 4'hd == io_ar_addr ? btb_13_pc : _GEN_204; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_206 = 4'he == io_ar_addr ? btb_14_pc : _GEN_205; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_221 = 4'h1 == io_aw_addr ? btb_1_pc : btb_0_pc; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_222 = 4'h1 == io_aw_addr ? btb_1_inst : btb_0_inst; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_223 = 4'h1 == io_aw_addr ? btb_1_exception_type : btb_0_exception_type; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_224 = 4'h1 == io_aw_addr ? btb_1_pre_pc_target : btb_0_pre_pc_target; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_225 = 4'h1 == io_aw_addr ? btb_1_pre_lookup_data : btb_0_pre_lookup_data; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_226 = 4'h1 == io_aw_addr ? btb_1_pre_hashcode : btb_0_pre_hashcode; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_227 = 4'h1 == io_aw_addr ? btb_1_pre_pht : btb_0_pre_pht; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_228 = 4'h1 == io_aw_addr ? btb_1_pre_bht : btb_0_pre_bht; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_229 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_branchD_flag : btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_230 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_jump : btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_231 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_branchdata : btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_232 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_jr : btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_233 = 4'h1 == io_aw_addr ? btb_1_true_branch_state : btb_0_true_branch_state; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_234 = 4'h2 == io_aw_addr ? btb_2_pc : _GEN_221; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_235 = 4'h2 == io_aw_addr ? btb_2_inst : _GEN_222; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_236 = 4'h2 == io_aw_addr ? btb_2_exception_type : _GEN_223; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_237 = 4'h2 == io_aw_addr ? btb_2_pre_pc_target : _GEN_224; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_238 = 4'h2 == io_aw_addr ? btb_2_pre_lookup_data : _GEN_225; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_239 = 4'h2 == io_aw_addr ? btb_2_pre_hashcode : _GEN_226; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_240 = 4'h2 == io_aw_addr ? btb_2_pre_pht : _GEN_227; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_241 = 4'h2 == io_aw_addr ? btb_2_pre_bht : _GEN_228; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_242 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_branchD_flag : _GEN_229; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_243 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_jump : _GEN_230; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_244 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_branchdata : _GEN_231; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_245 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_jr : _GEN_232; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_246 = 4'h2 == io_aw_addr ? btb_2_true_branch_state : _GEN_233; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_247 = 4'h3 == io_aw_addr ? btb_3_pc : _GEN_234; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_248 = 4'h3 == io_aw_addr ? btb_3_inst : _GEN_235; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_249 = 4'h3 == io_aw_addr ? btb_3_exception_type : _GEN_236; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_250 = 4'h3 == io_aw_addr ? btb_3_pre_pc_target : _GEN_237; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_251 = 4'h3 == io_aw_addr ? btb_3_pre_lookup_data : _GEN_238; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_252 = 4'h3 == io_aw_addr ? btb_3_pre_hashcode : _GEN_239; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_253 = 4'h3 == io_aw_addr ? btb_3_pre_pht : _GEN_240; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_254 = 4'h3 == io_aw_addr ? btb_3_pre_bht : _GEN_241; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_255 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_branchD_flag : _GEN_242; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_256 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_jump : _GEN_243; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_257 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_branchdata : _GEN_244; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_258 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_jr : _GEN_245; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_259 = 4'h3 == io_aw_addr ? btb_3_true_branch_state : _GEN_246; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_260 = 4'h4 == io_aw_addr ? btb_4_pc : _GEN_247; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_261 = 4'h4 == io_aw_addr ? btb_4_inst : _GEN_248; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_262 = 4'h4 == io_aw_addr ? btb_4_exception_type : _GEN_249; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_263 = 4'h4 == io_aw_addr ? btb_4_pre_pc_target : _GEN_250; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_264 = 4'h4 == io_aw_addr ? btb_4_pre_lookup_data : _GEN_251; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_265 = 4'h4 == io_aw_addr ? btb_4_pre_hashcode : _GEN_252; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_266 = 4'h4 == io_aw_addr ? btb_4_pre_pht : _GEN_253; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_267 = 4'h4 == io_aw_addr ? btb_4_pre_bht : _GEN_254; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_268 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_branchD_flag : _GEN_255; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_269 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_jump : _GEN_256; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_270 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_branchdata : _GEN_257; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_271 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_jr : _GEN_258; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_272 = 4'h4 == io_aw_addr ? btb_4_true_branch_state : _GEN_259; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_273 = 4'h5 == io_aw_addr ? btb_5_pc : _GEN_260; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_274 = 4'h5 == io_aw_addr ? btb_5_inst : _GEN_261; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_275 = 4'h5 == io_aw_addr ? btb_5_exception_type : _GEN_262; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_276 = 4'h5 == io_aw_addr ? btb_5_pre_pc_target : _GEN_263; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_277 = 4'h5 == io_aw_addr ? btb_5_pre_lookup_data : _GEN_264; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_278 = 4'h5 == io_aw_addr ? btb_5_pre_hashcode : _GEN_265; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_279 = 4'h5 == io_aw_addr ? btb_5_pre_pht : _GEN_266; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_280 = 4'h5 == io_aw_addr ? btb_5_pre_bht : _GEN_267; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_281 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_branchD_flag : _GEN_268; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_282 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_jump : _GEN_269; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_283 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_branchdata : _GEN_270; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_284 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_jr : _GEN_271; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_285 = 4'h5 == io_aw_addr ? btb_5_true_branch_state : _GEN_272; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_286 = 4'h6 == io_aw_addr ? btb_6_pc : _GEN_273; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_287 = 4'h6 == io_aw_addr ? btb_6_inst : _GEN_274; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_288 = 4'h6 == io_aw_addr ? btb_6_exception_type : _GEN_275; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_289 = 4'h6 == io_aw_addr ? btb_6_pre_pc_target : _GEN_276; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_290 = 4'h6 == io_aw_addr ? btb_6_pre_lookup_data : _GEN_277; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_291 = 4'h6 == io_aw_addr ? btb_6_pre_hashcode : _GEN_278; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_292 = 4'h6 == io_aw_addr ? btb_6_pre_pht : _GEN_279; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_293 = 4'h6 == io_aw_addr ? btb_6_pre_bht : _GEN_280; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_294 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_branchD_flag : _GEN_281; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_295 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_jump : _GEN_282; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_296 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_branchdata : _GEN_283; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_297 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_jr : _GEN_284; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_298 = 4'h6 == io_aw_addr ? btb_6_true_branch_state : _GEN_285; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_299 = 4'h7 == io_aw_addr ? btb_7_pc : _GEN_286; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_300 = 4'h7 == io_aw_addr ? btb_7_inst : _GEN_287; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_301 = 4'h7 == io_aw_addr ? btb_7_exception_type : _GEN_288; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_302 = 4'h7 == io_aw_addr ? btb_7_pre_pc_target : _GEN_289; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_303 = 4'h7 == io_aw_addr ? btb_7_pre_lookup_data : _GEN_290; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_304 = 4'h7 == io_aw_addr ? btb_7_pre_hashcode : _GEN_291; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_305 = 4'h7 == io_aw_addr ? btb_7_pre_pht : _GEN_292; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_306 = 4'h7 == io_aw_addr ? btb_7_pre_bht : _GEN_293; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_307 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_branchD_flag : _GEN_294; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_308 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_jump : _GEN_295; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_309 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_branchdata : _GEN_296; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_310 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_jr : _GEN_297; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_311 = 4'h7 == io_aw_addr ? btb_7_true_branch_state : _GEN_298; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_312 = 4'h8 == io_aw_addr ? btb_8_pc : _GEN_299; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_313 = 4'h8 == io_aw_addr ? btb_8_inst : _GEN_300; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_314 = 4'h8 == io_aw_addr ? btb_8_exception_type : _GEN_301; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_315 = 4'h8 == io_aw_addr ? btb_8_pre_pc_target : _GEN_302; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_316 = 4'h8 == io_aw_addr ? btb_8_pre_lookup_data : _GEN_303; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_317 = 4'h8 == io_aw_addr ? btb_8_pre_hashcode : _GEN_304; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_318 = 4'h8 == io_aw_addr ? btb_8_pre_pht : _GEN_305; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_319 = 4'h8 == io_aw_addr ? btb_8_pre_bht : _GEN_306; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_320 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_branchD_flag : _GEN_307; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_321 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_jump : _GEN_308; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_322 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_branchdata : _GEN_309; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_323 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_jr : _GEN_310; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_324 = 4'h8 == io_aw_addr ? btb_8_true_branch_state : _GEN_311; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_325 = 4'h9 == io_aw_addr ? btb_9_pc : _GEN_312; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_326 = 4'h9 == io_aw_addr ? btb_9_inst : _GEN_313; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_327 = 4'h9 == io_aw_addr ? btb_9_exception_type : _GEN_314; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_328 = 4'h9 == io_aw_addr ? btb_9_pre_pc_target : _GEN_315; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_329 = 4'h9 == io_aw_addr ? btb_9_pre_lookup_data : _GEN_316; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_330 = 4'h9 == io_aw_addr ? btb_9_pre_hashcode : _GEN_317; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_331 = 4'h9 == io_aw_addr ? btb_9_pre_pht : _GEN_318; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_332 = 4'h9 == io_aw_addr ? btb_9_pre_bht : _GEN_319; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_333 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_branchD_flag : _GEN_320; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_334 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_jump : _GEN_321; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_335 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_branchdata : _GEN_322; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_336 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_jr : _GEN_323; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_337 = 4'h9 == io_aw_addr ? btb_9_true_branch_state : _GEN_324; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_338 = 4'ha == io_aw_addr ? btb_10_pc : _GEN_325; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_339 = 4'ha == io_aw_addr ? btb_10_inst : _GEN_326; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_340 = 4'ha == io_aw_addr ? btb_10_exception_type : _GEN_327; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_341 = 4'ha == io_aw_addr ? btb_10_pre_pc_target : _GEN_328; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_342 = 4'ha == io_aw_addr ? btb_10_pre_lookup_data : _GEN_329; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_343 = 4'ha == io_aw_addr ? btb_10_pre_hashcode : _GEN_330; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_344 = 4'ha == io_aw_addr ? btb_10_pre_pht : _GEN_331; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_345 = 4'ha == io_aw_addr ? btb_10_pre_bht : _GEN_332; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_346 = 4'ha == io_aw_addr ? btb_10_pre_decoder_branchD_flag : _GEN_333; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_347 = 4'ha == io_aw_addr ? btb_10_pre_decoder_jump : _GEN_334; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_348 = 4'ha == io_aw_addr ? btb_10_pre_decoder_branchdata : _GEN_335; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_349 = 4'ha == io_aw_addr ? btb_10_pre_decoder_jr : _GEN_336; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_350 = 4'ha == io_aw_addr ? btb_10_true_branch_state : _GEN_337; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_351 = 4'hb == io_aw_addr ? btb_11_pc : _GEN_338; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_352 = 4'hb == io_aw_addr ? btb_11_inst : _GEN_339; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_353 = 4'hb == io_aw_addr ? btb_11_exception_type : _GEN_340; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_354 = 4'hb == io_aw_addr ? btb_11_pre_pc_target : _GEN_341; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_355 = 4'hb == io_aw_addr ? btb_11_pre_lookup_data : _GEN_342; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_356 = 4'hb == io_aw_addr ? btb_11_pre_hashcode : _GEN_343; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_357 = 4'hb == io_aw_addr ? btb_11_pre_pht : _GEN_344; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_358 = 4'hb == io_aw_addr ? btb_11_pre_bht : _GEN_345; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_359 = 4'hb == io_aw_addr ? btb_11_pre_decoder_branchD_flag : _GEN_346; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_360 = 4'hb == io_aw_addr ? btb_11_pre_decoder_jump : _GEN_347; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_361 = 4'hb == io_aw_addr ? btb_11_pre_decoder_branchdata : _GEN_348; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_362 = 4'hb == io_aw_addr ? btb_11_pre_decoder_jr : _GEN_349; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_363 = 4'hb == io_aw_addr ? btb_11_true_branch_state : _GEN_350; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_364 = 4'hc == io_aw_addr ? btb_12_pc : _GEN_351; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_365 = 4'hc == io_aw_addr ? btb_12_inst : _GEN_352; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_366 = 4'hc == io_aw_addr ? btb_12_exception_type : _GEN_353; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_367 = 4'hc == io_aw_addr ? btb_12_pre_pc_target : _GEN_354; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_368 = 4'hc == io_aw_addr ? btb_12_pre_lookup_data : _GEN_355; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_369 = 4'hc == io_aw_addr ? btb_12_pre_hashcode : _GEN_356; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_370 = 4'hc == io_aw_addr ? btb_12_pre_pht : _GEN_357; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_371 = 4'hc == io_aw_addr ? btb_12_pre_bht : _GEN_358; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_372 = 4'hc == io_aw_addr ? btb_12_pre_decoder_branchD_flag : _GEN_359; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_373 = 4'hc == io_aw_addr ? btb_12_pre_decoder_jump : _GEN_360; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_374 = 4'hc == io_aw_addr ? btb_12_pre_decoder_branchdata : _GEN_361; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_375 = 4'hc == io_aw_addr ? btb_12_pre_decoder_jr : _GEN_362; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_376 = 4'hc == io_aw_addr ? btb_12_true_branch_state : _GEN_363; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_377 = 4'hd == io_aw_addr ? btb_13_pc : _GEN_364; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_378 = 4'hd == io_aw_addr ? btb_13_inst : _GEN_365; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_379 = 4'hd == io_aw_addr ? btb_13_exception_type : _GEN_366; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_380 = 4'hd == io_aw_addr ? btb_13_pre_pc_target : _GEN_367; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_381 = 4'hd == io_aw_addr ? btb_13_pre_lookup_data : _GEN_368; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_382 = 4'hd == io_aw_addr ? btb_13_pre_hashcode : _GEN_369; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_383 = 4'hd == io_aw_addr ? btb_13_pre_pht : _GEN_370; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_384 = 4'hd == io_aw_addr ? btb_13_pre_bht : _GEN_371; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_385 = 4'hd == io_aw_addr ? btb_13_pre_decoder_branchD_flag : _GEN_372; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_386 = 4'hd == io_aw_addr ? btb_13_pre_decoder_jump : _GEN_373; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_387 = 4'hd == io_aw_addr ? btb_13_pre_decoder_branchdata : _GEN_374; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_388 = 4'hd == io_aw_addr ? btb_13_pre_decoder_jr : _GEN_375; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_389 = 4'hd == io_aw_addr ? btb_13_true_branch_state : _GEN_376; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_390 = 4'he == io_aw_addr ? btb_14_pc : _GEN_377; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_391 = 4'he == io_aw_addr ? btb_14_inst : _GEN_378; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_392 = 4'he == io_aw_addr ? btb_14_exception_type : _GEN_379; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_393 = 4'he == io_aw_addr ? btb_14_pre_pc_target : _GEN_380; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_394 = 4'he == io_aw_addr ? btb_14_pre_lookup_data : _GEN_381; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_395 = 4'he == io_aw_addr ? btb_14_pre_hashcode : _GEN_382; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_396 = 4'he == io_aw_addr ? btb_14_pre_pht : _GEN_383; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_397 = 4'he == io_aw_addr ? btb_14_pre_bht : _GEN_384; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_398 = 4'he == io_aw_addr ? btb_14_pre_decoder_branchD_flag : _GEN_385; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_399 = 4'he == io_aw_addr ? btb_14_pre_decoder_jump : _GEN_386; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_400 = 4'he == io_aw_addr ? btb_14_pre_decoder_branchdata : _GEN_387; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_401 = 4'he == io_aw_addr ? btb_14_pre_decoder_jr : _GEN_388; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_402 = 4'he == io_aw_addr ? btb_14_true_branch_state : _GEN_389; // @[ports_lookup_table.scala 107:{27,27}]
  assign io_out_pc = 4'hf == io_ar_addr ? btb_15_pc : _GEN_206; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_inst = 4'hf == io_ar_addr ? btb_15_inst : _GEN_190; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_exception_type = 4'hf == io_ar_addr ? btb_15_exception_type : _GEN_174; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_pc_target = 4'hf == io_ar_addr ? btb_15_pre_pc_target : _GEN_158; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_lookup_data = 4'hf == io_ar_addr ? btb_15_pre_lookup_data : _GEN_142; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_hashcode = 4'hf == io_ar_addr ? btb_15_pre_hashcode : _GEN_126; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_pht = 4'hf == io_ar_addr ? btb_15_pre_pht : _GEN_110; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_bht = 4'hf == io_ar_addr ? btb_15_pre_bht : _GEN_94; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_branchD_flag = 4'hf == io_ar_addr ? btb_15_pre_decoder_branchD_flag : _GEN_78; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_jump = 4'hf == io_ar_addr ? btb_15_pre_decoder_jump : _GEN_62; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_branchdata = 4'hf == io_ar_addr ? btb_15_pre_decoder_branchdata : _GEN_46; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_jr = 4'hf == io_ar_addr ? btb_15_pre_decoder_jr : _GEN_30; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_true_branch_state = 4'hf == io_ar_addr ? btb_15_true_branch_state : _GEN_14; // @[ports_lookup_table.scala 106:{12,12}]
  always @(posedge clock) begin
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_0_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_0_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_0_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_0_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_1_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_1_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_1_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_1_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_2_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_2_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_2_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_2_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_3_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_3_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_3_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_3_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_4_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_4_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_4_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_4_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_5_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_5_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_5_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_5_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_6_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_6_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_6_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_6_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_7_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_7_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_7_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_7_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_8_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_8_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_8_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_8_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_9_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_9_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_9_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_9_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_10_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_10_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_10_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_10_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_11_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_11_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_11_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_11_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_12_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_12_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_12_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_12_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_13_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_13_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_13_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_13_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pc <= btb_15_pc; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_inst <= btb_15_inst; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_exception_type <= btb_15_exception_type; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_pc_target <= btb_15_pre_pc_target; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_lookup_data <= btb_15_pre_lookup_data; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_hashcode <= btb_15_pre_hashcode; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_pht <= btb_15_pre_pht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_bht <= btb_15_pre_bht; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_jump <= btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_pre_decoder_jr <= btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_14_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_14_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:27]
        btb_14_true_branch_state <= btb_15_true_branch_state; // @[ports_lookup_table.scala 107:27]
      end else begin
        btb_14_true_branch_state <= _GEN_402;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pc <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pc <= io_in_pc;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pc <= _GEN_390;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_inst <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_inst <= io_in_inst;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_inst <= _GEN_391;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_exception_type <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_exception_type <= 2'h0;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_exception_type <= _GEN_392;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_pc_target <= 32'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_pc_target <= io_in_pre_pc_target;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_pc_target <= _GEN_393;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_lookup_data <= _GEN_394;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_hashcode <= io_in_pre_hashcode;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_hashcode <= _GEN_395;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_pht <= 2'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_pht <= io_in_pre_pht;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_pht <= _GEN_396;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_bht <= 7'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_bht <= io_in_pre_bht;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_bht <= _GEN_397;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_branchD_flag <= _GEN_398;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_jump <= _GEN_399;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_branchdata <= _GEN_400;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_pre_decoder_jr <= _GEN_401;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 105:22]
      btb_15_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 105:22]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 107:21]
      if (io_write) begin // @[ports_lookup_table.scala 107:27]
        btb_15_true_branch_state <= io_in_true_branch_state;
      end else if (!(4'hf == io_aw_addr)) begin // @[ports_lookup_table.scala 107:27]
        btb_15_true_branch_state <= _GEN_402;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  btb_0_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  btb_0_exception_type = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  btb_0_pre_pc_target = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  btb_0_pre_lookup_data = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  btb_0_pre_hashcode = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  btb_0_pre_pht = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  btb_0_pre_bht = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  btb_0_pre_decoder_branchD_flag = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btb_0_pre_decoder_jump = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btb_0_pre_decoder_branchdata = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  btb_0_pre_decoder_jr = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  btb_0_true_branch_state = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btb_1_pc = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  btb_1_inst = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  btb_1_exception_type = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  btb_1_pre_pc_target = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  btb_1_pre_lookup_data = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  btb_1_pre_hashcode = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  btb_1_pre_pht = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  btb_1_pre_bht = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  btb_1_pre_decoder_branchD_flag = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  btb_1_pre_decoder_jump = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  btb_1_pre_decoder_branchdata = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  btb_1_pre_decoder_jr = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  btb_1_true_branch_state = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  btb_2_pc = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  btb_2_inst = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  btb_2_exception_type = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  btb_2_pre_pc_target = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  btb_2_pre_lookup_data = _RAND_30[6:0];
  _RAND_31 = {1{`RANDOM}};
  btb_2_pre_hashcode = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  btb_2_pre_pht = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  btb_2_pre_bht = _RAND_33[6:0];
  _RAND_34 = {1{`RANDOM}};
  btb_2_pre_decoder_branchD_flag = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  btb_2_pre_decoder_jump = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  btb_2_pre_decoder_branchdata = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  btb_2_pre_decoder_jr = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  btb_2_true_branch_state = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  btb_3_pc = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  btb_3_inst = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  btb_3_exception_type = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  btb_3_pre_pc_target = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  btb_3_pre_lookup_data = _RAND_43[6:0];
  _RAND_44 = {1{`RANDOM}};
  btb_3_pre_hashcode = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  btb_3_pre_pht = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  btb_3_pre_bht = _RAND_46[6:0];
  _RAND_47 = {1{`RANDOM}};
  btb_3_pre_decoder_branchD_flag = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  btb_3_pre_decoder_jump = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  btb_3_pre_decoder_branchdata = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  btb_3_pre_decoder_jr = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  btb_3_true_branch_state = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  btb_4_pc = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  btb_4_inst = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  btb_4_exception_type = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  btb_4_pre_pc_target = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  btb_4_pre_lookup_data = _RAND_56[6:0];
  _RAND_57 = {1{`RANDOM}};
  btb_4_pre_hashcode = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  btb_4_pre_pht = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  btb_4_pre_bht = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  btb_4_pre_decoder_branchD_flag = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  btb_4_pre_decoder_jump = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  btb_4_pre_decoder_branchdata = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  btb_4_pre_decoder_jr = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  btb_4_true_branch_state = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  btb_5_pc = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  btb_5_inst = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  btb_5_exception_type = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  btb_5_pre_pc_target = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  btb_5_pre_lookup_data = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  btb_5_pre_hashcode = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  btb_5_pre_pht = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  btb_5_pre_bht = _RAND_72[6:0];
  _RAND_73 = {1{`RANDOM}};
  btb_5_pre_decoder_branchD_flag = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  btb_5_pre_decoder_jump = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  btb_5_pre_decoder_branchdata = _RAND_75[5:0];
  _RAND_76 = {1{`RANDOM}};
  btb_5_pre_decoder_jr = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  btb_5_true_branch_state = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  btb_6_pc = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  btb_6_inst = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  btb_6_exception_type = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  btb_6_pre_pc_target = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  btb_6_pre_lookup_data = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  btb_6_pre_hashcode = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  btb_6_pre_pht = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  btb_6_pre_bht = _RAND_85[6:0];
  _RAND_86 = {1{`RANDOM}};
  btb_6_pre_decoder_branchD_flag = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  btb_6_pre_decoder_jump = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  btb_6_pre_decoder_branchdata = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  btb_6_pre_decoder_jr = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  btb_6_true_branch_state = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  btb_7_pc = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  btb_7_inst = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  btb_7_exception_type = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  btb_7_pre_pc_target = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  btb_7_pre_lookup_data = _RAND_95[6:0];
  _RAND_96 = {1{`RANDOM}};
  btb_7_pre_hashcode = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  btb_7_pre_pht = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  btb_7_pre_bht = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  btb_7_pre_decoder_branchD_flag = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  btb_7_pre_decoder_jump = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  btb_7_pre_decoder_branchdata = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  btb_7_pre_decoder_jr = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  btb_7_true_branch_state = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  btb_8_pc = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  btb_8_inst = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  btb_8_exception_type = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  btb_8_pre_pc_target = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  btb_8_pre_lookup_data = _RAND_108[6:0];
  _RAND_109 = {1{`RANDOM}};
  btb_8_pre_hashcode = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  btb_8_pre_pht = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  btb_8_pre_bht = _RAND_111[6:0];
  _RAND_112 = {1{`RANDOM}};
  btb_8_pre_decoder_branchD_flag = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  btb_8_pre_decoder_jump = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  btb_8_pre_decoder_branchdata = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  btb_8_pre_decoder_jr = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  btb_8_true_branch_state = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  btb_9_pc = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  btb_9_inst = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  btb_9_exception_type = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  btb_9_pre_pc_target = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  btb_9_pre_lookup_data = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  btb_9_pre_hashcode = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  btb_9_pre_pht = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  btb_9_pre_bht = _RAND_124[6:0];
  _RAND_125 = {1{`RANDOM}};
  btb_9_pre_decoder_branchD_flag = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  btb_9_pre_decoder_jump = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  btb_9_pre_decoder_branchdata = _RAND_127[5:0];
  _RAND_128 = {1{`RANDOM}};
  btb_9_pre_decoder_jr = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  btb_9_true_branch_state = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  btb_10_pc = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  btb_10_inst = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  btb_10_exception_type = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  btb_10_pre_pc_target = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  btb_10_pre_lookup_data = _RAND_134[6:0];
  _RAND_135 = {1{`RANDOM}};
  btb_10_pre_hashcode = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  btb_10_pre_pht = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  btb_10_pre_bht = _RAND_137[6:0];
  _RAND_138 = {1{`RANDOM}};
  btb_10_pre_decoder_branchD_flag = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  btb_10_pre_decoder_jump = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  btb_10_pre_decoder_branchdata = _RAND_140[5:0];
  _RAND_141 = {1{`RANDOM}};
  btb_10_pre_decoder_jr = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  btb_10_true_branch_state = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  btb_11_pc = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  btb_11_inst = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  btb_11_exception_type = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  btb_11_pre_pc_target = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  btb_11_pre_lookup_data = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  btb_11_pre_hashcode = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  btb_11_pre_pht = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  btb_11_pre_bht = _RAND_150[6:0];
  _RAND_151 = {1{`RANDOM}};
  btb_11_pre_decoder_branchD_flag = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  btb_11_pre_decoder_jump = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  btb_11_pre_decoder_branchdata = _RAND_153[5:0];
  _RAND_154 = {1{`RANDOM}};
  btb_11_pre_decoder_jr = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  btb_11_true_branch_state = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  btb_12_pc = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  btb_12_inst = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  btb_12_exception_type = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  btb_12_pre_pc_target = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  btb_12_pre_lookup_data = _RAND_160[6:0];
  _RAND_161 = {1{`RANDOM}};
  btb_12_pre_hashcode = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  btb_12_pre_pht = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  btb_12_pre_bht = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  btb_12_pre_decoder_branchD_flag = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  btb_12_pre_decoder_jump = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  btb_12_pre_decoder_branchdata = _RAND_166[5:0];
  _RAND_167 = {1{`RANDOM}};
  btb_12_pre_decoder_jr = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  btb_12_true_branch_state = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  btb_13_pc = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  btb_13_inst = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  btb_13_exception_type = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  btb_13_pre_pc_target = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  btb_13_pre_lookup_data = _RAND_173[6:0];
  _RAND_174 = {1{`RANDOM}};
  btb_13_pre_hashcode = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  btb_13_pre_pht = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  btb_13_pre_bht = _RAND_176[6:0];
  _RAND_177 = {1{`RANDOM}};
  btb_13_pre_decoder_branchD_flag = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  btb_13_pre_decoder_jump = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  btb_13_pre_decoder_branchdata = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  btb_13_pre_decoder_jr = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  btb_13_true_branch_state = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  btb_14_pc = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  btb_14_inst = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  btb_14_exception_type = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  btb_14_pre_pc_target = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  btb_14_pre_lookup_data = _RAND_186[6:0];
  _RAND_187 = {1{`RANDOM}};
  btb_14_pre_hashcode = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  btb_14_pre_pht = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  btb_14_pre_bht = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  btb_14_pre_decoder_branchD_flag = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  btb_14_pre_decoder_jump = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  btb_14_pre_decoder_branchdata = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  btb_14_pre_decoder_jr = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  btb_14_true_branch_state = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  btb_15_pc = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  btb_15_inst = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  btb_15_exception_type = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  btb_15_pre_pc_target = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  btb_15_pre_lookup_data = _RAND_199[6:0];
  _RAND_200 = {1{`RANDOM}};
  btb_15_pre_hashcode = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  btb_15_pre_pht = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  btb_15_pre_bht = _RAND_202[6:0];
  _RAND_203 = {1{`RANDOM}};
  btb_15_pre_decoder_branchD_flag = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  btb_15_pre_decoder_jump = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  btb_15_pre_decoder_branchdata = _RAND_205[5:0];
  _RAND_206 = {1{`RANDOM}};
  btb_15_pre_decoder_jr = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  btb_15_true_branch_state = _RAND_207[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_fifo_with_bundle(
  input         clock,
  input         reset,
  input         io_read_en,
  input         io_write_en,
  output [31:0] io_read_out_0_pc,
  output [31:0] io_read_out_0_inst,
  output [1:0]  io_read_out_0_exception_type,
  output [31:0] io_read_out_0_pre_pc_target,
  output [6:0]  io_read_out_0_pre_lookup_data,
  output [3:0]  io_read_out_0_pre_hashcode,
  output [1:0]  io_read_out_0_pre_pht,
  output [6:0]  io_read_out_0_pre_bht,
  output        io_read_out_0_pre_decoder_branchD_flag,
  output        io_read_out_0_pre_decoder_jump,
  output [5:0]  io_read_out_0_pre_decoder_branchdata,
  output        io_read_out_0_pre_decoder_jr,
  output        io_read_out_0_true_branch_state,
  input  [31:0] io_write_in_0_pc,
  input  [31:0] io_write_in_0_inst,
  input  [31:0] io_write_in_0_pre_pc_target,
  input  [6:0]  io_write_in_0_pre_lookup_data,
  input  [3:0]  io_write_in_0_pre_hashcode,
  input  [1:0]  io_write_in_0_pre_pht,
  input  [6:0]  io_write_in_0_pre_bht,
  input         io_write_in_0_pre_decoder_branchD_flag,
  input         io_write_in_0_pre_decoder_jump,
  input  [5:0]  io_write_in_0_pre_decoder_branchdata,
  input         io_write_in_0_pre_decoder_jr,
  input         io_write_in_0_true_branch_state,
  output        io_full,
  output        io_empty,
  input         io_point_write_en,
  input         io_point_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  Look_up_table_read_first_with_bundle_clock; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_reset; // @[fifo.scala 118:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_ar_addr; // @[fifo.scala 118:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_aw_addr; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_write; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_in_pc; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_in_inst; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_in_pre_pc_target; // @[fifo.scala 118:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_in_pre_lookup_data; // @[fifo.scala 118:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_in_pre_hashcode; // @[fifo.scala 118:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_in_pre_pht; // @[fifo.scala 118:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_in_pre_bht; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump; // @[fifo.scala 118:55]
  wire [5:0] Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_in_true_branch_state; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_out_pc; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_out_inst; // @[fifo.scala 118:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_out_exception_type; // @[fifo.scala 118:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_out_pre_pc_target; // @[fifo.scala 118:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_out_pre_lookup_data; // @[fifo.scala 118:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_out_pre_hashcode; // @[fifo.scala 118:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_out_pre_pht; // @[fifo.scala 118:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_out_pre_bht; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump; // @[fifo.scala 118:55]
  wire [5:0] Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr; // @[fifo.scala 118:55]
  wire  Look_up_table_read_first_with_bundle_io_out_true_branch_state; // @[fifo.scala 118:55]
  reg [3:0] write_length_points; // @[fifo.scala 121:38]
  reg [3:0] read_length_points; // @[fifo.scala 123:37]
  wire [1:0] _GEN_0 = {{1'd0}, io_write_en}; // @[Mux.scala 81:61]
  wire  _write_length_points_T = io_point_flush | io_point_write_en; // @[fifo.scala 147:47]
  wire [2:0] _write_length_points_T_2 = {{1'd0}, _GEN_0}; // @[fifo.scala 147:134]
  wire [3:0] _GEN_3 = {{3'd0}, _write_length_points_T_2[0]}; // @[fifo.scala 147:93]
  wire [3:0] _write_length_points_T_7 = write_length_points + _GEN_3; // @[fifo.scala 147:93]
  wire [1:0] _GEN_4 = {{1'd0}, io_read_en}; // @[fifo.scala 149:131]
  wire [2:0] _read_length_points_T_2 = {{1'd0}, _GEN_4}; // @[fifo.scala 149:131]
  wire [3:0] _GEN_5 = {{3'd0}, _read_length_points_T_2[0]}; // @[fifo.scala 149:92]
  wire [3:0] _read_length_points_T_7 = read_length_points + _GEN_5; // @[fifo.scala 149:92]
  wire [31:0] fifo_banks_0_out_pc = Look_up_table_read_first_with_bundle_io_out_pc; // @[fifo.scala 118:{29,29}]
  wire [31:0] fifo_banks_0_out_inst = Look_up_table_read_first_with_bundle_io_out_inst; // @[fifo.scala 118:{29,29}]
  wire [1:0] fifo_banks_0_out_exception_type = Look_up_table_read_first_with_bundle_io_out_exception_type; // @[fifo.scala 118:{29,29}]
  wire [31:0] fifo_banks_0_out_pre_pc_target = Look_up_table_read_first_with_bundle_io_out_pre_pc_target; // @[fifo.scala 118:{29,29}]
  wire [6:0] fifo_banks_0_out_pre_lookup_data = Look_up_table_read_first_with_bundle_io_out_pre_lookup_data; // @[fifo.scala 118:{29,29}]
  wire [3:0] fifo_banks_0_out_pre_hashcode = Look_up_table_read_first_with_bundle_io_out_pre_hashcode; // @[fifo.scala 118:{29,29}]
  wire [1:0] fifo_banks_0_out_pre_pht = Look_up_table_read_first_with_bundle_io_out_pre_pht; // @[fifo.scala 118:{29,29}]
  wire [6:0] fifo_banks_0_out_pre_bht = Look_up_table_read_first_with_bundle_io_out_pre_bht; // @[fifo.scala 118:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_branchD_flag = Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag
    ; // @[fifo.scala 118:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_jump = Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump; // @[fifo.scala 118:{29,29}]
  wire [5:0] fifo_banks_0_out_pre_decoder_branchdata =
    Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata; // @[fifo.scala 118:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_jr = Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr; // @[fifo.scala 118:{29,29}]
  wire  fifo_banks_0_out_true_branch_state = Look_up_table_read_first_with_bundle_io_out_true_branch_state; // @[fifo.scala 118:{29,29}]
  wire [3:0] _io_full_T_1 = write_length_points + 4'h1; // @[fifo.scala 160:37]
  ysyx_22040886_Look_up_table_read_first_with_bundle Look_up_table_read_first_with_bundle ( // @[fifo.scala 118:55]
    .clock(Look_up_table_read_first_with_bundle_clock),
    .reset(Look_up_table_read_first_with_bundle_reset),
    .io_ar_addr(Look_up_table_read_first_with_bundle_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first_with_bundle_io_aw_addr),
    .io_write(Look_up_table_read_first_with_bundle_io_write),
    .io_in_pc(Look_up_table_read_first_with_bundle_io_in_pc),
    .io_in_inst(Look_up_table_read_first_with_bundle_io_in_inst),
    .io_in_pre_pc_target(Look_up_table_read_first_with_bundle_io_in_pre_pc_target),
    .io_in_pre_lookup_data(Look_up_table_read_first_with_bundle_io_in_pre_lookup_data),
    .io_in_pre_hashcode(Look_up_table_read_first_with_bundle_io_in_pre_hashcode),
    .io_in_pre_pht(Look_up_table_read_first_with_bundle_io_in_pre_pht),
    .io_in_pre_bht(Look_up_table_read_first_with_bundle_io_in_pre_bht),
    .io_in_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag),
    .io_in_pre_decoder_jump(Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump),
    .io_in_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata),
    .io_in_pre_decoder_jr(Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr),
    .io_in_true_branch_state(Look_up_table_read_first_with_bundle_io_in_true_branch_state),
    .io_out_pc(Look_up_table_read_first_with_bundle_io_out_pc),
    .io_out_inst(Look_up_table_read_first_with_bundle_io_out_inst),
    .io_out_exception_type(Look_up_table_read_first_with_bundle_io_out_exception_type),
    .io_out_pre_pc_target(Look_up_table_read_first_with_bundle_io_out_pre_pc_target),
    .io_out_pre_lookup_data(Look_up_table_read_first_with_bundle_io_out_pre_lookup_data),
    .io_out_pre_hashcode(Look_up_table_read_first_with_bundle_io_out_pre_hashcode),
    .io_out_pre_pht(Look_up_table_read_first_with_bundle_io_out_pre_pht),
    .io_out_pre_bht(Look_up_table_read_first_with_bundle_io_out_pre_bht),
    .io_out_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag),
    .io_out_pre_decoder_jump(Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump),
    .io_out_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata),
    .io_out_pre_decoder_jr(Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr),
    .io_out_true_branch_state(Look_up_table_read_first_with_bundle_io_out_true_branch_state)
  );
  assign io_read_out_0_pc = io_empty ? 32'h0 : fifo_banks_0_out_pc; // @[fifo.scala 151:30]
  assign io_read_out_0_inst = io_empty ? 32'h0 : fifo_banks_0_out_inst; // @[fifo.scala 151:30]
  assign io_read_out_0_exception_type = io_empty ? 2'h0 : fifo_banks_0_out_exception_type; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_pc_target = io_empty ? 32'h0 : fifo_banks_0_out_pre_pc_target; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_lookup_data = io_empty ? 7'h0 : fifo_banks_0_out_pre_lookup_data; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_hashcode = io_empty ? 4'h0 : fifo_banks_0_out_pre_hashcode; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_pht = io_empty ? 2'h0 : fifo_banks_0_out_pre_pht; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_bht = io_empty ? 7'h0 : fifo_banks_0_out_pre_bht; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_decoder_branchD_flag = io_empty ? 1'h0 : fifo_banks_0_out_pre_decoder_branchD_flag; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_decoder_jump = io_empty ? 1'h0 : fifo_banks_0_out_pre_decoder_jump; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_decoder_branchdata = io_empty ? 6'h0 : fifo_banks_0_out_pre_decoder_branchdata; // @[fifo.scala 151:30]
  assign io_read_out_0_pre_decoder_jr = io_empty ? 1'h0 : fifo_banks_0_out_pre_decoder_jr; // @[fifo.scala 151:30]
  assign io_read_out_0_true_branch_state = io_empty ? 1'h0 : fifo_banks_0_out_true_branch_state; // @[fifo.scala 151:30]
  assign io_full = _io_full_T_1 == read_length_points; // @[fifo.scala 160:43]
  assign io_empty = write_length_points == read_length_points | io_point_write_en; // @[fifo.scala 158:106]
  assign Look_up_table_read_first_with_bundle_clock = clock;
  assign Look_up_table_read_first_with_bundle_reset = reset;
  assign Look_up_table_read_first_with_bundle_io_ar_addr = read_length_points; // @[fifo.scala 118:29 128:38]
  assign Look_up_table_read_first_with_bundle_io_aw_addr = write_length_points; // @[fifo.scala 118:29 127:38]
  assign Look_up_table_read_first_with_bundle_io_write = io_write_en; // @[fifo.scala 132:28]
  assign Look_up_table_read_first_with_bundle_io_in_pc = io_write_in_0_pc; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_inst = io_write_in_0_inst; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_pc_target = io_write_in_0_pre_pc_target; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_lookup_data = io_write_in_0_pre_lookup_data; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_hashcode = io_write_in_0_pre_hashcode; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_pht = io_write_in_0_pre_pht; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_bht = io_write_in_0_pre_bht; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag = io_write_in_0_pre_decoder_branchD_flag; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump = io_write_in_0_pre_decoder_jump; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata = io_write_in_0_pre_decoder_branchdata; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr = io_write_in_0_pre_decoder_jr; // @[fifo.scala 118:29 129:38]
  assign Look_up_table_read_first_with_bundle_io_in_true_branch_state = io_write_in_0_true_branch_state; // @[fifo.scala 118:29 129:38]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 121:38]
      write_length_points <= 4'h0; // @[fifo.scala 121:38]
    end else if (io_point_flush | io_point_write_en) begin // @[fifo.scala 147:31]
      write_length_points <= 4'h0;
    end else begin
      write_length_points <= _write_length_points_T_7;
    end
    if (reset) begin // @[fifo.scala 123:37]
      read_length_points <= 4'h0; // @[fifo.scala 123:37]
    end else if (_write_length_points_T) begin // @[fifo.scala 149:30]
      read_length_points <= 4'h0;
    end else begin
      read_length_points <= _read_length_points_T_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  write_length_points = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  read_length_points = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_pc_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [31:0] io_in_pc_value_in,
  output [31:0] io_out_pc_value_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_value; // @[myCPU.scala 328:23]
  assign io_out_pc_value_out = pc_value; // @[myCPU.scala 331:25]
  always @(posedge clock) begin
    if (reset) begin // @[myCPU.scala 330:20]
      pc_value <= 32'h2ffffffc;
    end else if (io_flush) begin // @[myCPU.scala 330:60]
      pc_value <= 32'h0;
    end else if (io_stall) begin // @[myCPU.scala 330:77]
      pc_value <= io_in_pc_value_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_value = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_PHT(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [1:0] io_in,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] put_0; // @[PHTS.scala 18:22]
  reg [1:0] put_1; // @[PHTS.scala 18:22]
  reg [1:0] put_2; // @[PHTS.scala 18:22]
  reg [1:0] put_3; // @[PHTS.scala 18:22]
  reg [1:0] put_4; // @[PHTS.scala 18:22]
  reg [1:0] put_5; // @[PHTS.scala 18:22]
  reg [1:0] put_6; // @[PHTS.scala 18:22]
  reg [1:0] put_7; // @[PHTS.scala 18:22]
  reg [1:0] put_8; // @[PHTS.scala 18:22]
  reg [1:0] put_9; // @[PHTS.scala 18:22]
  reg [1:0] put_10; // @[PHTS.scala 18:22]
  reg [1:0] put_11; // @[PHTS.scala 18:22]
  reg [1:0] put_12; // @[PHTS.scala 18:22]
  reg [1:0] put_13; // @[PHTS.scala 18:22]
  reg [1:0] put_14; // @[PHTS.scala 18:22]
  reg [1:0] put_15; // @[PHTS.scala 18:22]
  reg [1:0] put_16; // @[PHTS.scala 18:22]
  reg [1:0] put_17; // @[PHTS.scala 18:22]
  reg [1:0] put_18; // @[PHTS.scala 18:22]
  reg [1:0] put_19; // @[PHTS.scala 18:22]
  reg [1:0] put_20; // @[PHTS.scala 18:22]
  reg [1:0] put_21; // @[PHTS.scala 18:22]
  reg [1:0] put_22; // @[PHTS.scala 18:22]
  reg [1:0] put_23; // @[PHTS.scala 18:22]
  reg [1:0] put_24; // @[PHTS.scala 18:22]
  reg [1:0] put_25; // @[PHTS.scala 18:22]
  reg [1:0] put_26; // @[PHTS.scala 18:22]
  reg [1:0] put_27; // @[PHTS.scala 18:22]
  reg [1:0] put_28; // @[PHTS.scala 18:22]
  reg [1:0] put_29; // @[PHTS.scala 18:22]
  reg [1:0] put_30; // @[PHTS.scala 18:22]
  reg [1:0] put_31; // @[PHTS.scala 18:22]
  reg [1:0] put_32; // @[PHTS.scala 18:22]
  reg [1:0] put_33; // @[PHTS.scala 18:22]
  reg [1:0] put_34; // @[PHTS.scala 18:22]
  reg [1:0] put_35; // @[PHTS.scala 18:22]
  reg [1:0] put_36; // @[PHTS.scala 18:22]
  reg [1:0] put_37; // @[PHTS.scala 18:22]
  reg [1:0] put_38; // @[PHTS.scala 18:22]
  reg [1:0] put_39; // @[PHTS.scala 18:22]
  reg [1:0] put_40; // @[PHTS.scala 18:22]
  reg [1:0] put_41; // @[PHTS.scala 18:22]
  reg [1:0] put_42; // @[PHTS.scala 18:22]
  reg [1:0] put_43; // @[PHTS.scala 18:22]
  reg [1:0] put_44; // @[PHTS.scala 18:22]
  reg [1:0] put_45; // @[PHTS.scala 18:22]
  reg [1:0] put_46; // @[PHTS.scala 18:22]
  reg [1:0] put_47; // @[PHTS.scala 18:22]
  reg [1:0] put_48; // @[PHTS.scala 18:22]
  reg [1:0] put_49; // @[PHTS.scala 18:22]
  reg [1:0] put_50; // @[PHTS.scala 18:22]
  reg [1:0] put_51; // @[PHTS.scala 18:22]
  reg [1:0] put_52; // @[PHTS.scala 18:22]
  reg [1:0] put_53; // @[PHTS.scala 18:22]
  reg [1:0] put_54; // @[PHTS.scala 18:22]
  reg [1:0] put_55; // @[PHTS.scala 18:22]
  reg [1:0] put_56; // @[PHTS.scala 18:22]
  reg [1:0] put_57; // @[PHTS.scala 18:22]
  reg [1:0] put_58; // @[PHTS.scala 18:22]
  reg [1:0] put_59; // @[PHTS.scala 18:22]
  reg [1:0] put_60; // @[PHTS.scala 18:22]
  reg [1:0] put_61; // @[PHTS.scala 18:22]
  reg [1:0] put_62; // @[PHTS.scala 18:22]
  reg [1:0] put_63; // @[PHTS.scala 18:22]
  reg [1:0] put_64; // @[PHTS.scala 18:22]
  reg [1:0] put_65; // @[PHTS.scala 18:22]
  reg [1:0] put_66; // @[PHTS.scala 18:22]
  reg [1:0] put_67; // @[PHTS.scala 18:22]
  reg [1:0] put_68; // @[PHTS.scala 18:22]
  reg [1:0] put_69; // @[PHTS.scala 18:22]
  reg [1:0] put_70; // @[PHTS.scala 18:22]
  reg [1:0] put_71; // @[PHTS.scala 18:22]
  reg [1:0] put_72; // @[PHTS.scala 18:22]
  reg [1:0] put_73; // @[PHTS.scala 18:22]
  reg [1:0] put_74; // @[PHTS.scala 18:22]
  reg [1:0] put_75; // @[PHTS.scala 18:22]
  reg [1:0] put_76; // @[PHTS.scala 18:22]
  reg [1:0] put_77; // @[PHTS.scala 18:22]
  reg [1:0] put_78; // @[PHTS.scala 18:22]
  reg [1:0] put_79; // @[PHTS.scala 18:22]
  reg [1:0] put_80; // @[PHTS.scala 18:22]
  reg [1:0] put_81; // @[PHTS.scala 18:22]
  reg [1:0] put_82; // @[PHTS.scala 18:22]
  reg [1:0] put_83; // @[PHTS.scala 18:22]
  reg [1:0] put_84; // @[PHTS.scala 18:22]
  reg [1:0] put_85; // @[PHTS.scala 18:22]
  reg [1:0] put_86; // @[PHTS.scala 18:22]
  reg [1:0] put_87; // @[PHTS.scala 18:22]
  reg [1:0] put_88; // @[PHTS.scala 18:22]
  reg [1:0] put_89; // @[PHTS.scala 18:22]
  reg [1:0] put_90; // @[PHTS.scala 18:22]
  reg [1:0] put_91; // @[PHTS.scala 18:22]
  reg [1:0] put_92; // @[PHTS.scala 18:22]
  reg [1:0] put_93; // @[PHTS.scala 18:22]
  reg [1:0] put_94; // @[PHTS.scala 18:22]
  reg [1:0] put_95; // @[PHTS.scala 18:22]
  reg [1:0] put_96; // @[PHTS.scala 18:22]
  reg [1:0] put_97; // @[PHTS.scala 18:22]
  reg [1:0] put_98; // @[PHTS.scala 18:22]
  reg [1:0] put_99; // @[PHTS.scala 18:22]
  reg [1:0] put_100; // @[PHTS.scala 18:22]
  reg [1:0] put_101; // @[PHTS.scala 18:22]
  reg [1:0] put_102; // @[PHTS.scala 18:22]
  reg [1:0] put_103; // @[PHTS.scala 18:22]
  reg [1:0] put_104; // @[PHTS.scala 18:22]
  reg [1:0] put_105; // @[PHTS.scala 18:22]
  reg [1:0] put_106; // @[PHTS.scala 18:22]
  reg [1:0] put_107; // @[PHTS.scala 18:22]
  reg [1:0] put_108; // @[PHTS.scala 18:22]
  reg [1:0] put_109; // @[PHTS.scala 18:22]
  reg [1:0] put_110; // @[PHTS.scala 18:22]
  reg [1:0] put_111; // @[PHTS.scala 18:22]
  reg [1:0] put_112; // @[PHTS.scala 18:22]
  reg [1:0] put_113; // @[PHTS.scala 18:22]
  reg [1:0] put_114; // @[PHTS.scala 18:22]
  reg [1:0] put_115; // @[PHTS.scala 18:22]
  reg [1:0] put_116; // @[PHTS.scala 18:22]
  reg [1:0] put_117; // @[PHTS.scala 18:22]
  reg [1:0] put_118; // @[PHTS.scala 18:22]
  reg [1:0] put_119; // @[PHTS.scala 18:22]
  reg [1:0] put_120; // @[PHTS.scala 18:22]
  reg [1:0] put_121; // @[PHTS.scala 18:22]
  reg [1:0] put_122; // @[PHTS.scala 18:22]
  reg [1:0] put_123; // @[PHTS.scala 18:22]
  reg [1:0] put_124; // @[PHTS.scala 18:22]
  reg [1:0] put_125; // @[PHTS.scala 18:22]
  reg [1:0] put_126; // @[PHTS.scala 18:22]
  reg [1:0] put_127; // @[PHTS.scala 18:22]
  wire [1:0] _GEN_1 = 7'h1 == io_ar_addr ? put_1 : put_0; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_2 = 7'h2 == io_ar_addr ? put_2 : _GEN_1; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_3 = 7'h3 == io_ar_addr ? put_3 : _GEN_2; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_4 = 7'h4 == io_ar_addr ? put_4 : _GEN_3; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_5 = 7'h5 == io_ar_addr ? put_5 : _GEN_4; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_6 = 7'h6 == io_ar_addr ? put_6 : _GEN_5; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_7 = 7'h7 == io_ar_addr ? put_7 : _GEN_6; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_8 = 7'h8 == io_ar_addr ? put_8 : _GEN_7; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_9 = 7'h9 == io_ar_addr ? put_9 : _GEN_8; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_10 = 7'ha == io_ar_addr ? put_10 : _GEN_9; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_11 = 7'hb == io_ar_addr ? put_11 : _GEN_10; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_12 = 7'hc == io_ar_addr ? put_12 : _GEN_11; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_13 = 7'hd == io_ar_addr ? put_13 : _GEN_12; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_14 = 7'he == io_ar_addr ? put_14 : _GEN_13; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_15 = 7'hf == io_ar_addr ? put_15 : _GEN_14; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_16 = 7'h10 == io_ar_addr ? put_16 : _GEN_15; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_17 = 7'h11 == io_ar_addr ? put_17 : _GEN_16; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_18 = 7'h12 == io_ar_addr ? put_18 : _GEN_17; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_19 = 7'h13 == io_ar_addr ? put_19 : _GEN_18; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_20 = 7'h14 == io_ar_addr ? put_20 : _GEN_19; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_21 = 7'h15 == io_ar_addr ? put_21 : _GEN_20; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_22 = 7'h16 == io_ar_addr ? put_22 : _GEN_21; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_23 = 7'h17 == io_ar_addr ? put_23 : _GEN_22; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_24 = 7'h18 == io_ar_addr ? put_24 : _GEN_23; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_25 = 7'h19 == io_ar_addr ? put_25 : _GEN_24; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_26 = 7'h1a == io_ar_addr ? put_26 : _GEN_25; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_27 = 7'h1b == io_ar_addr ? put_27 : _GEN_26; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_28 = 7'h1c == io_ar_addr ? put_28 : _GEN_27; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_29 = 7'h1d == io_ar_addr ? put_29 : _GEN_28; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_30 = 7'h1e == io_ar_addr ? put_30 : _GEN_29; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_31 = 7'h1f == io_ar_addr ? put_31 : _GEN_30; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_32 = 7'h20 == io_ar_addr ? put_32 : _GEN_31; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_33 = 7'h21 == io_ar_addr ? put_33 : _GEN_32; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_34 = 7'h22 == io_ar_addr ? put_34 : _GEN_33; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_35 = 7'h23 == io_ar_addr ? put_35 : _GEN_34; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_36 = 7'h24 == io_ar_addr ? put_36 : _GEN_35; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_37 = 7'h25 == io_ar_addr ? put_37 : _GEN_36; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_38 = 7'h26 == io_ar_addr ? put_38 : _GEN_37; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_39 = 7'h27 == io_ar_addr ? put_39 : _GEN_38; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_40 = 7'h28 == io_ar_addr ? put_40 : _GEN_39; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_41 = 7'h29 == io_ar_addr ? put_41 : _GEN_40; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_42 = 7'h2a == io_ar_addr ? put_42 : _GEN_41; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_43 = 7'h2b == io_ar_addr ? put_43 : _GEN_42; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_44 = 7'h2c == io_ar_addr ? put_44 : _GEN_43; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_45 = 7'h2d == io_ar_addr ? put_45 : _GEN_44; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_46 = 7'h2e == io_ar_addr ? put_46 : _GEN_45; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_47 = 7'h2f == io_ar_addr ? put_47 : _GEN_46; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_48 = 7'h30 == io_ar_addr ? put_48 : _GEN_47; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_49 = 7'h31 == io_ar_addr ? put_49 : _GEN_48; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_50 = 7'h32 == io_ar_addr ? put_50 : _GEN_49; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_51 = 7'h33 == io_ar_addr ? put_51 : _GEN_50; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_52 = 7'h34 == io_ar_addr ? put_52 : _GEN_51; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_53 = 7'h35 == io_ar_addr ? put_53 : _GEN_52; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_54 = 7'h36 == io_ar_addr ? put_54 : _GEN_53; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_55 = 7'h37 == io_ar_addr ? put_55 : _GEN_54; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_56 = 7'h38 == io_ar_addr ? put_56 : _GEN_55; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_57 = 7'h39 == io_ar_addr ? put_57 : _GEN_56; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_58 = 7'h3a == io_ar_addr ? put_58 : _GEN_57; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_59 = 7'h3b == io_ar_addr ? put_59 : _GEN_58; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_60 = 7'h3c == io_ar_addr ? put_60 : _GEN_59; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_61 = 7'h3d == io_ar_addr ? put_61 : _GEN_60; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_62 = 7'h3e == io_ar_addr ? put_62 : _GEN_61; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_63 = 7'h3f == io_ar_addr ? put_63 : _GEN_62; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_64 = 7'h40 == io_ar_addr ? put_64 : _GEN_63; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_65 = 7'h41 == io_ar_addr ? put_65 : _GEN_64; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_66 = 7'h42 == io_ar_addr ? put_66 : _GEN_65; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_67 = 7'h43 == io_ar_addr ? put_67 : _GEN_66; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_68 = 7'h44 == io_ar_addr ? put_68 : _GEN_67; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_69 = 7'h45 == io_ar_addr ? put_69 : _GEN_68; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_70 = 7'h46 == io_ar_addr ? put_70 : _GEN_69; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_71 = 7'h47 == io_ar_addr ? put_71 : _GEN_70; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_72 = 7'h48 == io_ar_addr ? put_72 : _GEN_71; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_73 = 7'h49 == io_ar_addr ? put_73 : _GEN_72; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_74 = 7'h4a == io_ar_addr ? put_74 : _GEN_73; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_75 = 7'h4b == io_ar_addr ? put_75 : _GEN_74; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_76 = 7'h4c == io_ar_addr ? put_76 : _GEN_75; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_77 = 7'h4d == io_ar_addr ? put_77 : _GEN_76; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_78 = 7'h4e == io_ar_addr ? put_78 : _GEN_77; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_79 = 7'h4f == io_ar_addr ? put_79 : _GEN_78; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_80 = 7'h50 == io_ar_addr ? put_80 : _GEN_79; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_81 = 7'h51 == io_ar_addr ? put_81 : _GEN_80; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_82 = 7'h52 == io_ar_addr ? put_82 : _GEN_81; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_83 = 7'h53 == io_ar_addr ? put_83 : _GEN_82; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_84 = 7'h54 == io_ar_addr ? put_84 : _GEN_83; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_85 = 7'h55 == io_ar_addr ? put_85 : _GEN_84; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_86 = 7'h56 == io_ar_addr ? put_86 : _GEN_85; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_87 = 7'h57 == io_ar_addr ? put_87 : _GEN_86; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_88 = 7'h58 == io_ar_addr ? put_88 : _GEN_87; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_89 = 7'h59 == io_ar_addr ? put_89 : _GEN_88; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_90 = 7'h5a == io_ar_addr ? put_90 : _GEN_89; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_91 = 7'h5b == io_ar_addr ? put_91 : _GEN_90; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_92 = 7'h5c == io_ar_addr ? put_92 : _GEN_91; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_93 = 7'h5d == io_ar_addr ? put_93 : _GEN_92; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_94 = 7'h5e == io_ar_addr ? put_94 : _GEN_93; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_95 = 7'h5f == io_ar_addr ? put_95 : _GEN_94; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_96 = 7'h60 == io_ar_addr ? put_96 : _GEN_95; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_97 = 7'h61 == io_ar_addr ? put_97 : _GEN_96; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_98 = 7'h62 == io_ar_addr ? put_98 : _GEN_97; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_99 = 7'h63 == io_ar_addr ? put_99 : _GEN_98; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_100 = 7'h64 == io_ar_addr ? put_100 : _GEN_99; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_101 = 7'h65 == io_ar_addr ? put_101 : _GEN_100; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_102 = 7'h66 == io_ar_addr ? put_102 : _GEN_101; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_103 = 7'h67 == io_ar_addr ? put_103 : _GEN_102; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_104 = 7'h68 == io_ar_addr ? put_104 : _GEN_103; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_105 = 7'h69 == io_ar_addr ? put_105 : _GEN_104; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_106 = 7'h6a == io_ar_addr ? put_106 : _GEN_105; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_107 = 7'h6b == io_ar_addr ? put_107 : _GEN_106; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_108 = 7'h6c == io_ar_addr ? put_108 : _GEN_107; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_109 = 7'h6d == io_ar_addr ? put_109 : _GEN_108; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_110 = 7'h6e == io_ar_addr ? put_110 : _GEN_109; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_111 = 7'h6f == io_ar_addr ? put_111 : _GEN_110; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_112 = 7'h70 == io_ar_addr ? put_112 : _GEN_111; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_113 = 7'h71 == io_ar_addr ? put_113 : _GEN_112; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_114 = 7'h72 == io_ar_addr ? put_114 : _GEN_113; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_115 = 7'h73 == io_ar_addr ? put_115 : _GEN_114; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_116 = 7'h74 == io_ar_addr ? put_116 : _GEN_115; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_117 = 7'h75 == io_ar_addr ? put_117 : _GEN_116; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_118 = 7'h76 == io_ar_addr ? put_118 : _GEN_117; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_119 = 7'h77 == io_ar_addr ? put_119 : _GEN_118; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_120 = 7'h78 == io_ar_addr ? put_120 : _GEN_119; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_121 = 7'h79 == io_ar_addr ? put_121 : _GEN_120; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_122 = 7'h7a == io_ar_addr ? put_122 : _GEN_121; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_123 = 7'h7b == io_ar_addr ? put_123 : _GEN_122; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_124 = 7'h7c == io_ar_addr ? put_124 : _GEN_123; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_125 = 7'h7d == io_ar_addr ? put_125 : _GEN_124; // @[PHTS.scala 19:{12,12}]
  wire [1:0] _GEN_126 = 7'h7e == io_ar_addr ? put_126 : _GEN_125; // @[PHTS.scala 19:{12,12}]
  assign io_out = 7'h7f == io_ar_addr ? put_127 : _GEN_126; // @[PHTS.scala 19:{12,12}]
  always @(posedge clock) begin
    if (reset) begin // @[PHTS.scala 18:22]
      put_0 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h0 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_0 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_1 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_1 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_2 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_2 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_3 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_3 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_4 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_4 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_5 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_5 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_6 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_6 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_7 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_7 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_8 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h8 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_8 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_9 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h9 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_9 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_10 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'ha == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_10 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_11 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'hb == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_11 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_12 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'hc == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_12 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_13 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'hd == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_13 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_14 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'he == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_14 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_15 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'hf == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_15 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_16 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h10 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_16 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_17 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h11 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_17 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_18 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h12 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_18 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_19 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h13 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_19 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_20 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h14 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_20 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_21 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h15 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_21 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_22 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h16 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_22 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_23 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h17 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_23 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_24 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h18 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_24 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_25 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h19 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_25 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_26 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_26 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_27 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_27 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_28 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_28 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_29 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_29 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_30 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_30 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_31 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h1f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_31 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_32 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h20 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_32 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_33 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h21 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_33 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_34 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h22 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_34 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_35 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h23 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_35 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_36 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h24 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_36 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_37 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h25 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_37 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_38 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h26 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_38 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_39 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h27 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_39 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_40 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h28 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_40 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_41 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h29 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_41 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_42 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_42 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_43 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_43 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_44 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_44 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_45 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_45 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_46 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_46 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_47 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h2f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_47 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_48 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h30 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_48 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_49 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h31 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_49 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_50 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h32 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_50 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_51 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h33 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_51 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_52 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h34 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_52 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_53 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h35 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_53 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_54 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h36 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_54 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_55 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h37 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_55 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_56 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h38 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_56 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_57 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h39 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_57 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_58 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_58 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_59 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_59 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_60 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_60 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_61 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_61 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_62 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_62 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_63 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h3f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_63 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_64 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h40 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_64 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_65 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h41 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_65 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_66 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h42 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_66 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_67 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h43 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_67 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_68 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h44 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_68 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_69 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h45 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_69 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_70 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h46 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_70 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_71 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h47 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_71 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_72 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h48 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_72 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_73 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h49 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_73 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_74 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_74 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_75 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_75 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_76 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_76 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_77 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_77 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_78 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_78 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_79 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h4f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_79 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_80 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h50 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_80 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_81 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h51 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_81 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_82 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h52 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_82 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_83 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h53 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_83 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_84 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h54 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_84 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_85 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h55 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_85 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_86 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h56 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_86 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_87 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h57 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_87 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_88 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h58 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_88 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_89 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h59 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_89 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_90 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_90 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_91 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_91 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_92 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_92 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_93 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_93 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_94 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_94 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_95 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h5f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_95 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_96 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h60 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_96 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_97 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h61 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_97 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_98 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h62 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_98 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_99 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h63 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_99 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_100 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h64 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_100 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_101 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h65 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_101 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_102 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h66 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_102 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_103 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h67 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_103 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_104 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h68 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_104 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_105 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h69 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_105 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_106 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_106 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_107 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_107 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_108 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_108 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_109 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_109 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_110 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_110 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_111 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h6f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_111 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_112 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h70 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_112 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_113 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h71 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_113 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_114 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h72 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_114 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_115 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h73 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_115 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_116 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h74 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_116 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_117 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h75 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_117 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_118 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h76 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_118 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_119 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h77 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_119 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_120 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h78 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_120 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_121 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h79 == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_121 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_122 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7a == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_122 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_123 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7b == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_123 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_124 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7c == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_124 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_125 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7d == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_125 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_126 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7e == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_126 <= io_in;
    end
    if (reset) begin // @[PHTS.scala 18:22]
      put_127 <= 2'h0; // @[PHTS.scala 18:22]
    end else if (io_write & 7'h7f == io_aw_addr) begin // @[PHTS.scala 22:22]
      put_127 <= io_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  put_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  put_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  put_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  put_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  put_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  put_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  put_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  put_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  put_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  put_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  put_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  put_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  put_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  put_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  put_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  put_15 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  put_16 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  put_17 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  put_18 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  put_19 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  put_20 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  put_21 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  put_22 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  put_23 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  put_24 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  put_25 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  put_26 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  put_27 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  put_28 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  put_29 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  put_30 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  put_31 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  put_32 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  put_33 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  put_34 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  put_35 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  put_36 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  put_37 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  put_38 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  put_39 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  put_40 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  put_41 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  put_42 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  put_43 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  put_44 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  put_45 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  put_46 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  put_47 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  put_48 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  put_49 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  put_50 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  put_51 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  put_52 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  put_53 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  put_54 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  put_55 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  put_56 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  put_57 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  put_58 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  put_59 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  put_60 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  put_61 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  put_62 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  put_63 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  put_64 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  put_65 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  put_66 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  put_67 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  put_68 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  put_69 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  put_70 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  put_71 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  put_72 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  put_73 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  put_74 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  put_75 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  put_76 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  put_77 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  put_78 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  put_79 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  put_80 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  put_81 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  put_82 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  put_83 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  put_84 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  put_85 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  put_86 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  put_87 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  put_88 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  put_89 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  put_90 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  put_91 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  put_92 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  put_93 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  put_94 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  put_95 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  put_96 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  put_97 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  put_98 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  put_99 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  put_100 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  put_101 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  put_102 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  put_103 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  put_104 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  put_105 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  put_106 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  put_107 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  put_108 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  put_109 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  put_110 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  put_111 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  put_112 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  put_113 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  put_114 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  put_115 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  put_116 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  put_117 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  put_118 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  put_119 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  put_120 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  put_121 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  put_122 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  put_123 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  put_124 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  put_125 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  put_126 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  put_127 = _RAND_127[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_PHTS(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [1:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [1:0] io_aw_pht_addr,
  input        io_write,
  input  [1:0] io_in,
  output [1:0] io_out
);
  wire  PHT_clock; // @[PHTS.scala 42:45]
  wire  PHT_reset; // @[PHTS.scala 42:45]
  wire [6:0] PHT_io_ar_addr; // @[PHTS.scala 42:45]
  wire [6:0] PHT_io_aw_addr; // @[PHTS.scala 42:45]
  wire  PHT_io_write; // @[PHTS.scala 42:45]
  wire [1:0] PHT_io_in; // @[PHTS.scala 42:45]
  wire [1:0] PHT_io_out; // @[PHTS.scala 42:45]
  wire  PHT_1_clock; // @[PHTS.scala 42:45]
  wire  PHT_1_reset; // @[PHTS.scala 42:45]
  wire [6:0] PHT_1_io_ar_addr; // @[PHTS.scala 42:45]
  wire [6:0] PHT_1_io_aw_addr; // @[PHTS.scala 42:45]
  wire  PHT_1_io_write; // @[PHTS.scala 42:45]
  wire [1:0] PHT_1_io_in; // @[PHTS.scala 42:45]
  wire [1:0] PHT_1_io_out; // @[PHTS.scala 42:45]
  wire  PHT_2_clock; // @[PHTS.scala 42:45]
  wire  PHT_2_reset; // @[PHTS.scala 42:45]
  wire [6:0] PHT_2_io_ar_addr; // @[PHTS.scala 42:45]
  wire [6:0] PHT_2_io_aw_addr; // @[PHTS.scala 42:45]
  wire  PHT_2_io_write; // @[PHTS.scala 42:45]
  wire [1:0] PHT_2_io_in; // @[PHTS.scala 42:45]
  wire [1:0] PHT_2_io_out; // @[PHTS.scala 42:45]
  wire  PHT_3_clock; // @[PHTS.scala 42:45]
  wire  PHT_3_reset; // @[PHTS.scala 42:45]
  wire [6:0] PHT_3_io_ar_addr; // @[PHTS.scala 42:45]
  wire [6:0] PHT_3_io_aw_addr; // @[PHTS.scala 42:45]
  wire  PHT_3_io_write; // @[PHTS.scala 42:45]
  wire [1:0] PHT_3_io_in; // @[PHTS.scala 42:45]
  wire [1:0] PHT_3_io_out; // @[PHTS.scala 42:45]
  wire [1:0] phts_0_out = PHT_io_out; // @[PHTS.scala 42:{23,23}]
  wire [1:0] phts_1_out = PHT_1_io_out; // @[PHTS.scala 42:{23,23}]
  wire [1:0] _GEN_1 = 2'h1 == io_ar_pht_addr ? phts_1_out : phts_0_out; // @[PHTS.scala 49:{12,12}]
  wire [1:0] phts_2_out = PHT_2_io_out; // @[PHTS.scala 42:{23,23}]
  wire [1:0] _GEN_2 = 2'h2 == io_ar_pht_addr ? phts_2_out : _GEN_1; // @[PHTS.scala 49:{12,12}]
  wire [1:0] phts_3_out = PHT_3_io_out; // @[PHTS.scala 42:{23,23}]
  ysyx_22040886_PHT PHT ( // @[PHTS.scala 42:45]
    .clock(PHT_clock),
    .reset(PHT_reset),
    .io_ar_addr(PHT_io_ar_addr),
    .io_aw_addr(PHT_io_aw_addr),
    .io_write(PHT_io_write),
    .io_in(PHT_io_in),
    .io_out(PHT_io_out)
  );
  ysyx_22040886_PHT PHT_1 ( // @[PHTS.scala 42:45]
    .clock(PHT_1_clock),
    .reset(PHT_1_reset),
    .io_ar_addr(PHT_1_io_ar_addr),
    .io_aw_addr(PHT_1_io_aw_addr),
    .io_write(PHT_1_io_write),
    .io_in(PHT_1_io_in),
    .io_out(PHT_1_io_out)
  );
  ysyx_22040886_PHT PHT_2 ( // @[PHTS.scala 42:45]
    .clock(PHT_2_clock),
    .reset(PHT_2_reset),
    .io_ar_addr(PHT_2_io_ar_addr),
    .io_aw_addr(PHT_2_io_aw_addr),
    .io_write(PHT_2_io_write),
    .io_in(PHT_2_io_in),
    .io_out(PHT_2_io_out)
  );
  ysyx_22040886_PHT PHT_3 ( // @[PHTS.scala 42:45]
    .clock(PHT_3_clock),
    .reset(PHT_3_reset),
    .io_ar_addr(PHT_3_io_ar_addr),
    .io_aw_addr(PHT_3_io_aw_addr),
    .io_write(PHT_3_io_write),
    .io_in(PHT_3_io_in),
    .io_out(PHT_3_io_out)
  );
  assign io_out = 2'h3 == io_ar_pht_addr ? phts_3_out : _GEN_2; // @[PHTS.scala 49:{12,12}]
  assign PHT_clock = clock;
  assign PHT_reset = reset;
  assign PHT_io_ar_addr = io_ar_addr; // @[PHTS.scala 42:23 46:25]
  assign PHT_io_aw_addr = io_aw_addr; // @[PHTS.scala 42:23 47:25]
  assign PHT_io_write = io_aw_pht_addr == 2'h0 & io_write; // @[PHTS.scala 44:54]
  assign PHT_io_in = io_in; // @[PHTS.scala 42:23 45:20]
  assign PHT_1_clock = clock;
  assign PHT_1_reset = reset;
  assign PHT_1_io_ar_addr = io_ar_addr; // @[PHTS.scala 42:23 46:25]
  assign PHT_1_io_aw_addr = io_aw_addr; // @[PHTS.scala 42:23 47:25]
  assign PHT_1_io_write = io_aw_pht_addr == 2'h1 & io_write; // @[PHTS.scala 44:54]
  assign PHT_1_io_in = io_in; // @[PHTS.scala 42:23 45:20]
  assign PHT_2_clock = clock;
  assign PHT_2_reset = reset;
  assign PHT_2_io_ar_addr = io_ar_addr; // @[PHTS.scala 42:23 46:25]
  assign PHT_2_io_aw_addr = io_aw_addr; // @[PHTS.scala 42:23 47:25]
  assign PHT_2_io_write = io_aw_pht_addr == 2'h2 & io_write; // @[PHTS.scala 44:54]
  assign PHT_2_io_in = io_in; // @[PHTS.scala 42:23 45:20]
  assign PHT_3_clock = clock;
  assign PHT_3_reset = reset;
  assign PHT_3_io_ar_addr = io_ar_addr; // @[PHTS.scala 42:23 46:25]
  assign PHT_3_io_aw_addr = io_aw_addr; // @[PHTS.scala 42:23 47:25]
  assign PHT_3_io_write = io_aw_pht_addr == 2'h3 & io_write; // @[PHTS.scala 44:54]
  assign PHT_3_io_in = io_in; // @[PHTS.scala 42:23 45:20]
endmodule
module ysyx_22040886_PHTS_banks_oneissue(
  input        clock,
  input        reset,
  input        io_ar_bank_sel,
  input  [6:0] io_ar_addr,
  input  [1:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [1:0] io_aw_pht_addr,
  input        io_aw_bank_sel,
  input        io_write,
  input  [1:0] io_in,
  output [1:0] io_out
);
  wire  PHTS_clock; // @[PHTS.scala 122:55]
  wire  PHTS_reset; // @[PHTS.scala 122:55]
  wire [6:0] PHTS_io_ar_addr; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_io_ar_pht_addr; // @[PHTS.scala 122:55]
  wire [6:0] PHTS_io_aw_addr; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_io_aw_pht_addr; // @[PHTS.scala 122:55]
  wire  PHTS_io_write; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_io_in; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_io_out; // @[PHTS.scala 122:55]
  wire  PHTS_1_clock; // @[PHTS.scala 122:55]
  wire  PHTS_1_reset; // @[PHTS.scala 122:55]
  wire [6:0] PHTS_1_io_ar_addr; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_1_io_ar_pht_addr; // @[PHTS.scala 122:55]
  wire [6:0] PHTS_1_io_aw_addr; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_1_io_aw_pht_addr; // @[PHTS.scala 122:55]
  wire  PHTS_1_io_write; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_1_io_in; // @[PHTS.scala 122:55]
  wire [1:0] PHTS_1_io_out; // @[PHTS.scala 122:55]
  wire [1:0] phts_banks_0_out = PHTS_io_out; // @[PHTS.scala 122:{29,29}]
  wire [1:0] phts_banks_1_out = PHTS_1_io_out; // @[PHTS.scala 122:{29,29}]
  ysyx_22040886_PHTS PHTS ( // @[PHTS.scala 122:55]
    .clock(PHTS_clock),
    .reset(PHTS_reset),
    .io_ar_addr(PHTS_io_ar_addr),
    .io_ar_pht_addr(PHTS_io_ar_pht_addr),
    .io_aw_addr(PHTS_io_aw_addr),
    .io_aw_pht_addr(PHTS_io_aw_pht_addr),
    .io_write(PHTS_io_write),
    .io_in(PHTS_io_in),
    .io_out(PHTS_io_out)
  );
  ysyx_22040886_PHTS PHTS_1 ( // @[PHTS.scala 122:55]
    .clock(PHTS_1_clock),
    .reset(PHTS_1_reset),
    .io_ar_addr(PHTS_1_io_ar_addr),
    .io_ar_pht_addr(PHTS_1_io_ar_pht_addr),
    .io_aw_addr(PHTS_1_io_aw_addr),
    .io_aw_pht_addr(PHTS_1_io_aw_pht_addr),
    .io_write(PHTS_1_io_write),
    .io_in(PHTS_1_io_in),
    .io_out(PHTS_1_io_out)
  );
  assign io_out = io_ar_bank_sel ? phts_banks_1_out : phts_banks_0_out; // @[PHTS.scala 133:{12,12}]
  assign PHTS_clock = clock;
  assign PHTS_reset = reset;
  assign PHTS_io_ar_addr = io_ar_addr; // @[PHTS.scala 122:29 126:31]
  assign PHTS_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 122:29 129:35]
  assign PHTS_io_aw_addr = io_aw_addr; // @[PHTS.scala 122:29 130:31]
  assign PHTS_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 122:29 131:35]
  assign PHTS_io_write = ~io_aw_bank_sel & io_write; // @[PHTS.scala 124:60]
  assign PHTS_io_in = io_in; // @[PHTS.scala 122:29 125:26]
  assign PHTS_1_clock = clock;
  assign PHTS_1_reset = reset;
  assign PHTS_1_io_ar_addr = io_ar_addr; // @[PHTS.scala 122:29 126:31]
  assign PHTS_1_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 122:29 129:35]
  assign PHTS_1_io_aw_addr = io_aw_addr; // @[PHTS.scala 122:29 130:31]
  assign PHTS_1_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 122:29 131:35]
  assign PHTS_1_io_write = io_aw_bank_sel & io_write; // @[PHTS.scala 124:60]
  assign PHTS_1_io_in = io_in; // @[PHTS.scala 122:29 125:26]
endmodule
module ysyx_22040886_BHT(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] bht_0; // @[BHT.scala 20:22]
  reg [2:0] bht_1; // @[BHT.scala 20:22]
  reg [2:0] bht_2; // @[BHT.scala 20:22]
  reg [2:0] bht_3; // @[BHT.scala 20:22]
  reg [2:0] bht_4; // @[BHT.scala 20:22]
  reg [2:0] bht_5; // @[BHT.scala 20:22]
  reg [2:0] bht_6; // @[BHT.scala 20:22]
  reg [2:0] bht_7; // @[BHT.scala 20:22]
  reg [2:0] bht_8; // @[BHT.scala 20:22]
  reg [2:0] bht_9; // @[BHT.scala 20:22]
  reg [2:0] bht_10; // @[BHT.scala 20:22]
  reg [2:0] bht_11; // @[BHT.scala 20:22]
  reg [2:0] bht_12; // @[BHT.scala 20:22]
  reg [2:0] bht_13; // @[BHT.scala 20:22]
  reg [2:0] bht_14; // @[BHT.scala 20:22]
  reg [2:0] bht_15; // @[BHT.scala 20:22]
  reg [2:0] bht_16; // @[BHT.scala 20:22]
  reg [2:0] bht_17; // @[BHT.scala 20:22]
  reg [2:0] bht_18; // @[BHT.scala 20:22]
  reg [2:0] bht_19; // @[BHT.scala 20:22]
  reg [2:0] bht_20; // @[BHT.scala 20:22]
  reg [2:0] bht_21; // @[BHT.scala 20:22]
  reg [2:0] bht_22; // @[BHT.scala 20:22]
  reg [2:0] bht_23; // @[BHT.scala 20:22]
  reg [2:0] bht_24; // @[BHT.scala 20:22]
  reg [2:0] bht_25; // @[BHT.scala 20:22]
  reg [2:0] bht_26; // @[BHT.scala 20:22]
  reg [2:0] bht_27; // @[BHT.scala 20:22]
  reg [2:0] bht_28; // @[BHT.scala 20:22]
  reg [2:0] bht_29; // @[BHT.scala 20:22]
  reg [2:0] bht_30; // @[BHT.scala 20:22]
  reg [2:0] bht_31; // @[BHT.scala 20:22]
  reg [2:0] bht_32; // @[BHT.scala 20:22]
  reg [2:0] bht_33; // @[BHT.scala 20:22]
  reg [2:0] bht_34; // @[BHT.scala 20:22]
  reg [2:0] bht_35; // @[BHT.scala 20:22]
  reg [2:0] bht_36; // @[BHT.scala 20:22]
  reg [2:0] bht_37; // @[BHT.scala 20:22]
  reg [2:0] bht_38; // @[BHT.scala 20:22]
  reg [2:0] bht_39; // @[BHT.scala 20:22]
  reg [2:0] bht_40; // @[BHT.scala 20:22]
  reg [2:0] bht_41; // @[BHT.scala 20:22]
  reg [2:0] bht_42; // @[BHT.scala 20:22]
  reg [2:0] bht_43; // @[BHT.scala 20:22]
  reg [2:0] bht_44; // @[BHT.scala 20:22]
  reg [2:0] bht_45; // @[BHT.scala 20:22]
  reg [2:0] bht_46; // @[BHT.scala 20:22]
  reg [2:0] bht_47; // @[BHT.scala 20:22]
  reg [2:0] bht_48; // @[BHT.scala 20:22]
  reg [2:0] bht_49; // @[BHT.scala 20:22]
  reg [2:0] bht_50; // @[BHT.scala 20:22]
  reg [2:0] bht_51; // @[BHT.scala 20:22]
  reg [2:0] bht_52; // @[BHT.scala 20:22]
  reg [2:0] bht_53; // @[BHT.scala 20:22]
  reg [2:0] bht_54; // @[BHT.scala 20:22]
  reg [2:0] bht_55; // @[BHT.scala 20:22]
  reg [2:0] bht_56; // @[BHT.scala 20:22]
  reg [2:0] bht_57; // @[BHT.scala 20:22]
  reg [2:0] bht_58; // @[BHT.scala 20:22]
  reg [2:0] bht_59; // @[BHT.scala 20:22]
  reg [2:0] bht_60; // @[BHT.scala 20:22]
  reg [2:0] bht_61; // @[BHT.scala 20:22]
  reg [2:0] bht_62; // @[BHT.scala 20:22]
  reg [2:0] bht_63; // @[BHT.scala 20:22]
  reg [2:0] bht_64; // @[BHT.scala 20:22]
  reg [2:0] bht_65; // @[BHT.scala 20:22]
  reg [2:0] bht_66; // @[BHT.scala 20:22]
  reg [2:0] bht_67; // @[BHT.scala 20:22]
  reg [2:0] bht_68; // @[BHT.scala 20:22]
  reg [2:0] bht_69; // @[BHT.scala 20:22]
  reg [2:0] bht_70; // @[BHT.scala 20:22]
  reg [2:0] bht_71; // @[BHT.scala 20:22]
  reg [2:0] bht_72; // @[BHT.scala 20:22]
  reg [2:0] bht_73; // @[BHT.scala 20:22]
  reg [2:0] bht_74; // @[BHT.scala 20:22]
  reg [2:0] bht_75; // @[BHT.scala 20:22]
  reg [2:0] bht_76; // @[BHT.scala 20:22]
  reg [2:0] bht_77; // @[BHT.scala 20:22]
  reg [2:0] bht_78; // @[BHT.scala 20:22]
  reg [2:0] bht_79; // @[BHT.scala 20:22]
  reg [2:0] bht_80; // @[BHT.scala 20:22]
  reg [2:0] bht_81; // @[BHT.scala 20:22]
  reg [2:0] bht_82; // @[BHT.scala 20:22]
  reg [2:0] bht_83; // @[BHT.scala 20:22]
  reg [2:0] bht_84; // @[BHT.scala 20:22]
  reg [2:0] bht_85; // @[BHT.scala 20:22]
  reg [2:0] bht_86; // @[BHT.scala 20:22]
  reg [2:0] bht_87; // @[BHT.scala 20:22]
  reg [2:0] bht_88; // @[BHT.scala 20:22]
  reg [2:0] bht_89; // @[BHT.scala 20:22]
  reg [2:0] bht_90; // @[BHT.scala 20:22]
  reg [2:0] bht_91; // @[BHT.scala 20:22]
  reg [2:0] bht_92; // @[BHT.scala 20:22]
  reg [2:0] bht_93; // @[BHT.scala 20:22]
  reg [2:0] bht_94; // @[BHT.scala 20:22]
  reg [2:0] bht_95; // @[BHT.scala 20:22]
  reg [2:0] bht_96; // @[BHT.scala 20:22]
  reg [2:0] bht_97; // @[BHT.scala 20:22]
  reg [2:0] bht_98; // @[BHT.scala 20:22]
  reg [2:0] bht_99; // @[BHT.scala 20:22]
  reg [2:0] bht_100; // @[BHT.scala 20:22]
  reg [2:0] bht_101; // @[BHT.scala 20:22]
  reg [2:0] bht_102; // @[BHT.scala 20:22]
  reg [2:0] bht_103; // @[BHT.scala 20:22]
  reg [2:0] bht_104; // @[BHT.scala 20:22]
  reg [2:0] bht_105; // @[BHT.scala 20:22]
  reg [2:0] bht_106; // @[BHT.scala 20:22]
  reg [2:0] bht_107; // @[BHT.scala 20:22]
  reg [2:0] bht_108; // @[BHT.scala 20:22]
  reg [2:0] bht_109; // @[BHT.scala 20:22]
  reg [2:0] bht_110; // @[BHT.scala 20:22]
  reg [2:0] bht_111; // @[BHT.scala 20:22]
  reg [2:0] bht_112; // @[BHT.scala 20:22]
  reg [2:0] bht_113; // @[BHT.scala 20:22]
  reg [2:0] bht_114; // @[BHT.scala 20:22]
  reg [2:0] bht_115; // @[BHT.scala 20:22]
  reg [2:0] bht_116; // @[BHT.scala 20:22]
  reg [2:0] bht_117; // @[BHT.scala 20:22]
  reg [2:0] bht_118; // @[BHT.scala 20:22]
  reg [2:0] bht_119; // @[BHT.scala 20:22]
  reg [2:0] bht_120; // @[BHT.scala 20:22]
  reg [2:0] bht_121; // @[BHT.scala 20:22]
  reg [2:0] bht_122; // @[BHT.scala 20:22]
  reg [2:0] bht_123; // @[BHT.scala 20:22]
  reg [2:0] bht_124; // @[BHT.scala 20:22]
  reg [2:0] bht_125; // @[BHT.scala 20:22]
  reg [2:0] bht_126; // @[BHT.scala 20:22]
  reg [2:0] bht_127; // @[BHT.scala 20:22]
  wire [2:0] _GEN_1 = 7'h1 == io_ar_addr ? bht_1 : bht_0; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_2 = 7'h2 == io_ar_addr ? bht_2 : _GEN_1; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_3 = 7'h3 == io_ar_addr ? bht_3 : _GEN_2; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_4 = 7'h4 == io_ar_addr ? bht_4 : _GEN_3; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_5 = 7'h5 == io_ar_addr ? bht_5 : _GEN_4; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_6 = 7'h6 == io_ar_addr ? bht_6 : _GEN_5; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_7 = 7'h7 == io_ar_addr ? bht_7 : _GEN_6; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_8 = 7'h8 == io_ar_addr ? bht_8 : _GEN_7; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_9 = 7'h9 == io_ar_addr ? bht_9 : _GEN_8; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_10 = 7'ha == io_ar_addr ? bht_10 : _GEN_9; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_11 = 7'hb == io_ar_addr ? bht_11 : _GEN_10; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_12 = 7'hc == io_ar_addr ? bht_12 : _GEN_11; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_13 = 7'hd == io_ar_addr ? bht_13 : _GEN_12; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_14 = 7'he == io_ar_addr ? bht_14 : _GEN_13; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_15 = 7'hf == io_ar_addr ? bht_15 : _GEN_14; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_16 = 7'h10 == io_ar_addr ? bht_16 : _GEN_15; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_17 = 7'h11 == io_ar_addr ? bht_17 : _GEN_16; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_18 = 7'h12 == io_ar_addr ? bht_18 : _GEN_17; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_19 = 7'h13 == io_ar_addr ? bht_19 : _GEN_18; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_20 = 7'h14 == io_ar_addr ? bht_20 : _GEN_19; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_21 = 7'h15 == io_ar_addr ? bht_21 : _GEN_20; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_22 = 7'h16 == io_ar_addr ? bht_22 : _GEN_21; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_23 = 7'h17 == io_ar_addr ? bht_23 : _GEN_22; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_24 = 7'h18 == io_ar_addr ? bht_24 : _GEN_23; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_25 = 7'h19 == io_ar_addr ? bht_25 : _GEN_24; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_26 = 7'h1a == io_ar_addr ? bht_26 : _GEN_25; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_27 = 7'h1b == io_ar_addr ? bht_27 : _GEN_26; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_28 = 7'h1c == io_ar_addr ? bht_28 : _GEN_27; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_29 = 7'h1d == io_ar_addr ? bht_29 : _GEN_28; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_30 = 7'h1e == io_ar_addr ? bht_30 : _GEN_29; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_31 = 7'h1f == io_ar_addr ? bht_31 : _GEN_30; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_32 = 7'h20 == io_ar_addr ? bht_32 : _GEN_31; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_33 = 7'h21 == io_ar_addr ? bht_33 : _GEN_32; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_34 = 7'h22 == io_ar_addr ? bht_34 : _GEN_33; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_35 = 7'h23 == io_ar_addr ? bht_35 : _GEN_34; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_36 = 7'h24 == io_ar_addr ? bht_36 : _GEN_35; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_37 = 7'h25 == io_ar_addr ? bht_37 : _GEN_36; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_38 = 7'h26 == io_ar_addr ? bht_38 : _GEN_37; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_39 = 7'h27 == io_ar_addr ? bht_39 : _GEN_38; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_40 = 7'h28 == io_ar_addr ? bht_40 : _GEN_39; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_41 = 7'h29 == io_ar_addr ? bht_41 : _GEN_40; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_42 = 7'h2a == io_ar_addr ? bht_42 : _GEN_41; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_43 = 7'h2b == io_ar_addr ? bht_43 : _GEN_42; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_44 = 7'h2c == io_ar_addr ? bht_44 : _GEN_43; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_45 = 7'h2d == io_ar_addr ? bht_45 : _GEN_44; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_46 = 7'h2e == io_ar_addr ? bht_46 : _GEN_45; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_47 = 7'h2f == io_ar_addr ? bht_47 : _GEN_46; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_48 = 7'h30 == io_ar_addr ? bht_48 : _GEN_47; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_49 = 7'h31 == io_ar_addr ? bht_49 : _GEN_48; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_50 = 7'h32 == io_ar_addr ? bht_50 : _GEN_49; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_51 = 7'h33 == io_ar_addr ? bht_51 : _GEN_50; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_52 = 7'h34 == io_ar_addr ? bht_52 : _GEN_51; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_53 = 7'h35 == io_ar_addr ? bht_53 : _GEN_52; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_54 = 7'h36 == io_ar_addr ? bht_54 : _GEN_53; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_55 = 7'h37 == io_ar_addr ? bht_55 : _GEN_54; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_56 = 7'h38 == io_ar_addr ? bht_56 : _GEN_55; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_57 = 7'h39 == io_ar_addr ? bht_57 : _GEN_56; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_58 = 7'h3a == io_ar_addr ? bht_58 : _GEN_57; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_59 = 7'h3b == io_ar_addr ? bht_59 : _GEN_58; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_60 = 7'h3c == io_ar_addr ? bht_60 : _GEN_59; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_61 = 7'h3d == io_ar_addr ? bht_61 : _GEN_60; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_62 = 7'h3e == io_ar_addr ? bht_62 : _GEN_61; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_63 = 7'h3f == io_ar_addr ? bht_63 : _GEN_62; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_64 = 7'h40 == io_ar_addr ? bht_64 : _GEN_63; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_65 = 7'h41 == io_ar_addr ? bht_65 : _GEN_64; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_66 = 7'h42 == io_ar_addr ? bht_66 : _GEN_65; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_67 = 7'h43 == io_ar_addr ? bht_67 : _GEN_66; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_68 = 7'h44 == io_ar_addr ? bht_68 : _GEN_67; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_69 = 7'h45 == io_ar_addr ? bht_69 : _GEN_68; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_70 = 7'h46 == io_ar_addr ? bht_70 : _GEN_69; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_71 = 7'h47 == io_ar_addr ? bht_71 : _GEN_70; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_72 = 7'h48 == io_ar_addr ? bht_72 : _GEN_71; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_73 = 7'h49 == io_ar_addr ? bht_73 : _GEN_72; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_74 = 7'h4a == io_ar_addr ? bht_74 : _GEN_73; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_75 = 7'h4b == io_ar_addr ? bht_75 : _GEN_74; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_76 = 7'h4c == io_ar_addr ? bht_76 : _GEN_75; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_77 = 7'h4d == io_ar_addr ? bht_77 : _GEN_76; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_78 = 7'h4e == io_ar_addr ? bht_78 : _GEN_77; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_79 = 7'h4f == io_ar_addr ? bht_79 : _GEN_78; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_80 = 7'h50 == io_ar_addr ? bht_80 : _GEN_79; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_81 = 7'h51 == io_ar_addr ? bht_81 : _GEN_80; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_82 = 7'h52 == io_ar_addr ? bht_82 : _GEN_81; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_83 = 7'h53 == io_ar_addr ? bht_83 : _GEN_82; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_84 = 7'h54 == io_ar_addr ? bht_84 : _GEN_83; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_85 = 7'h55 == io_ar_addr ? bht_85 : _GEN_84; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_86 = 7'h56 == io_ar_addr ? bht_86 : _GEN_85; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_87 = 7'h57 == io_ar_addr ? bht_87 : _GEN_86; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_88 = 7'h58 == io_ar_addr ? bht_88 : _GEN_87; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_89 = 7'h59 == io_ar_addr ? bht_89 : _GEN_88; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_90 = 7'h5a == io_ar_addr ? bht_90 : _GEN_89; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_91 = 7'h5b == io_ar_addr ? bht_91 : _GEN_90; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_92 = 7'h5c == io_ar_addr ? bht_92 : _GEN_91; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_93 = 7'h5d == io_ar_addr ? bht_93 : _GEN_92; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_94 = 7'h5e == io_ar_addr ? bht_94 : _GEN_93; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_95 = 7'h5f == io_ar_addr ? bht_95 : _GEN_94; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_96 = 7'h60 == io_ar_addr ? bht_96 : _GEN_95; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_97 = 7'h61 == io_ar_addr ? bht_97 : _GEN_96; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_98 = 7'h62 == io_ar_addr ? bht_98 : _GEN_97; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_99 = 7'h63 == io_ar_addr ? bht_99 : _GEN_98; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_100 = 7'h64 == io_ar_addr ? bht_100 : _GEN_99; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_101 = 7'h65 == io_ar_addr ? bht_101 : _GEN_100; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_102 = 7'h66 == io_ar_addr ? bht_102 : _GEN_101; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_103 = 7'h67 == io_ar_addr ? bht_103 : _GEN_102; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_104 = 7'h68 == io_ar_addr ? bht_104 : _GEN_103; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_105 = 7'h69 == io_ar_addr ? bht_105 : _GEN_104; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_106 = 7'h6a == io_ar_addr ? bht_106 : _GEN_105; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_107 = 7'h6b == io_ar_addr ? bht_107 : _GEN_106; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_108 = 7'h6c == io_ar_addr ? bht_108 : _GEN_107; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_109 = 7'h6d == io_ar_addr ? bht_109 : _GEN_108; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_110 = 7'h6e == io_ar_addr ? bht_110 : _GEN_109; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_111 = 7'h6f == io_ar_addr ? bht_111 : _GEN_110; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_112 = 7'h70 == io_ar_addr ? bht_112 : _GEN_111; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_113 = 7'h71 == io_ar_addr ? bht_113 : _GEN_112; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_114 = 7'h72 == io_ar_addr ? bht_114 : _GEN_113; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_115 = 7'h73 == io_ar_addr ? bht_115 : _GEN_114; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_116 = 7'h74 == io_ar_addr ? bht_116 : _GEN_115; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_117 = 7'h75 == io_ar_addr ? bht_117 : _GEN_116; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_118 = 7'h76 == io_ar_addr ? bht_118 : _GEN_117; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_119 = 7'h77 == io_ar_addr ? bht_119 : _GEN_118; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_120 = 7'h78 == io_ar_addr ? bht_120 : _GEN_119; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_121 = 7'h79 == io_ar_addr ? bht_121 : _GEN_120; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_122 = 7'h7a == io_ar_addr ? bht_122 : _GEN_121; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_123 = 7'h7b == io_ar_addr ? bht_123 : _GEN_122; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_124 = 7'h7c == io_ar_addr ? bht_124 : _GEN_123; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_125 = 7'h7d == io_ar_addr ? bht_125 : _GEN_124; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_126 = 7'h7e == io_ar_addr ? bht_126 : _GEN_125; // @[BHT.scala 21:{12,12}]
  assign io_out = 7'h7f == io_ar_addr ? bht_127 : _GEN_126; // @[BHT.scala 21:{12,12}]
  always @(posedge clock) begin
    if (reset) begin // @[BHT.scala 20:22]
      bht_0 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h0 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_0 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_1 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_1 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_2 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_2 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_3 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_3 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_4 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_4 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_5 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_5 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_6 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_6 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_7 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_7 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_8 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h8 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_8 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_9 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h9 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_9 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_10 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'ha == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_10 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_11 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'hb == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_11 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_12 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'hc == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_12 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_13 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'hd == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_13 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_14 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'he == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_14 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_15 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'hf == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_15 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_16 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h10 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_16 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_17 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h11 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_17 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_18 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h12 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_18 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_19 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h13 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_19 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_20 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h14 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_20 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_21 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h15 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_21 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_22 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h16 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_22 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_23 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h17 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_23 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_24 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h18 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_24 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_25 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h19 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_25 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_26 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_26 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_27 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_27 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_28 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_28 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_29 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_29 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_30 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_30 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_31 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h1f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_31 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_32 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h20 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_32 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_33 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h21 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_33 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_34 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h22 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_34 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_35 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h23 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_35 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_36 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h24 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_36 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_37 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h25 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_37 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_38 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h26 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_38 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_39 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h27 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_39 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_40 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h28 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_40 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_41 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h29 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_41 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_42 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_42 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_43 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_43 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_44 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_44 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_45 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_45 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_46 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_46 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_47 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h2f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_47 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_48 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h30 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_48 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_49 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h31 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_49 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_50 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h32 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_50 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_51 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h33 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_51 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_52 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h34 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_52 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_53 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h35 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_53 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_54 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h36 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_54 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_55 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h37 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_55 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_56 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h38 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_56 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_57 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h39 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_57 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_58 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_58 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_59 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_59 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_60 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_60 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_61 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_61 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_62 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_62 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_63 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h3f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_63 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_64 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h40 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_64 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_65 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h41 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_65 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_66 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h42 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_66 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_67 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h43 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_67 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_68 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h44 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_68 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_69 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h45 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_69 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_70 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h46 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_70 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_71 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h47 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_71 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_72 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h48 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_72 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_73 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h49 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_73 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_74 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_74 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_75 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_75 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_76 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_76 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_77 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_77 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_78 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_78 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_79 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h4f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_79 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_80 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h50 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_80 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_81 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h51 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_81 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_82 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h52 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_82 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_83 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h53 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_83 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_84 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h54 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_84 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_85 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h55 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_85 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_86 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h56 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_86 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_87 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h57 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_87 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_88 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h58 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_88 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_89 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h59 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_89 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_90 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_90 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_91 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_91 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_92 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_92 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_93 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_93 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_94 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_94 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_95 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h5f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_95 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_96 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h60 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_96 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_97 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h61 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_97 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_98 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h62 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_98 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_99 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h63 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_99 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_100 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h64 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_100 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_101 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h65 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_101 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_102 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h66 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_102 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_103 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h67 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_103 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_104 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h68 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_104 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_105 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h69 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_105 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_106 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_106 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_107 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_107 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_108 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_108 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_109 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_109 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_110 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_110 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_111 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h6f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_111 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_112 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h70 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_112 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_113 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h71 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_113 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_114 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h72 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_114 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_115 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h73 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_115 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_116 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h74 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_116 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_117 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h75 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_117 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_118 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h76 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_118 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_119 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h77 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_119 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_120 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h78 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_120 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_121 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h79 == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_121 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_122 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7a == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_122 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_123 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7b == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_123 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_124 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7c == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_124 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_125 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7d == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_125 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_126 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7e == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_126 <= io_in;
    end
    if (reset) begin // @[BHT.scala 20:22]
      bht_127 <= 3'h0; // @[BHT.scala 20:22]
    end else if (io_write & 7'h7f == io_aw_addr) begin // @[BHT.scala 23:22]
      bht_127 <= io_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bht_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  bht_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  bht_3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  bht_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bht_5 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  bht_6 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  bht_7 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  bht_8 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  bht_9 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  bht_10 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  bht_11 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  bht_12 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  bht_13 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  bht_14 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  bht_15 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  bht_16 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  bht_17 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  bht_18 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  bht_19 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  bht_20 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  bht_21 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  bht_22 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  bht_23 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  bht_24 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  bht_25 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  bht_26 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  bht_27 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  bht_28 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  bht_29 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  bht_30 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  bht_31 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  bht_32 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  bht_33 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  bht_34 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  bht_35 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  bht_36 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  bht_37 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  bht_38 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  bht_39 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  bht_40 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  bht_41 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  bht_42 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  bht_43 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  bht_44 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  bht_45 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  bht_46 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  bht_47 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  bht_48 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  bht_49 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  bht_50 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  bht_51 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  bht_52 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  bht_53 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  bht_54 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  bht_55 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  bht_56 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  bht_57 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  bht_58 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  bht_59 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  bht_60 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  bht_61 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  bht_62 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  bht_63 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  bht_64 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  bht_65 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  bht_66 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  bht_67 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  bht_68 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  bht_69 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  bht_70 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  bht_71 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  bht_72 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  bht_73 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  bht_74 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  bht_75 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  bht_76 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  bht_77 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  bht_78 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  bht_79 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  bht_80 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  bht_81 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  bht_82 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  bht_83 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  bht_84 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  bht_85 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  bht_86 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  bht_87 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  bht_88 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  bht_89 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  bht_90 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  bht_91 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  bht_92 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  bht_93 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  bht_94 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  bht_95 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  bht_96 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  bht_97 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  bht_98 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  bht_99 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  bht_100 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  bht_101 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  bht_102 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  bht_103 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  bht_104 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  bht_105 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  bht_106 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  bht_107 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  bht_108 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  bht_109 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  bht_110 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  bht_111 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  bht_112 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  bht_113 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  bht_114 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  bht_115 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  bht_116 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  bht_117 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  bht_118 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  bht_119 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  bht_120 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  bht_121 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  bht_122 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  bht_123 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  bht_124 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  bht_125 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  bht_126 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  bht_127 = _RAND_127[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_BHT_banks_oneissue(
  input        clock,
  input        reset,
  input  [1:0] io_ar_bank_sel,
  input  [6:0] io_ar_addr,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out
);
  wire  BHT_clock; // @[BHT.scala 80:54]
  wire  BHT_reset; // @[BHT.scala 80:54]
  wire [6:0] BHT_io_ar_addr; // @[BHT.scala 80:54]
  wire [6:0] BHT_io_aw_addr; // @[BHT.scala 80:54]
  wire  BHT_io_write; // @[BHT.scala 80:54]
  wire [2:0] BHT_io_in; // @[BHT.scala 80:54]
  wire [2:0] BHT_io_out; // @[BHT.scala 80:54]
  wire  BHT_1_clock; // @[BHT.scala 80:54]
  wire  BHT_1_reset; // @[BHT.scala 80:54]
  wire [6:0] BHT_1_io_ar_addr; // @[BHT.scala 80:54]
  wire [6:0] BHT_1_io_aw_addr; // @[BHT.scala 80:54]
  wire  BHT_1_io_write; // @[BHT.scala 80:54]
  wire [2:0] BHT_1_io_in; // @[BHT.scala 80:54]
  wire [2:0] BHT_1_io_out; // @[BHT.scala 80:54]
  wire  BHT_2_clock; // @[BHT.scala 80:54]
  wire  BHT_2_reset; // @[BHT.scala 80:54]
  wire [6:0] BHT_2_io_ar_addr; // @[BHT.scala 80:54]
  wire [6:0] BHT_2_io_aw_addr; // @[BHT.scala 80:54]
  wire  BHT_2_io_write; // @[BHT.scala 80:54]
  wire [2:0] BHT_2_io_in; // @[BHT.scala 80:54]
  wire [2:0] BHT_2_io_out; // @[BHT.scala 80:54]
  wire  BHT_3_clock; // @[BHT.scala 80:54]
  wire  BHT_3_reset; // @[BHT.scala 80:54]
  wire [6:0] BHT_3_io_ar_addr; // @[BHT.scala 80:54]
  wire [6:0] BHT_3_io_aw_addr; // @[BHT.scala 80:54]
  wire  BHT_3_io_write; // @[BHT.scala 80:54]
  wire [2:0] BHT_3_io_in; // @[BHT.scala 80:54]
  wire [2:0] BHT_3_io_out; // @[BHT.scala 80:54]
  wire [2:0] bht_banks_0_out = BHT_io_out; // @[BHT.scala 80:{28,28}]
  wire [2:0] bht_banks_1_out = BHT_1_io_out; // @[BHT.scala 80:{28,28}]
  wire [2:0] _GEN_1 = 2'h1 == io_ar_bank_sel ? bht_banks_1_out : bht_banks_0_out; // @[BHT.scala 87:{12,12}]
  wire [2:0] bht_banks_2_out = BHT_2_io_out; // @[BHT.scala 80:{28,28}]
  wire [2:0] _GEN_2 = 2'h2 == io_ar_bank_sel ? bht_banks_2_out : _GEN_1; // @[BHT.scala 87:{12,12}]
  wire [2:0] bht_banks_3_out = BHT_3_io_out; // @[BHT.scala 80:{28,28}]
  ysyx_22040886_BHT BHT ( // @[BHT.scala 80:54]
    .clock(BHT_clock),
    .reset(BHT_reset),
    .io_ar_addr(BHT_io_ar_addr),
    .io_aw_addr(BHT_io_aw_addr),
    .io_write(BHT_io_write),
    .io_in(BHT_io_in),
    .io_out(BHT_io_out)
  );
  ysyx_22040886_BHT BHT_1 ( // @[BHT.scala 80:54]
    .clock(BHT_1_clock),
    .reset(BHT_1_reset),
    .io_ar_addr(BHT_1_io_ar_addr),
    .io_aw_addr(BHT_1_io_aw_addr),
    .io_write(BHT_1_io_write),
    .io_in(BHT_1_io_in),
    .io_out(BHT_1_io_out)
  );
  ysyx_22040886_BHT BHT_2 ( // @[BHT.scala 80:54]
    .clock(BHT_2_clock),
    .reset(BHT_2_reset),
    .io_ar_addr(BHT_2_io_ar_addr),
    .io_aw_addr(BHT_2_io_aw_addr),
    .io_write(BHT_2_io_write),
    .io_in(BHT_2_io_in),
    .io_out(BHT_2_io_out)
  );
  ysyx_22040886_BHT BHT_3 ( // @[BHT.scala 80:54]
    .clock(BHT_3_clock),
    .reset(BHT_3_reset),
    .io_ar_addr(BHT_3_io_ar_addr),
    .io_aw_addr(BHT_3_io_aw_addr),
    .io_write(BHT_3_io_write),
    .io_in(BHT_3_io_in),
    .io_out(BHT_3_io_out)
  );
  assign io_out = 2'h3 == io_ar_bank_sel ? bht_banks_3_out : _GEN_2; // @[BHT.scala 87:{12,12}]
  assign BHT_clock = clock;
  assign BHT_reset = reset;
  assign BHT_io_ar_addr = io_ar_addr; // @[BHT.scala 80:28 84:30]
  assign BHT_io_aw_addr = io_aw_addr; // @[BHT.scala 80:28 85:30]
  assign BHT_io_write = io_ar_bank_sel == 2'h0 & io_write; // @[BHT.scala 82:59]
  assign BHT_io_in = io_in; // @[BHT.scala 80:28 83:25]
  assign BHT_1_clock = clock;
  assign BHT_1_reset = reset;
  assign BHT_1_io_ar_addr = io_ar_addr; // @[BHT.scala 80:28 84:30]
  assign BHT_1_io_aw_addr = io_aw_addr; // @[BHT.scala 80:28 85:30]
  assign BHT_1_io_write = io_ar_bank_sel == 2'h1 & io_write; // @[BHT.scala 82:59]
  assign BHT_1_io_in = io_in; // @[BHT.scala 80:28 83:25]
  assign BHT_2_clock = clock;
  assign BHT_2_reset = reset;
  assign BHT_2_io_ar_addr = io_ar_addr; // @[BHT.scala 80:28 84:30]
  assign BHT_2_io_aw_addr = io_aw_addr; // @[BHT.scala 80:28 85:30]
  assign BHT_2_io_write = io_ar_bank_sel == 2'h2 & io_write; // @[BHT.scala 82:59]
  assign BHT_2_io_in = io_in; // @[BHT.scala 80:28 83:25]
  assign BHT_3_clock = clock;
  assign BHT_3_reset = reset;
  assign BHT_3_io_ar_addr = io_ar_addr; // @[BHT.scala 80:28 84:30]
  assign BHT_3_io_aw_addr = io_aw_addr; // @[BHT.scala 80:28 85:30]
  assign BHT_3_io_write = io_ar_bank_sel == 2'h3 & io_write; // @[BHT.scala 82:59]
  assign BHT_3_io_in = io_in; // @[BHT.scala 80:28 83:25]
endmodule
module ysyx_22040886_Look_up_table_read_first_(
  input        clock,
  input        reset,
  input  [5:0] io_ar_addr,
  input  [5:0] io_aw_addr,
  input        io_write,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_15; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_16; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_17; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_18; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_19; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_20; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_21; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_22; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_23; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_24; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_25; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_26; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_27; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_28; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_29; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_30; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_31; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_32; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_33; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_34; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_35; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_36; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_37; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_38; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_39; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_40; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_41; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_42; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_43; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_44; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_45; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_46; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_47; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_48; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_49; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_50; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_51; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_52; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_53; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_54; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_55; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_56; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_57; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_58; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_59; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_60; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_61; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_62; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_63; // @[ports_lookup_table.scala 81:22]
  wire [7:0] _GEN_1 = 6'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_2 = 6'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_3 = 6'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_4 = 6'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_5 = 6'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_6 = 6'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_7 = 6'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_8 = 6'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_9 = 6'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_10 = 6'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_11 = 6'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_12 = 6'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_13 = 6'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_14 = 6'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_15 = 6'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_16 = 6'h10 == io_ar_addr ? btb_16 : _GEN_15; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_17 = 6'h11 == io_ar_addr ? btb_17 : _GEN_16; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_18 = 6'h12 == io_ar_addr ? btb_18 : _GEN_17; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_19 = 6'h13 == io_ar_addr ? btb_19 : _GEN_18; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_20 = 6'h14 == io_ar_addr ? btb_20 : _GEN_19; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_21 = 6'h15 == io_ar_addr ? btb_21 : _GEN_20; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_22 = 6'h16 == io_ar_addr ? btb_22 : _GEN_21; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_23 = 6'h17 == io_ar_addr ? btb_23 : _GEN_22; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_24 = 6'h18 == io_ar_addr ? btb_24 : _GEN_23; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_25 = 6'h19 == io_ar_addr ? btb_25 : _GEN_24; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_26 = 6'h1a == io_ar_addr ? btb_26 : _GEN_25; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_27 = 6'h1b == io_ar_addr ? btb_27 : _GEN_26; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_28 = 6'h1c == io_ar_addr ? btb_28 : _GEN_27; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_29 = 6'h1d == io_ar_addr ? btb_29 : _GEN_28; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_30 = 6'h1e == io_ar_addr ? btb_30 : _GEN_29; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_31 = 6'h1f == io_ar_addr ? btb_31 : _GEN_30; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_32 = 6'h20 == io_ar_addr ? btb_32 : _GEN_31; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_33 = 6'h21 == io_ar_addr ? btb_33 : _GEN_32; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_34 = 6'h22 == io_ar_addr ? btb_34 : _GEN_33; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_35 = 6'h23 == io_ar_addr ? btb_35 : _GEN_34; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_36 = 6'h24 == io_ar_addr ? btb_36 : _GEN_35; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_37 = 6'h25 == io_ar_addr ? btb_37 : _GEN_36; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_38 = 6'h26 == io_ar_addr ? btb_38 : _GEN_37; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_39 = 6'h27 == io_ar_addr ? btb_39 : _GEN_38; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_40 = 6'h28 == io_ar_addr ? btb_40 : _GEN_39; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_41 = 6'h29 == io_ar_addr ? btb_41 : _GEN_40; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_42 = 6'h2a == io_ar_addr ? btb_42 : _GEN_41; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_43 = 6'h2b == io_ar_addr ? btb_43 : _GEN_42; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_44 = 6'h2c == io_ar_addr ? btb_44 : _GEN_43; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_45 = 6'h2d == io_ar_addr ? btb_45 : _GEN_44; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_46 = 6'h2e == io_ar_addr ? btb_46 : _GEN_45; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_47 = 6'h2f == io_ar_addr ? btb_47 : _GEN_46; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_48 = 6'h30 == io_ar_addr ? btb_48 : _GEN_47; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_49 = 6'h31 == io_ar_addr ? btb_49 : _GEN_48; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_50 = 6'h32 == io_ar_addr ? btb_50 : _GEN_49; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_51 = 6'h33 == io_ar_addr ? btb_51 : _GEN_50; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_52 = 6'h34 == io_ar_addr ? btb_52 : _GEN_51; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_53 = 6'h35 == io_ar_addr ? btb_53 : _GEN_52; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_54 = 6'h36 == io_ar_addr ? btb_54 : _GEN_53; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_55 = 6'h37 == io_ar_addr ? btb_55 : _GEN_54; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_56 = 6'h38 == io_ar_addr ? btb_56 : _GEN_55; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_57 = 6'h39 == io_ar_addr ? btb_57 : _GEN_56; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_58 = 6'h3a == io_ar_addr ? btb_58 : _GEN_57; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_59 = 6'h3b == io_ar_addr ? btb_59 : _GEN_58; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_60 = 6'h3c == io_ar_addr ? btb_60 : _GEN_59; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_61 = 6'h3d == io_ar_addr ? btb_61 : _GEN_60; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_62 = 6'h3e == io_ar_addr ? btb_62 : _GEN_61; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_65 = 6'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_66 = 6'h2 == io_aw_addr ? btb_2 : _GEN_65; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_67 = 6'h3 == io_aw_addr ? btb_3 : _GEN_66; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_68 = 6'h4 == io_aw_addr ? btb_4 : _GEN_67; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_69 = 6'h5 == io_aw_addr ? btb_5 : _GEN_68; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_70 = 6'h6 == io_aw_addr ? btb_6 : _GEN_69; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_71 = 6'h7 == io_aw_addr ? btb_7 : _GEN_70; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_72 = 6'h8 == io_aw_addr ? btb_8 : _GEN_71; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_73 = 6'h9 == io_aw_addr ? btb_9 : _GEN_72; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_74 = 6'ha == io_aw_addr ? btb_10 : _GEN_73; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_75 = 6'hb == io_aw_addr ? btb_11 : _GEN_74; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_76 = 6'hc == io_aw_addr ? btb_12 : _GEN_75; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_77 = 6'hd == io_aw_addr ? btb_13 : _GEN_76; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_78 = 6'he == io_aw_addr ? btb_14 : _GEN_77; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_79 = 6'hf == io_aw_addr ? btb_15 : _GEN_78; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_80 = 6'h10 == io_aw_addr ? btb_16 : _GEN_79; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_81 = 6'h11 == io_aw_addr ? btb_17 : _GEN_80; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_82 = 6'h12 == io_aw_addr ? btb_18 : _GEN_81; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_83 = 6'h13 == io_aw_addr ? btb_19 : _GEN_82; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_84 = 6'h14 == io_aw_addr ? btb_20 : _GEN_83; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_85 = 6'h15 == io_aw_addr ? btb_21 : _GEN_84; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_86 = 6'h16 == io_aw_addr ? btb_22 : _GEN_85; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_87 = 6'h17 == io_aw_addr ? btb_23 : _GEN_86; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_88 = 6'h18 == io_aw_addr ? btb_24 : _GEN_87; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_89 = 6'h19 == io_aw_addr ? btb_25 : _GEN_88; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_90 = 6'h1a == io_aw_addr ? btb_26 : _GEN_89; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_91 = 6'h1b == io_aw_addr ? btb_27 : _GEN_90; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_92 = 6'h1c == io_aw_addr ? btb_28 : _GEN_91; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_93 = 6'h1d == io_aw_addr ? btb_29 : _GEN_92; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_94 = 6'h1e == io_aw_addr ? btb_30 : _GEN_93; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_95 = 6'h1f == io_aw_addr ? btb_31 : _GEN_94; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_96 = 6'h20 == io_aw_addr ? btb_32 : _GEN_95; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_97 = 6'h21 == io_aw_addr ? btb_33 : _GEN_96; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_98 = 6'h22 == io_aw_addr ? btb_34 : _GEN_97; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_99 = 6'h23 == io_aw_addr ? btb_35 : _GEN_98; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_100 = 6'h24 == io_aw_addr ? btb_36 : _GEN_99; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_101 = 6'h25 == io_aw_addr ? btb_37 : _GEN_100; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_102 = 6'h26 == io_aw_addr ? btb_38 : _GEN_101; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_103 = 6'h27 == io_aw_addr ? btb_39 : _GEN_102; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_104 = 6'h28 == io_aw_addr ? btb_40 : _GEN_103; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_105 = 6'h29 == io_aw_addr ? btb_41 : _GEN_104; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_106 = 6'h2a == io_aw_addr ? btb_42 : _GEN_105; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_107 = 6'h2b == io_aw_addr ? btb_43 : _GEN_106; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_108 = 6'h2c == io_aw_addr ? btb_44 : _GEN_107; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_109 = 6'h2d == io_aw_addr ? btb_45 : _GEN_108; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_110 = 6'h2e == io_aw_addr ? btb_46 : _GEN_109; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_111 = 6'h2f == io_aw_addr ? btb_47 : _GEN_110; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_112 = 6'h30 == io_aw_addr ? btb_48 : _GEN_111; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_113 = 6'h31 == io_aw_addr ? btb_49 : _GEN_112; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_114 = 6'h32 == io_aw_addr ? btb_50 : _GEN_113; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_115 = 6'h33 == io_aw_addr ? btb_51 : _GEN_114; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_116 = 6'h34 == io_aw_addr ? btb_52 : _GEN_115; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_117 = 6'h35 == io_aw_addr ? btb_53 : _GEN_116; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_118 = 6'h36 == io_aw_addr ? btb_54 : _GEN_117; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_119 = 6'h37 == io_aw_addr ? btb_55 : _GEN_118; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_120 = 6'h38 == io_aw_addr ? btb_56 : _GEN_119; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_121 = 6'h39 == io_aw_addr ? btb_57 : _GEN_120; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_122 = 6'h3a == io_aw_addr ? btb_58 : _GEN_121; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_123 = 6'h3b == io_aw_addr ? btb_59 : _GEN_122; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_124 = 6'h3c == io_aw_addr ? btb_60 : _GEN_123; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_125 = 6'h3d == io_aw_addr ? btb_61 : _GEN_124; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_126 = 6'h3e == io_aw_addr ? btb_62 : _GEN_125; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 6'h3f == io_ar_addr ? btb_63 : _GEN_62; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock) begin
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_0 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_0 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_0 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_0 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_1 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_1 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_1 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_1 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_2 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_2 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_2 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_2 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_3 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_3 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_3 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_3 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_4 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_4 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_4 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_4 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_5 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_5 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_5 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_5 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_6 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_6 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_6 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_6 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_7 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_7 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_7 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_7 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_8 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_8 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_8 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_8 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_9 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_9 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_9 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_9 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_10 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'ha == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_10 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_10 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_10 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_11 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hb == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_11 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_11 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_11 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_12 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hc == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_12 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_12 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_12 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_13 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hd == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_13 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_13 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_13 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_14 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'he == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_14 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_14 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_14 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_15 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hf == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_15 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_15 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_15 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_16 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h10 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_16 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_16 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_16 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_17 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h11 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_17 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_17 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_17 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_18 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h12 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_18 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_18 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_18 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_19 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h13 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_19 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_19 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_19 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_20 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h14 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_20 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_20 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_20 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_21 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h15 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_21 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_21 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_21 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_22 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h16 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_22 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_22 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_22 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_23 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h17 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_23 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_23 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_23 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_24 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h18 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_24 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_24 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_24 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_25 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h19 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_25 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_25 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_25 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_26 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_26 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_26 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_26 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_27 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_27 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_27 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_27 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_28 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_28 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_28 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_28 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_29 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_29 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_29 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_29 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_30 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_30 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_30 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_30 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_31 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_31 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_31 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_31 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_32 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h20 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_32 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_32 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_32 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_33 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h21 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_33 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_33 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_33 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_34 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h22 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_34 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_34 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_34 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_35 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h23 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_35 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_35 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_35 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_36 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h24 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_36 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_36 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_36 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_37 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h25 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_37 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_37 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_37 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_38 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h26 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_38 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_38 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_38 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_39 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h27 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_39 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_39 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_39 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_40 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h28 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_40 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_40 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_40 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_41 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h29 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_41 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_41 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_41 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_42 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_42 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_42 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_42 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_43 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_43 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_43 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_43 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_44 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_44 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_44 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_44 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_45 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_45 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_45 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_45 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_46 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_46 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_46 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_46 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_47 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_47 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_47 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_47 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_48 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h30 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_48 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_48 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_48 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_49 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h31 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_49 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_49 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_49 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_50 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h32 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_50 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_50 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_50 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_51 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h33 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_51 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_51 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_51 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_52 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h34 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_52 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_52 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_52 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_53 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h35 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_53 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_53 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_53 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_54 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h36 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_54 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_54 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_54 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_55 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h37 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_55 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_55 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_55 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_56 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h38 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_56 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_56 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_56 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_57 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h39 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_57 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_57 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_57 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_58 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_58 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_58 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_58 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_59 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_59 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_59 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_59 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_60 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_60 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_60 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_60 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_61 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_61 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_61 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_61 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_62 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_62 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_62 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_62 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_63 <= 8'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_63 <= io_in;
      end else if (!(6'h3f == io_aw_addr)) begin // @[ports_lookup_table.scala 83:27]
        btb_63 <= _GEN_126;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  btb_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  btb_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  btb_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  btb_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  btb_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  btb_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  btb_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  btb_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  btb_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  btb_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  btb_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  btb_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  btb_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  btb_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  btb_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  btb_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  btb_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  btb_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  btb_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  btb_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  btb_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  btb_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  btb_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  btb_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  btb_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  btb_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  btb_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  btb_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  btb_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  btb_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  btb_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  btb_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  btb_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  btb_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  btb_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  btb_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  btb_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  btb_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  btb_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  btb_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  btb_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  btb_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  btb_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  btb_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  btb_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  btb_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  btb_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  btb_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  btb_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  btb_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  btb_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  btb_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  btb_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  btb_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  btb_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  btb_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  btb_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  btb_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  btb_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  btb_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  btb_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  btb_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  btb_63 = _RAND_63[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_Look_up_table_read_first__4(
  input         clock,
  input         reset,
  input  [5:0]  io_ar_addr,
  input  [5:0]  io_aw_addr,
  input         io_write,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_15; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_16; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_17; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_18; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_19; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_20; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_21; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_22; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_23; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_24; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_25; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_26; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_27; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_28; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_29; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_30; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_31; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_32; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_33; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_34; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_35; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_36; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_37; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_38; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_39; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_40; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_41; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_42; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_43; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_44; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_45; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_46; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_47; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_48; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_49; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_50; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_51; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_52; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_53; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_54; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_55; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_56; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_57; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_58; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_59; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_60; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_61; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_62; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_63; // @[ports_lookup_table.scala 81:22]
  wire [31:0] _GEN_1 = 6'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_2 = 6'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_3 = 6'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_4 = 6'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_5 = 6'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_6 = 6'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_7 = 6'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_8 = 6'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_9 = 6'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_10 = 6'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_11 = 6'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_12 = 6'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_13 = 6'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_14 = 6'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_15 = 6'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_16 = 6'h10 == io_ar_addr ? btb_16 : _GEN_15; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_17 = 6'h11 == io_ar_addr ? btb_17 : _GEN_16; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_18 = 6'h12 == io_ar_addr ? btb_18 : _GEN_17; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_19 = 6'h13 == io_ar_addr ? btb_19 : _GEN_18; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_20 = 6'h14 == io_ar_addr ? btb_20 : _GEN_19; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_21 = 6'h15 == io_ar_addr ? btb_21 : _GEN_20; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_22 = 6'h16 == io_ar_addr ? btb_22 : _GEN_21; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_23 = 6'h17 == io_ar_addr ? btb_23 : _GEN_22; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_24 = 6'h18 == io_ar_addr ? btb_24 : _GEN_23; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_25 = 6'h19 == io_ar_addr ? btb_25 : _GEN_24; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_26 = 6'h1a == io_ar_addr ? btb_26 : _GEN_25; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_27 = 6'h1b == io_ar_addr ? btb_27 : _GEN_26; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_28 = 6'h1c == io_ar_addr ? btb_28 : _GEN_27; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_29 = 6'h1d == io_ar_addr ? btb_29 : _GEN_28; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_30 = 6'h1e == io_ar_addr ? btb_30 : _GEN_29; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_31 = 6'h1f == io_ar_addr ? btb_31 : _GEN_30; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_32 = 6'h20 == io_ar_addr ? btb_32 : _GEN_31; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_33 = 6'h21 == io_ar_addr ? btb_33 : _GEN_32; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_34 = 6'h22 == io_ar_addr ? btb_34 : _GEN_33; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_35 = 6'h23 == io_ar_addr ? btb_35 : _GEN_34; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_36 = 6'h24 == io_ar_addr ? btb_36 : _GEN_35; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_37 = 6'h25 == io_ar_addr ? btb_37 : _GEN_36; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_38 = 6'h26 == io_ar_addr ? btb_38 : _GEN_37; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_39 = 6'h27 == io_ar_addr ? btb_39 : _GEN_38; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_40 = 6'h28 == io_ar_addr ? btb_40 : _GEN_39; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_41 = 6'h29 == io_ar_addr ? btb_41 : _GEN_40; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_42 = 6'h2a == io_ar_addr ? btb_42 : _GEN_41; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_43 = 6'h2b == io_ar_addr ? btb_43 : _GEN_42; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_44 = 6'h2c == io_ar_addr ? btb_44 : _GEN_43; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_45 = 6'h2d == io_ar_addr ? btb_45 : _GEN_44; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_46 = 6'h2e == io_ar_addr ? btb_46 : _GEN_45; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_47 = 6'h2f == io_ar_addr ? btb_47 : _GEN_46; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_48 = 6'h30 == io_ar_addr ? btb_48 : _GEN_47; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_49 = 6'h31 == io_ar_addr ? btb_49 : _GEN_48; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_50 = 6'h32 == io_ar_addr ? btb_50 : _GEN_49; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_51 = 6'h33 == io_ar_addr ? btb_51 : _GEN_50; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_52 = 6'h34 == io_ar_addr ? btb_52 : _GEN_51; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_53 = 6'h35 == io_ar_addr ? btb_53 : _GEN_52; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_54 = 6'h36 == io_ar_addr ? btb_54 : _GEN_53; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_55 = 6'h37 == io_ar_addr ? btb_55 : _GEN_54; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_56 = 6'h38 == io_ar_addr ? btb_56 : _GEN_55; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_57 = 6'h39 == io_ar_addr ? btb_57 : _GEN_56; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_58 = 6'h3a == io_ar_addr ? btb_58 : _GEN_57; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_59 = 6'h3b == io_ar_addr ? btb_59 : _GEN_58; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_60 = 6'h3c == io_ar_addr ? btb_60 : _GEN_59; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_61 = 6'h3d == io_ar_addr ? btb_61 : _GEN_60; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_62 = 6'h3e == io_ar_addr ? btb_62 : _GEN_61; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_65 = 6'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_66 = 6'h2 == io_aw_addr ? btb_2 : _GEN_65; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_67 = 6'h3 == io_aw_addr ? btb_3 : _GEN_66; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_68 = 6'h4 == io_aw_addr ? btb_4 : _GEN_67; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_69 = 6'h5 == io_aw_addr ? btb_5 : _GEN_68; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_70 = 6'h6 == io_aw_addr ? btb_6 : _GEN_69; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_71 = 6'h7 == io_aw_addr ? btb_7 : _GEN_70; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_72 = 6'h8 == io_aw_addr ? btb_8 : _GEN_71; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_73 = 6'h9 == io_aw_addr ? btb_9 : _GEN_72; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_74 = 6'ha == io_aw_addr ? btb_10 : _GEN_73; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_75 = 6'hb == io_aw_addr ? btb_11 : _GEN_74; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_76 = 6'hc == io_aw_addr ? btb_12 : _GEN_75; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_77 = 6'hd == io_aw_addr ? btb_13 : _GEN_76; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_78 = 6'he == io_aw_addr ? btb_14 : _GEN_77; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_79 = 6'hf == io_aw_addr ? btb_15 : _GEN_78; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_80 = 6'h10 == io_aw_addr ? btb_16 : _GEN_79; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_81 = 6'h11 == io_aw_addr ? btb_17 : _GEN_80; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_82 = 6'h12 == io_aw_addr ? btb_18 : _GEN_81; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_83 = 6'h13 == io_aw_addr ? btb_19 : _GEN_82; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_84 = 6'h14 == io_aw_addr ? btb_20 : _GEN_83; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_85 = 6'h15 == io_aw_addr ? btb_21 : _GEN_84; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_86 = 6'h16 == io_aw_addr ? btb_22 : _GEN_85; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_87 = 6'h17 == io_aw_addr ? btb_23 : _GEN_86; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_88 = 6'h18 == io_aw_addr ? btb_24 : _GEN_87; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_89 = 6'h19 == io_aw_addr ? btb_25 : _GEN_88; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_90 = 6'h1a == io_aw_addr ? btb_26 : _GEN_89; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_91 = 6'h1b == io_aw_addr ? btb_27 : _GEN_90; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_92 = 6'h1c == io_aw_addr ? btb_28 : _GEN_91; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_93 = 6'h1d == io_aw_addr ? btb_29 : _GEN_92; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_94 = 6'h1e == io_aw_addr ? btb_30 : _GEN_93; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_95 = 6'h1f == io_aw_addr ? btb_31 : _GEN_94; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_96 = 6'h20 == io_aw_addr ? btb_32 : _GEN_95; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_97 = 6'h21 == io_aw_addr ? btb_33 : _GEN_96; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_98 = 6'h22 == io_aw_addr ? btb_34 : _GEN_97; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_99 = 6'h23 == io_aw_addr ? btb_35 : _GEN_98; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_100 = 6'h24 == io_aw_addr ? btb_36 : _GEN_99; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_101 = 6'h25 == io_aw_addr ? btb_37 : _GEN_100; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_102 = 6'h26 == io_aw_addr ? btb_38 : _GEN_101; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_103 = 6'h27 == io_aw_addr ? btb_39 : _GEN_102; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_104 = 6'h28 == io_aw_addr ? btb_40 : _GEN_103; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_105 = 6'h29 == io_aw_addr ? btb_41 : _GEN_104; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_106 = 6'h2a == io_aw_addr ? btb_42 : _GEN_105; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_107 = 6'h2b == io_aw_addr ? btb_43 : _GEN_106; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_108 = 6'h2c == io_aw_addr ? btb_44 : _GEN_107; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_109 = 6'h2d == io_aw_addr ? btb_45 : _GEN_108; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_110 = 6'h2e == io_aw_addr ? btb_46 : _GEN_109; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_111 = 6'h2f == io_aw_addr ? btb_47 : _GEN_110; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_112 = 6'h30 == io_aw_addr ? btb_48 : _GEN_111; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_113 = 6'h31 == io_aw_addr ? btb_49 : _GEN_112; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_114 = 6'h32 == io_aw_addr ? btb_50 : _GEN_113; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_115 = 6'h33 == io_aw_addr ? btb_51 : _GEN_114; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_116 = 6'h34 == io_aw_addr ? btb_52 : _GEN_115; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_117 = 6'h35 == io_aw_addr ? btb_53 : _GEN_116; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_118 = 6'h36 == io_aw_addr ? btb_54 : _GEN_117; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_119 = 6'h37 == io_aw_addr ? btb_55 : _GEN_118; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_120 = 6'h38 == io_aw_addr ? btb_56 : _GEN_119; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_121 = 6'h39 == io_aw_addr ? btb_57 : _GEN_120; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_122 = 6'h3a == io_aw_addr ? btb_58 : _GEN_121; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_123 = 6'h3b == io_aw_addr ? btb_59 : _GEN_122; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_124 = 6'h3c == io_aw_addr ? btb_60 : _GEN_123; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_125 = 6'h3d == io_aw_addr ? btb_61 : _GEN_124; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_126 = 6'h3e == io_aw_addr ? btb_62 : _GEN_125; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 6'h3f == io_ar_addr ? btb_63 : _GEN_62; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock) begin
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_0 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_0 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_0 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_0 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_1 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_1 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_1 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_1 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_2 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_2 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_2 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_2 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_3 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_3 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_3 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_3 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_4 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_4 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_4 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_4 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_5 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_5 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_5 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_5 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_6 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_6 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_6 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_6 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_7 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_7 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_7 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_7 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_8 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_8 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_8 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_8 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_9 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_9 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_9 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_9 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_10 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'ha == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_10 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_10 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_10 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_11 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hb == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_11 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_11 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_11 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_12 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hc == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_12 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_12 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_12 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_13 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hd == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_13 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_13 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_13 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_14 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'he == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_14 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_14 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_14 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_15 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'hf == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_15 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_15 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_15 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_16 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h10 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_16 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_16 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_16 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_17 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h11 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_17 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_17 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_17 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_18 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h12 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_18 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_18 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_18 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_19 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h13 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_19 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_19 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_19 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_20 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h14 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_20 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_20 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_20 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_21 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h15 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_21 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_21 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_21 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_22 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h16 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_22 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_22 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_22 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_23 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h17 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_23 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_23 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_23 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_24 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h18 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_24 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_24 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_24 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_25 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h19 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_25 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_25 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_25 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_26 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_26 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_26 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_26 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_27 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_27 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_27 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_27 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_28 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_28 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_28 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_28 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_29 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_29 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_29 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_29 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_30 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_30 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_30 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_30 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_31 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h1f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_31 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_31 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_31 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_32 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h20 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_32 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_32 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_32 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_33 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h21 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_33 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_33 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_33 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_34 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h22 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_34 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_34 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_34 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_35 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h23 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_35 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_35 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_35 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_36 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h24 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_36 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_36 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_36 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_37 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h25 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_37 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_37 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_37 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_38 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h26 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_38 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_38 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_38 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_39 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h27 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_39 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_39 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_39 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_40 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h28 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_40 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_40 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_40 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_41 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h29 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_41 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_41 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_41 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_42 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_42 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_42 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_42 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_43 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_43 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_43 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_43 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_44 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_44 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_44 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_44 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_45 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_45 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_45 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_45 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_46 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_46 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_46 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_46 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_47 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h2f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_47 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_47 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_47 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_48 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h30 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_48 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_48 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_48 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_49 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h31 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_49 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_49 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_49 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_50 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h32 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_50 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_50 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_50 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_51 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h33 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_51 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_51 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_51 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_52 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h34 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_52 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_52 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_52 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_53 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h35 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_53 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_53 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_53 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_54 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h36 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_54 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_54 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_54 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_55 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h37 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_55 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_55 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_55 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_56 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h38 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_56 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_56 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_56 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_57 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h39 == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_57 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_57 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_57 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_58 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3a == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_58 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_58 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_58 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_59 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3b == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_59 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_59 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_59 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_60 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3c == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_60 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_60 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_60 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_61 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3d == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_61 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_61 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_61 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_62 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3e == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_62 <= io_in;
      end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:27]
        btb_62 <= btb_63; // @[ports_lookup_table.scala 83:27]
      end else begin
        btb_62 <= _GEN_126;
      end
    end
    if (reset) begin // @[ports_lookup_table.scala 81:22]
      btb_63 <= 32'h0; // @[ports_lookup_table.scala 81:22]
    end else if (6'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 83:21]
      if (io_write) begin // @[ports_lookup_table.scala 83:27]
        btb_63 <= io_in;
      end else if (!(6'h3f == io_aw_addr)) begin // @[ports_lookup_table.scala 83:27]
        btb_63 <= _GEN_126;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  btb_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  btb_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  btb_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  btb_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  btb_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  btb_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  btb_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  btb_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  btb_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  btb_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  btb_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  btb_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  btb_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  btb_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  btb_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  btb_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  btb_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  btb_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  btb_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  btb_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  btb_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  btb_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  btb_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  btb_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  btb_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  btb_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  btb_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  btb_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  btb_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  btb_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  btb_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  btb_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  btb_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  btb_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  btb_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  btb_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  btb_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  btb_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  btb_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  btb_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  btb_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  btb_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  btb_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  btb_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  btb_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  btb_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  btb_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  btb_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  btb_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  btb_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  btb_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  btb_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  btb_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  btb_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  btb_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  btb_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  btb_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  btb_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  btb_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  btb_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  btb_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  btb_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  btb_63 = _RAND_63[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_BTB_banks_oneissue(
  input         clock,
  input         reset,
  input  [31:0] io_ar_addr,
  input  [31:0] io_aw_addr,
  input  [31:0] io_aw_target_addr,
  input         io_write,
  output [31:0] io_out,
  output        io_hit
);
  wire  Look_up_table_read_first__clock; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__reset; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__io_ar_addr; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__io_aw_addr; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__io_write; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__io_in; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__io_out; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__1_clock; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__1_reset; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__1_io_ar_addr; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__1_io_aw_addr; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__1_io_write; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__1_io_in; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__1_io_out; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__2_clock; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__2_reset; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__2_io_ar_addr; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__2_io_aw_addr; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__2_io_write; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__2_io_in; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__2_io_out; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__3_clock; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__3_reset; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__3_io_ar_addr; // @[BTB.scala 86:54]
  wire [5:0] Look_up_table_read_first__3_io_aw_addr; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__3_io_write; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__3_io_in; // @[BTB.scala 86:54]
  wire [7:0] Look_up_table_read_first__3_io_out; // @[BTB.scala 86:54]
  wire  Look_up_table_read_first__4_clock; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__4_reset; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__4_io_ar_addr; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__4_io_aw_addr; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__4_io_write; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__4_io_in; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__4_io_out; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__5_clock; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__5_reset; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__5_io_ar_addr; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__5_io_aw_addr; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__5_io_write; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__5_io_in; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__5_io_out; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__6_clock; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__6_reset; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__6_io_ar_addr; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__6_io_aw_addr; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__6_io_write; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__6_io_in; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__6_io_out; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__7_clock; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__7_reset; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__7_io_ar_addr; // @[BTB.scala 88:54]
  wire [5:0] Look_up_table_read_first__7_io_aw_addr; // @[BTB.scala 88:54]
  wire  Look_up_table_read_first__7_io_write; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__7_io_in; // @[BTB.scala 88:54]
  wire [31:0] Look_up_table_read_first__7_io_out; // @[BTB.scala 88:54]
  wire  _btb_banks_0_write_T_1 = io_aw_addr[3:2] == 2'h0; // @[BTB.scala 90:64]
  wire  _btb_banks_1_write_T_1 = io_aw_addr[3:2] == 2'h1; // @[BTB.scala 90:64]
  wire  _btb_banks_2_write_T_1 = io_aw_addr[3:2] == 2'h2; // @[BTB.scala 90:64]
  wire  _btb_banks_3_write_T_1 = io_aw_addr[3:2] == 2'h3; // @[BTB.scala 90:64]
  wire [31:0] btb_banks_0_out = Look_up_table_read_first__4_io_out; // @[BTB.scala 88:{28,28}]
  wire [31:0] btb_banks_1_out = Look_up_table_read_first__5_io_out; // @[BTB.scala 88:{28,28}]
  wire [31:0] _GEN_1 = 2'h1 == io_ar_addr[3:2] ? btb_banks_1_out : btb_banks_0_out; // @[BTB.scala 109:{12,12}]
  wire [31:0] btb_banks_2_out = Look_up_table_read_first__6_io_out; // @[BTB.scala 88:{28,28}]
  wire [31:0] _GEN_2 = 2'h2 == io_ar_addr[3:2] ? btb_banks_2_out : _GEN_1; // @[BTB.scala 109:{12,12}]
  wire [31:0] btb_banks_3_out = Look_up_table_read_first__7_io_out; // @[BTB.scala 88:{28,28}]
  wire [7:0] tag_banks_0_out = Look_up_table_read_first__io_out; // @[BTB.scala 86:{28,28}]
  wire [7:0] tag_banks_1_out = Look_up_table_read_first__1_io_out; // @[BTB.scala 86:{28,28}]
  wire [7:0] _GEN_5 = 2'h1 == io_ar_addr[3:2] ? tag_banks_1_out : tag_banks_0_out; // @[BTB.scala 112:{62,62}]
  wire [7:0] tag_banks_2_out = Look_up_table_read_first__2_io_out; // @[BTB.scala 86:{28,28}]
  wire [7:0] _GEN_6 = 2'h2 == io_ar_addr[3:2] ? tag_banks_2_out : _GEN_5; // @[BTB.scala 112:{62,62}]
  wire [7:0] tag_banks_3_out = Look_up_table_read_first__3_io_out; // @[BTB.scala 86:{28,28}]
  wire [7:0] _GEN_7 = 2'h3 == io_ar_addr[3:2] ? tag_banks_3_out : _GEN_6; // @[BTB.scala 112:{62,62}]
  ysyx_22040886_Look_up_table_read_first_ Look_up_table_read_first_ ( // @[BTB.scala 86:54]
    .clock(Look_up_table_read_first__clock),
    .reset(Look_up_table_read_first__reset),
    .io_ar_addr(Look_up_table_read_first__io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__io_aw_addr),
    .io_write(Look_up_table_read_first__io_write),
    .io_in(Look_up_table_read_first__io_in),
    .io_out(Look_up_table_read_first__io_out)
  );
  ysyx_22040886_Look_up_table_read_first_ Look_up_table_read_first__1 ( // @[BTB.scala 86:54]
    .clock(Look_up_table_read_first__1_clock),
    .reset(Look_up_table_read_first__1_reset),
    .io_ar_addr(Look_up_table_read_first__1_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__1_io_aw_addr),
    .io_write(Look_up_table_read_first__1_io_write),
    .io_in(Look_up_table_read_first__1_io_in),
    .io_out(Look_up_table_read_first__1_io_out)
  );
  ysyx_22040886_Look_up_table_read_first_ Look_up_table_read_first__2 ( // @[BTB.scala 86:54]
    .clock(Look_up_table_read_first__2_clock),
    .reset(Look_up_table_read_first__2_reset),
    .io_ar_addr(Look_up_table_read_first__2_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__2_io_aw_addr),
    .io_write(Look_up_table_read_first__2_io_write),
    .io_in(Look_up_table_read_first__2_io_in),
    .io_out(Look_up_table_read_first__2_io_out)
  );
  ysyx_22040886_Look_up_table_read_first_ Look_up_table_read_first__3 ( // @[BTB.scala 86:54]
    .clock(Look_up_table_read_first__3_clock),
    .reset(Look_up_table_read_first__3_reset),
    .io_ar_addr(Look_up_table_read_first__3_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__3_io_aw_addr),
    .io_write(Look_up_table_read_first__3_io_write),
    .io_in(Look_up_table_read_first__3_io_in),
    .io_out(Look_up_table_read_first__3_io_out)
  );
  ysyx_22040886_Look_up_table_read_first__4 Look_up_table_read_first__4 ( // @[BTB.scala 88:54]
    .clock(Look_up_table_read_first__4_clock),
    .reset(Look_up_table_read_first__4_reset),
    .io_ar_addr(Look_up_table_read_first__4_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__4_io_aw_addr),
    .io_write(Look_up_table_read_first__4_io_write),
    .io_in(Look_up_table_read_first__4_io_in),
    .io_out(Look_up_table_read_first__4_io_out)
  );
  ysyx_22040886_Look_up_table_read_first__4 Look_up_table_read_first__5 ( // @[BTB.scala 88:54]
    .clock(Look_up_table_read_first__5_clock),
    .reset(Look_up_table_read_first__5_reset),
    .io_ar_addr(Look_up_table_read_first__5_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__5_io_aw_addr),
    .io_write(Look_up_table_read_first__5_io_write),
    .io_in(Look_up_table_read_first__5_io_in),
    .io_out(Look_up_table_read_first__5_io_out)
  );
  ysyx_22040886_Look_up_table_read_first__4 Look_up_table_read_first__6 ( // @[BTB.scala 88:54]
    .clock(Look_up_table_read_first__6_clock),
    .reset(Look_up_table_read_first__6_reset),
    .io_ar_addr(Look_up_table_read_first__6_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__6_io_aw_addr),
    .io_write(Look_up_table_read_first__6_io_write),
    .io_in(Look_up_table_read_first__6_io_in),
    .io_out(Look_up_table_read_first__6_io_out)
  );
  ysyx_22040886_Look_up_table_read_first__4 Look_up_table_read_first__7 ( // @[BTB.scala 88:54]
    .clock(Look_up_table_read_first__7_clock),
    .reset(Look_up_table_read_first__7_reset),
    .io_ar_addr(Look_up_table_read_first__7_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__7_io_aw_addr),
    .io_write(Look_up_table_read_first__7_io_write),
    .io_in(Look_up_table_read_first__7_io_in),
    .io_out(Look_up_table_read_first__7_io_out)
  );
  assign io_out = 2'h3 == io_ar_addr[3:2] ? btb_banks_3_out : _GEN_2; // @[BTB.scala 109:{12,12}]
  assign io_hit = _GEN_7[6:0] == io_ar_addr[16:10] & _GEN_7[7]; // @[BTB.scala 112:160]
  assign Look_up_table_read_first__clock = clock;
  assign Look_up_table_read_first__reset = reset;
  assign Look_up_table_read_first__io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 100:43]
  assign Look_up_table_read_first__io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 106:43]
  assign Look_up_table_read_first__io_write = _btb_banks_0_write_T_1 & io_write; // @[BTB.scala 98:77]
  assign Look_up_table_read_first__io_in = {1'h1,io_aw_addr[16:10]}; // @[Cat.scala 31:58]
  assign Look_up_table_read_first__1_clock = clock;
  assign Look_up_table_read_first__1_reset = reset;
  assign Look_up_table_read_first__1_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 100:43]
  assign Look_up_table_read_first__1_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 106:43]
  assign Look_up_table_read_first__1_io_write = _btb_banks_1_write_T_1 & io_write; // @[BTB.scala 98:77]
  assign Look_up_table_read_first__1_io_in = {1'h1,io_aw_addr[16:10]}; // @[Cat.scala 31:58]
  assign Look_up_table_read_first__2_clock = clock;
  assign Look_up_table_read_first__2_reset = reset;
  assign Look_up_table_read_first__2_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 100:43]
  assign Look_up_table_read_first__2_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 106:43]
  assign Look_up_table_read_first__2_io_write = _btb_banks_2_write_T_1 & io_write; // @[BTB.scala 98:77]
  assign Look_up_table_read_first__2_io_in = {1'h1,io_aw_addr[16:10]}; // @[Cat.scala 31:58]
  assign Look_up_table_read_first__3_clock = clock;
  assign Look_up_table_read_first__3_reset = reset;
  assign Look_up_table_read_first__3_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 100:43]
  assign Look_up_table_read_first__3_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 106:43]
  assign Look_up_table_read_first__3_io_write = _btb_banks_3_write_T_1 & io_write; // @[BTB.scala 98:77]
  assign Look_up_table_read_first__3_io_in = {1'h1,io_aw_addr[16:10]}; // @[Cat.scala 31:58]
  assign Look_up_table_read_first__4_clock = clock;
  assign Look_up_table_read_first__4_reset = reset;
  assign Look_up_table_read_first__4_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 92:43]
  assign Look_up_table_read_first__4_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 93:43]
  assign Look_up_table_read_first__4_io_write = io_aw_addr[3:2] == 2'h0 & io_write; // @[BTB.scala 90:77]
  assign Look_up_table_read_first__4_io_in = io_aw_target_addr; // @[BTB.scala 88:28 91:25]
  assign Look_up_table_read_first__5_clock = clock;
  assign Look_up_table_read_first__5_reset = reset;
  assign Look_up_table_read_first__5_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 92:43]
  assign Look_up_table_read_first__5_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 93:43]
  assign Look_up_table_read_first__5_io_write = io_aw_addr[3:2] == 2'h1 & io_write; // @[BTB.scala 90:77]
  assign Look_up_table_read_first__5_io_in = io_aw_target_addr; // @[BTB.scala 88:28 91:25]
  assign Look_up_table_read_first__6_clock = clock;
  assign Look_up_table_read_first__6_reset = reset;
  assign Look_up_table_read_first__6_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 92:43]
  assign Look_up_table_read_first__6_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 93:43]
  assign Look_up_table_read_first__6_io_write = io_aw_addr[3:2] == 2'h2 & io_write; // @[BTB.scala 90:77]
  assign Look_up_table_read_first__6_io_in = io_aw_target_addr; // @[BTB.scala 88:28 91:25]
  assign Look_up_table_read_first__7_clock = clock;
  assign Look_up_table_read_first__7_reset = reset;
  assign Look_up_table_read_first__7_io_ar_addr = io_ar_addr[9:4]; // @[BTB.scala 92:43]
  assign Look_up_table_read_first__7_io_aw_addr = io_aw_addr[9:4]; // @[BTB.scala 93:43]
  assign Look_up_table_read_first__7_io_write = io_aw_addr[3:2] == 2'h3 & io_write; // @[BTB.scala 90:77]
  assign Look_up_table_read_first__7_io_in = io_aw_target_addr; // @[BTB.scala 88:28 91:25]
endmodule
module ysyx_22040886_branch_prediction(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [31:0] io_write_pc,
  input  [3:0]  io_aw_pht_ways_addr,
  input  [6:0]  io_aw_pht_addr,
  input  [6:0]  io_aw_bht_addr,
  input  [31:0] io_aw_target_addr,
  input         io_btb_write,
  input         io_bht_write,
  input         io_pht_write,
  input  [6:0]  io_bht_in,
  input  [1:0]  io_pht_in,
  output [1:0]  io_out,
  output        io_pre,
  output [6:0]  io_bht,
  output        io_btb_hit,
  output [31:0] io_pre_target,
  input         io_stage2_stall,
  input         io_stage2_flush,
  output [6:0]  io_lookup_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  PHTS_banks_oneissue_clock; // @[branch_prediction.scala 42:28]
  wire  PHTS_banks_oneissue_reset; // @[branch_prediction.scala 42:28]
  wire  PHTS_banks_oneissue_io_ar_bank_sel; // @[branch_prediction.scala 42:28]
  wire [6:0] PHTS_banks_oneissue_io_ar_addr; // @[branch_prediction.scala 42:28]
  wire [1:0] PHTS_banks_oneissue_io_ar_pht_addr; // @[branch_prediction.scala 42:28]
  wire [6:0] PHTS_banks_oneissue_io_aw_addr; // @[branch_prediction.scala 42:28]
  wire [1:0] PHTS_banks_oneissue_io_aw_pht_addr; // @[branch_prediction.scala 42:28]
  wire  PHTS_banks_oneissue_io_aw_bank_sel; // @[branch_prediction.scala 42:28]
  wire  PHTS_banks_oneissue_io_write; // @[branch_prediction.scala 42:28]
  wire [1:0] PHTS_banks_oneissue_io_in; // @[branch_prediction.scala 42:28]
  wire [1:0] PHTS_banks_oneissue_io_out; // @[branch_prediction.scala 42:28]
  wire  BHT_banks_oneissue_clock; // @[branch_prediction.scala 43:28]
  wire  BHT_banks_oneissue_reset; // @[branch_prediction.scala 43:28]
  wire [1:0] BHT_banks_oneissue_io_ar_bank_sel; // @[branch_prediction.scala 43:28]
  wire [6:0] BHT_banks_oneissue_io_ar_addr; // @[branch_prediction.scala 43:28]
  wire [6:0] BHT_banks_oneissue_io_aw_addr; // @[branch_prediction.scala 43:28]
  wire  BHT_banks_oneissue_io_write; // @[branch_prediction.scala 43:28]
  wire [2:0] BHT_banks_oneissue_io_in; // @[branch_prediction.scala 43:28]
  wire [2:0] BHT_banks_oneissue_io_out; // @[branch_prediction.scala 43:28]
  wire  BTB_banks_oneissue_clock; // @[branch_prediction.scala 44:27]
  wire  BTB_banks_oneissue_reset; // @[branch_prediction.scala 44:27]
  wire [31:0] BTB_banks_oneissue_io_ar_addr; // @[branch_prediction.scala 44:27]
  wire [31:0] BTB_banks_oneissue_io_aw_addr; // @[branch_prediction.scala 44:27]
  wire [31:0] BTB_banks_oneissue_io_aw_target_addr; // @[branch_prediction.scala 44:27]
  wire  BTB_banks_oneissue_io_write; // @[branch_prediction.scala 44:27]
  wire [31:0] BTB_banks_oneissue_io_out; // @[branch_prediction.scala 44:27]
  wire  BTB_banks_oneissue_io_hit; // @[branch_prediction.scala 44:27]
  wire  pc_hash_num_array_0 = ^io_pc[7:4]; // @[macros.scala 455:45]
  wire  pc_hash_num_array_1 = ^io_pc[11:8]; // @[macros.scala 455:45]
  wire  pc_hash_num_array_2 = ^io_pc[15:12]; // @[macros.scala 455:45]
  wire  pc_hash_num_array_3 = ^io_pc[19:16]; // @[macros.scala 455:45]
  wire [3:0] pc_hash = {pc_hash_num_array_3,pc_hash_num_array_2,pc_hash_num_array_1,pc_hash_num_array_0}; // @[macros.scala 457:13]
  reg [6:0] stage_2_pht_lookup_0; // @[branch_prediction.scala 46:37]
  reg [63:0] stage_2_pc; // @[branch_prediction.scala 47:29]
  reg [3:0] stage_2_pc_hash; // @[branch_prediction.scala 48:34]
  reg  stage_2_btb_hit_0; // @[branch_prediction.scala 49:34]
  reg [31:0] stage_2_btb_target_pc; // @[branch_prediction.scala 50:40]
  wire [6:0] _GEN_0 = {{4'd0}, BHT_banks_oneissue_io_out}; // @[branch_prediction.scala 83:45]
  wire [6:0] stage_1_pht_lookup_0 = _GEN_0 ^ io_pc[16:10]; // @[branch_prediction.scala 83:45]
  reg [1:0] phts_out; // @[branch_prediction.scala 100:27]
  wire  _io_pre_T_3 = 2'h0 == phts_out ? 1'h0 : 2'h3 == phts_out; // @[Mux.scala 81:58]
  wire  _io_pre_T_5 = 2'h1 == phts_out ? 1'h0 : _io_pre_T_3; // @[Mux.scala 81:58]
  ysyx_22040886_PHTS_banks_oneissue PHTS_banks_oneissue ( // @[branch_prediction.scala 42:28]
    .clock(PHTS_banks_oneissue_clock),
    .reset(PHTS_banks_oneissue_reset),
    .io_ar_bank_sel(PHTS_banks_oneissue_io_ar_bank_sel),
    .io_ar_addr(PHTS_banks_oneissue_io_ar_addr),
    .io_ar_pht_addr(PHTS_banks_oneissue_io_ar_pht_addr),
    .io_aw_addr(PHTS_banks_oneissue_io_aw_addr),
    .io_aw_pht_addr(PHTS_banks_oneissue_io_aw_pht_addr),
    .io_aw_bank_sel(PHTS_banks_oneissue_io_aw_bank_sel),
    .io_write(PHTS_banks_oneissue_io_write),
    .io_in(PHTS_banks_oneissue_io_in),
    .io_out(PHTS_banks_oneissue_io_out)
  );
  ysyx_22040886_BHT_banks_oneissue BHT_banks_oneissue ( // @[branch_prediction.scala 43:28]
    .clock(BHT_banks_oneissue_clock),
    .reset(BHT_banks_oneissue_reset),
    .io_ar_bank_sel(BHT_banks_oneissue_io_ar_bank_sel),
    .io_ar_addr(BHT_banks_oneissue_io_ar_addr),
    .io_aw_addr(BHT_banks_oneissue_io_aw_addr),
    .io_write(BHT_banks_oneissue_io_write),
    .io_in(BHT_banks_oneissue_io_in),
    .io_out(BHT_banks_oneissue_io_out)
  );
  ysyx_22040886_BTB_banks_oneissue BTB_banks_oneissue ( // @[branch_prediction.scala 44:27]
    .clock(BTB_banks_oneissue_clock),
    .reset(BTB_banks_oneissue_reset),
    .io_ar_addr(BTB_banks_oneissue_io_ar_addr),
    .io_aw_addr(BTB_banks_oneissue_io_aw_addr),
    .io_aw_target_addr(BTB_banks_oneissue_io_aw_target_addr),
    .io_write(BTB_banks_oneissue_io_write),
    .io_out(BTB_banks_oneissue_io_out),
    .io_hit(BTB_banks_oneissue_io_hit)
  );
  assign io_out = phts_out; // @[branch_prediction.scala 101:12]
  assign io_pre = 2'h2 == phts_out | _io_pre_T_5; // @[Mux.scala 81:58]
  assign io_bht = {{4'd0}, BHT_banks_oneissue_io_out}; // @[branch_prediction.scala 102:12]
  assign io_btb_hit = stage_2_btb_hit_0; // @[branch_prediction.scala 51:16]
  assign io_pre_target = stage_2_btb_target_pc; // @[branch_prediction.scala 106:19]
  assign io_lookup_data = stage_2_pht_lookup_0; // @[branch_prediction.scala 66:20]
  assign PHTS_banks_oneissue_clock = clock;
  assign PHTS_banks_oneissue_reset = reset;
  assign PHTS_banks_oneissue_io_ar_bank_sel = stage_2_pc[2]; // @[branch_prediction.scala 77:28]
  assign PHTS_banks_oneissue_io_ar_addr = stage_2_pht_lookup_0; // @[branch_prediction.scala 80:24]
  assign PHTS_banks_oneissue_io_ar_pht_addr = stage_2_pc_hash[1:0]; // @[branch_prediction.scala 78:28]
  assign PHTS_banks_oneissue_io_aw_addr = io_aw_pht_addr; // @[branch_prediction.scala 85:24]
  assign PHTS_banks_oneissue_io_aw_pht_addr = io_aw_pht_ways_addr[1:0]; // @[branch_prediction.scala 86:28]
  assign PHTS_banks_oneissue_io_aw_bank_sel = io_write_pc[2]; // @[branch_prediction.scala 87:28]
  assign PHTS_banks_oneissue_io_write = io_pht_write; // @[branch_prediction.scala 88:22]
  assign PHTS_banks_oneissue_io_in = io_pht_in; // @[branch_prediction.scala 89:19]
  assign BHT_banks_oneissue_clock = clock;
  assign BHT_banks_oneissue_reset = reset;
  assign BHT_banks_oneissue_io_ar_bank_sel = io_pc[3:2]; // @[branch_prediction.scala 70:36]
  assign BHT_banks_oneissue_io_ar_addr = io_pc[10:4]; // @[branch_prediction.scala 72:32]
  assign BHT_banks_oneissue_io_aw_addr = io_aw_bht_addr; // @[branch_prediction.scala 75:24]
  assign BHT_banks_oneissue_io_write = io_bht_write; // @[branch_prediction.scala 71:22]
  assign BHT_banks_oneissue_io_in = io_bht_in[2:0]; // @[branch_prediction.scala 74:19]
  assign BTB_banks_oneissue_clock = clock;
  assign BTB_banks_oneissue_reset = reset;
  assign BTB_banks_oneissue_io_ar_addr = io_pc; // @[branch_prediction.scala 92:23]
  assign BTB_banks_oneissue_io_aw_addr = io_write_pc; // @[branch_prediction.scala 93:25]
  assign BTB_banks_oneissue_io_aw_target_addr = io_aw_target_addr; // @[branch_prediction.scala 94:30]
  assign BTB_banks_oneissue_io_write = io_btb_write; // @[branch_prediction.scala 95:21]
  always @(posedge clock) begin
    if (reset) begin // @[branch_prediction.scala 46:37]
      stage_2_pht_lookup_0 <= 7'h0; // @[branch_prediction.scala 46:37]
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 56:33]
      stage_2_pht_lookup_0 <= 7'h0;
    end else if (io_stage2_stall) begin // @[branch_prediction.scala 56:57]
      stage_2_pht_lookup_0 <= stage_1_pht_lookup_0;
    end
    if (reset) begin // @[branch_prediction.scala 47:29]
      stage_2_pc <= 64'h0; // @[branch_prediction.scala 47:29]
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 59:22]
      stage_2_pc <= 64'h0;
    end else if (io_stage2_stall) begin // @[branch_prediction.scala 59:46]
      stage_2_pc <= {{32'd0}, io_pc};
    end
    if (reset) begin // @[branch_prediction.scala 48:34]
      stage_2_pc_hash <= 4'h0; // @[branch_prediction.scala 48:34]
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 61:27]
      stage_2_pc_hash <= 4'h0;
    end else if (io_stage2_stall) begin // @[branch_prediction.scala 61:51]
      stage_2_pc_hash <= pc_hash;
    end
    if (reset) begin // @[branch_prediction.scala 49:34]
      stage_2_btb_hit_0 <= 1'h0; // @[branch_prediction.scala 49:34]
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 62:30]
      stage_2_btb_hit_0 <= 1'h0;
    end else if (io_stage2_stall) begin // @[branch_prediction.scala 62:54]
      stage_2_btb_hit_0 <= BTB_banks_oneissue_io_hit;
    end
    if (reset) begin // @[branch_prediction.scala 50:40]
      stage_2_btb_target_pc <= 32'h0; // @[branch_prediction.scala 50:40]
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 63:33]
      stage_2_btb_target_pc <= 32'h0;
    end else if (io_stage2_stall) begin // @[branch_prediction.scala 63:57]
      stage_2_btb_target_pc <= BTB_banks_oneissue_io_out;
    end
    phts_out <= PHTS_banks_oneissue_io_out; // @[branch_prediction.scala 100:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage_2_pht_lookup_0 = _RAND_0[6:0];
  _RAND_1 = {2{`RANDOM}};
  stage_2_pc = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  stage_2_pc_hash = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  stage_2_btb_hit_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  stage_2_btb_target_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  phts_out = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_bru_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [1:0]  io_in_pht,
  input  [6:0]  io_in_bht,
  input  [3:0]  io_in_hashcode,
  input  [63:0] io_in_target_pc,
  input  [6:0]  io_in_lookup_data,
  output [1:0]  io_out_pht,
  output [6:0]  io_out_bht,
  output [3:0]  io_out_hashcode,
  output [63:0] io_out_target_pc,
  output [6:0]  io_out_lookup_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pht_value; // @[myCPU.scala 641:45]
  reg [6:0] bht_value; // @[myCPU.scala 642:34]
  reg [3:0] hashcode_value; // @[myCPU.scala 643:39]
  reg [63:0] target_pc_value; // @[myCPU.scala 644:40]
  reg [6:0] lookup_data_value; // @[myCPU.scala 645:42]
  assign io_out_pht = pht_value; // @[myCPU.scala 655:20]
  assign io_out_bht = bht_value; // @[myCPU.scala 656:20]
  assign io_out_hashcode = hashcode_value; // @[myCPU.scala 657:25]
  assign io_out_target_pc = target_pc_value; // @[myCPU.scala 658:26]
  assign io_out_lookup_data = lookup_data_value; // @[myCPU.scala 659:28]
  always @(posedge clock) begin
    if (reset) begin // @[myCPU.scala 641:45]
      pht_value <= 2'h0; // @[myCPU.scala 641:45]
    end else if (io_flush) begin // @[myCPU.scala 647:25]
      pht_value <= 2'h0;
    end else if (io_stall) begin // @[myCPU.scala 647:42]
      pht_value <= io_in_pht;
    end
    if (reset) begin // @[myCPU.scala 642:34]
      bht_value <= 7'h0; // @[myCPU.scala 642:34]
    end else if (io_flush) begin // @[myCPU.scala 648:25]
      bht_value <= 7'h0;
    end else if (io_stall) begin // @[myCPU.scala 648:42]
      bht_value <= io_in_bht;
    end
    if (reset) begin // @[myCPU.scala 643:39]
      hashcode_value <= 4'h0; // @[myCPU.scala 643:39]
    end else if (io_flush) begin // @[myCPU.scala 649:30]
      hashcode_value <= 4'h0;
    end else if (io_stall) begin // @[myCPU.scala 649:47]
      hashcode_value <= io_in_hashcode;
    end
    if (reset) begin // @[myCPU.scala 644:40]
      target_pc_value <= 64'h0; // @[myCPU.scala 644:40]
    end else if (io_flush) begin // @[myCPU.scala 650:31]
      target_pc_value <= 64'h0;
    end else if (io_stall) begin // @[myCPU.scala 650:48]
      target_pc_value <= io_in_target_pc;
    end
    if (reset) begin // @[myCPU.scala 645:42]
      lookup_data_value <= 7'h0; // @[myCPU.scala 645:42]
    end else if (io_flush) begin // @[myCPU.scala 651:33]
      lookup_data_value <= 7'h0;
    end else if (io_stall) begin // @[myCPU.scala 651:50]
      lookup_data_value <= io_in_lookup_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pht_value = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  bht_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  hashcode_value = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  target_pc_value = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  lookup_data_value = _RAND_4[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_lys_cpu(
  input         clock,
  input         reset,
  input         ext_int_timer,
  input         ext_int_out_int,
  output        inst_cache,
  output        inst_sram_en,
  output [63:0] inst_sram_addr,
  input  [39:0] inst_sram_rdata_L,
  input  [1:0]  inst_write_en,
  output        stage2_flush,
  input         stage2_stall,
  output        stage1_valid_flush,
  output        inst_ready_to_use,
  output        inst_buffer_full,
  output        data_sram_en,
  output        data_sram_wen,
  output [1:0]  data_size,
  output [31:0] data_sram_addr,
  output [63:0] data_sram_wdata,
  output        data_cache,
  input  [63:0] data_sram_rdata,
  input         data_stage2_stall,
  output [7:0]  data_wstrb,
  output        data_fence_i_control,
  output        icache_tag_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] _alu_io_ctrl; // @[myCPU.scala 118:22]
  wire [63:0] _alu_io_in1; // @[myCPU.scala 118:22]
  wire [63:0] _alu_io_in2; // @[myCPU.scala 118:22]
  wire [63:0] _alu_io_result; // @[myCPU.scala 118:22]
  wire  _alu_io_overflow; // @[myCPU.scala 118:22]
  wire  _alu_io_data_w; // @[myCPU.scala 118:22]
  wire  _br_reset; // @[myCPU.scala 119:22]
  wire [63:0] _br_io_r1; // @[myCPU.scala 119:22]
  wire [63:0] _br_io_r2; // @[myCPU.scala 119:22]
  wire [5:0] _br_io_branch; // @[myCPU.scala 119:22]
  wire  _br_io_exe; // @[myCPU.scala 119:22]
  wire  _cfu_reset; // @[myCPU.scala 120:22]
  wire  _cfu_io_Inst_Fifo_Empty; // @[myCPU.scala 120:22]
  wire  _cfu_io_dmem_calD; // @[myCPU.scala 120:22]
  wire  _cfu_io_BranchD_Flag; // @[myCPU.scala 120:22]
  wire  _cfu_io_JRD; // @[myCPU.scala 120:22]
  wire  _cfu_io_CanBranchD; // @[myCPU.scala 120:22]
  wire  _cfu_io_DivPendingE; // @[myCPU.scala 120:22]
  wire  _cfu_io_DataPendingM; // @[myCPU.scala 120:22]
  wire  _cfu_io_InException; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_WriteRegE; // @[myCPU.scala 120:22]
  wire  _cfu_io_RegWriteE; // @[myCPU.scala 120:22]
  wire  _cfu_io_csrToRegE; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_WriteRegM; // @[myCPU.scala 120:22]
  wire  _cfu_io_MemToRegM; // @[myCPU.scala 120:22]
  wire  _cfu_io_RegWriteM; // @[myCPU.scala 120:22]
  wire  _cfu_io_csrWriteM; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_WriteRegM2; // @[myCPU.scala 120:22]
  wire  _cfu_io_MemToRegM2; // @[myCPU.scala 120:22]
  wire  _cfu_io_RegWriteM2; // @[myCPU.scala 120:22]
  wire  _cfu_io_csrWriteM2; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_WriteRegW; // @[myCPU.scala 120:22]
  wire  _cfu_io_RegWriteW; // @[myCPU.scala 120:22]
  wire [11:0] _cfu_io_ReadcsrAddrE; // @[myCPU.scala 120:22]
  wire [11:0] _cfu_io_WritecsrAddrM; // @[myCPU.scala 120:22]
  wire [11:0] _cfu_io_WritecsrAddrM2; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_R2D; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_R1D; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_R2E; // @[myCPU.scala 120:22]
  wire [4:0] _cfu_io_R1E; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallF; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallD; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallE; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallM; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallM2; // @[myCPU.scala 120:22]
  wire  _cfu_io_StallW; // @[myCPU.scala 120:22]
  wire  _cfu_io_FlushD; // @[myCPU.scala 120:22]
  wire  _cfu_io_FlushE; // @[myCPU.scala 120:22]
  wire  _cfu_io_FlushM; // @[myCPU.scala 120:22]
  wire  _cfu_io_FlushM2; // @[myCPU.scala 120:22]
  wire  _cfu_io_FlushW; // @[myCPU.scala 120:22]
  wire [1:0] _cfu_io_Forward1E; // @[myCPU.scala 120:22]
  wire [1:0] _cfu_io_Forward2E; // @[myCPU.scala 120:22]
  wire [1:0] _cfu_io_Forward1D; // @[myCPU.scala 120:22]
  wire [1:0] _cfu_io_Forward2D; // @[myCPU.scala 120:22]
  wire [1:0] _cfu_io_ForwardcsrE; // @[myCPU.scala 120:22]
  wire  _csr_clock; // @[myCPU.scala 121:22]
  wire  _csr_reset; // @[myCPU.scala 121:22]
  wire [11:0] _csr_io_csr_read_addr; // @[myCPU.scala 121:22]
  wire [11:0] _csr_io_csr_write_addr; // @[myCPU.scala 121:22]
  wire [63:0] _csr_io_csr_write_data; // @[myCPU.scala 121:22]
  wire  _csr_io_csr_write_en; // @[myCPU.scala 121:22]
  wire [63:0] _csr_io_pc; // @[myCPU.scala 121:22]
  wire [30:0] _csr_io_exception_type_i; // @[myCPU.scala 121:22]
  wire [63:0] _csr_io_return_pc; // @[myCPU.scala 121:22]
  wire  _csr_io_exception; // @[myCPU.scala 121:22]
  wire [63:0] _csr_io_csr_read_data; // @[myCPU.scala 121:22]
  wire  _csr_io_icache_tags_flush; // @[myCPU.scala 121:22]
  wire  _csr_io_int_type_timer; // @[myCPU.scala 121:22]
  wire  _csr_io_int_type_out_int; // @[myCPU.scala 121:22]
  wire [63:0] _csr_io_stageW_pc; // @[myCPU.scala 121:22]
  wire  _csr_io_Int_able; // @[myCPU.scala 121:22]
  wire  _csr_io_int_type_able_timer; // @[myCPU.scala 121:22]
  wire  _csr_io_int_type_able_out_int; // @[myCPU.scala 121:22]
  wire [31:0] _cu_io1_InstrD; // @[myCPU.scala 122:22]
  wire  _cu_io1_BadInstrD; // @[myCPU.scala 122:22]
  wire  _cu_io1_SysCallD; // @[myCPU.scala 122:22]
  wire  _cu_io1_EretD; // @[myCPU.scala 122:22]
  wire  _cu_io1_dmem_addr_cal; // @[myCPU.scala 122:22]
  wire  _cu_io_RegWriteD; // @[myCPU.scala 122:22]
  wire  _cu_io_MemToRegD; // @[myCPU.scala 122:22]
  wire  _cu_io_MemWriteD; // @[myCPU.scala 122:22]
  wire [15:0] _cu_io_ALUCtrlD; // @[myCPU.scala 122:22]
  wire  _cu_io_ALUSrcD_0; // @[myCPU.scala 122:22]
  wire  _cu_io_ALUSrcD_1; // @[myCPU.scala 122:22]
  wire [4:0] _cu_io_RegDstD; // @[myCPU.scala 122:22]
  wire  _cu_io_LinkD; // @[myCPU.scala 122:22]
  wire  _cu_io_csrWriteD; // @[myCPU.scala 122:22]
  wire  _cu_io_csrToRegD; // @[myCPU.scala 122:22]
  wire  _cu_io_LoadUnsignedD; // @[myCPU.scala 122:22]
  wire [1:0] _cu_io_MemWidthD; // @[myCPU.scala 122:22]
  wire [63:0] _cu_io_ImmD; // @[myCPU.scala 122:22]
  wire  _cu_io_data_wD; // @[myCPU.scala 122:22]
  wire [23:0] _cu_io_muldiv_control; // @[myCPU.scala 122:22]
  wire  _cu_io_muldiv_cal; // @[myCPU.scala 122:22]
  wire  _cu_io_alu_cal; // @[myCPU.scala 122:22]
  wire [2:0] _cu_io_csr_control; // @[myCPU.scala 122:22]
  wire  _cu_io_csr_Imm; // @[myCPU.scala 122:22]
  wire  _cu_io_fence_i_control; // @[myCPU.scala 122:22]
  wire  _dmem_io_data_ok; // @[myCPU.scala 123:23]
  wire [63:0] _dmem_io_rdata; // @[myCPU.scala 123:23]
  wire [2:0] _dmem_io_Physisc_Address; // @[myCPU.scala 123:23]
  wire [1:0] _dmem_io_WIDTH; // @[myCPU.scala 123:23]
  wire  _dmem_io_SIGN; // @[myCPU.scala 123:23]
  wire [63:0] _dmem_io_RD; // @[myCPU.scala 123:23]
  wire  _dmem_io_data_pending; // @[myCPU.scala 123:23]
  wire  _dmemreq_io_en; // @[myCPU.scala 124:26]
  wire  _dmemreq_io_MemWriteE; // @[myCPU.scala 124:26]
  wire  _dmemreq_io_MemToRegE; // @[myCPU.scala 124:26]
  wire [1:0] _dmemreq_io_MemWidthE; // @[myCPU.scala 124:26]
  wire [31:0] _dmemreq_io_VAddrE; // @[myCPU.scala 124:26]
  wire [63:0] _dmemreq_io_WriteDataE; // @[myCPU.scala 124:26]
  wire  _dmemreq_io_req; // @[myCPU.scala 124:26]
  wire  _dmemreq_io_wr; // @[myCPU.scala 124:26]
  wire [1:0] _dmemreq_io_size; // @[myCPU.scala 124:26]
  wire [31:0] _dmemreq_io_addr; // @[myCPU.scala 124:26]
  wire [63:0] _dmemreq_io_wdata; // @[myCPU.scala 124:26]
  wire [7:0] _dmemreq_io_wstrb; // @[myCPU.scala 124:26]
  wire  _ex2mem_clock; // @[myCPU.scala 125:26]
  wire  _ex2mem_reset; // @[myCPU.scala 125:26]
  wire  _ex2mem_io1_RegWriteE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io1_MemToRegE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io1_LoadUnsignedE; // @[myCPU.scala 125:26]
  wire [1:0] _ex2mem_io1_MemWidthE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io1_csrWriteE; // @[myCPU.scala 125:26]
  wire [11:0] _ex2mem_io1_WritecsrAddrE; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io1_PCE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io1_BranchJump_JrE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_en; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_clr; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_WriteDataE; // @[myCPU.scala 125:26]
  wire [4:0] _ex2mem_io_WriteRegE; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_PhyAddrE; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_CsrWritedataE; // @[myCPU.scala 125:26]
  wire [31:0] _ex2mem_io_ExceptionTypeE; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_RegWriteM; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_MemToRegM; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_WriteDataM; // @[myCPU.scala 125:26]
  wire [4:0] _ex2mem_io_WriteRegM; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 125:26]
  wire [1:0] _ex2mem_io_MemWidthM; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_PhyAddrM; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_csrWriteM; // @[myCPU.scala 125:26]
  wire [11:0] _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_PCM; // @[myCPU.scala 125:26]
  wire [31:0] _ex2mem_io_ExceptionTypeM_Out; // @[myCPU.scala 125:26]
  wire  _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 125:26]
  wire [63:0] _ex2mem_io_CsrWritedataM; // @[myCPU.scala 125:26]
  wire  _mem2mem2_clock; // @[myCPU.scala 126:28]
  wire  _mem2mem2_reset; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io1_RegWriteE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io1_MemToRegE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io1_LoadUnsignedE; // @[myCPU.scala 126:28]
  wire [1:0] _mem2mem2_io1_MemWidthE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io1_csrWriteE; // @[myCPU.scala 126:28]
  wire [11:0] _mem2mem2_io1_WritecsrAddrE; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io1_PCE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io1_BranchJump_JrE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_en; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_clr; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_WriteDataE; // @[myCPU.scala 126:28]
  wire [4:0] _mem2mem2_io_WriteRegE; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_PhyAddrE; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_CsrWritedataE; // @[myCPU.scala 126:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeE; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_RegWriteM; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_MemToRegM; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_WriteDataM; // @[myCPU.scala 126:28]
  wire [4:0] _mem2mem2_io_WriteRegM; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 126:28]
  wire [1:0] _mem2mem2_io_MemWidthM; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_PhyAddrM; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_csrWriteM; // @[myCPU.scala 126:28]
  wire [11:0] _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_PCM; // @[myCPU.scala 126:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeM_Out; // @[myCPU.scala 126:28]
  wire  _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 126:28]
  wire [63:0] _mem2mem2_io_CsrWritedataM; // @[myCPU.scala 126:28]
  wire  _id2ex_clock; // @[myCPU.scala 128:26]
  wire  _id2ex_reset; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_RegWriteD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_MemToRegD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_MemWriteD; // @[myCPU.scala 128:26]
  wire [15:0] _id2ex_io1_ALUCtrlD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_ALUSrcD_0; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_ALUSrcD_1; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io1_RegDstD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_LinkD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_csrWriteD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_csrToRegD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_LoadUnsignedD; // @[myCPU.scala 128:26]
  wire [1:0] _id2ex_io1_MemWidthD; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_data_wD; // @[myCPU.scala 128:26]
  wire [23:0] _id2ex_io1_muldiv_control; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_muldiv_cal; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_alu_cal; // @[myCPU.scala 128:26]
  wire [2:0] _id2ex_io1_csr_control; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_csr_Imm; // @[myCPU.scala 128:26]
  wire  _id2ex_io1_fence_i_control; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_RegWriteE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_MemToRegE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_MemWriteE; // @[myCPU.scala 128:26]
  wire [15:0] _id2ex_io2_ALUCtrlE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_ALUSrcE_0; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_ALUSrcE_1; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io2_RegDstE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_LinkE; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io2_PCPlus4E; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 128:26]
  wire [1:0] _id2ex_io2_MemWidthE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_csrWriteE; // @[myCPU.scala 128:26]
  wire [11:0] _id2ex_io2_WritecsrAddrE; // @[myCPU.scala 128:26]
  wire [11:0] _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io2_PCE; // @[myCPU.scala 128:26]
  wire  _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 128:26]
  wire  _id2ex_io_en; // @[myCPU.scala 128:26]
  wire  _id2ex_io_clr; // @[myCPU.scala 128:26]
  wire  _id2ex_io_csrToRegE_Out; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_RD1D; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_RD2D; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io_R2D; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io_R1D; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_ImmD; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_PCPlus4D; // @[myCPU.scala 128:26]
  wire [11:0] _id2ex_io_WritecsrAddrD; // @[myCPU.scala 128:26]
  wire [11:0] _id2ex_io_ReadcsrAddrD; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_PCD; // @[myCPU.scala 128:26]
  wire [31:0] _id2ex_io_ExceptionTypeD; // @[myCPU.scala 128:26]
  wire  _id2ex_io_BranchJump_JrD; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_RD1E; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_RD2E; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io_R2E; // @[myCPU.scala 128:26]
  wire [4:0] _id2ex_io_R1E; // @[myCPU.scala 128:26]
  wire [63:0] _id2ex_io_ImmE; // @[myCPU.scala 128:26]
  wire  _id2ex_io_data_wE; // @[myCPU.scala 128:26]
  wire [23:0] _id2ex_io_muldiv_control; // @[myCPU.scala 128:26]
  wire  _id2ex_io_alu_calE; // @[myCPU.scala 128:26]
  wire  _id2ex_io_muldiv_calE; // @[myCPU.scala 128:26]
  wire [31:0] _id2ex_io_ExceptionTypeE_Out; // @[myCPU.scala 128:26]
  wire [2:0] _id2ex_io_csr_controlE; // @[myCPU.scala 128:26]
  wire  _id2ex_io_csr_ImmE; // @[myCPU.scala 128:26]
  wire  _id2ex_io_fence_i_controlE; // @[myCPU.scala 128:26]
  wire  _if2id_clock; // @[myCPU.scala 129:26]
  wire  _if2id_reset; // @[myCPU.scala 129:26]
  wire  _if2id_io_en; // @[myCPU.scala 129:26]
  wire  _if2id_io_clr; // @[myCPU.scala 129:26]
  wire [31:0] _if2id_io_InstrF; // @[myCPU.scala 129:26]
  wire [63:0] _if2id_io_PCPlus4F; // @[myCPU.scala 129:26]
  wire [63:0] _if2id_io_PCF; // @[myCPU.scala 129:26]
  wire [1:0] _if2id_io_ExceptionTypeF; // @[myCPU.scala 129:26]
  wire [31:0] _if2id_io_InstrD; // @[myCPU.scala 129:26]
  wire [63:0] _if2id_io_PCPlus4D; // @[myCPU.scala 129:26]
  wire [63:0] _if2id_io_PCD; // @[myCPU.scala 129:26]
  wire [1:0] _if2id_io_ExceptionTypeD_Out; // @[myCPU.scala 129:26]
  wire  _mem22wb_clock; // @[myCPU.scala 131:27]
  wire  _mem22wb_reset; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_en; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_clr; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_RegWriteM; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_ResultM; // @[myCPU.scala 131:27]
  wire [4:0] _mem22wb_io_WriteRegM; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_csrWriteM; // @[myCPU.scala 131:27]
  wire [11:0] _mem22wb_io_WritecsrAddrM; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_CsrWritedataM; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_PCM; // @[myCPU.scala 131:27]
  wire [30:0] _mem22wb_io_ExceptionTypeM; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_BranchJump_JrM; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_ResultW; // @[myCPU.scala 131:27]
  wire [4:0] _mem22wb_io_WriteRegW; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_csrWriteW; // @[myCPU.scala 131:27]
  wire [11:0] _mem22wb_io_WritecsrAddrW; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_PCW; // @[myCPU.scala 131:27]
  wire [30:0] _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 131:27]
  wire  _mem22wb_io_BranchJump_JrW; // @[myCPU.scala 131:27]
  wire [63:0] _mem22wb_io_CsrWritedataW; // @[myCPU.scala 131:27]
  wire [31:0] _addr_cal_io_d_vaddr; // @[myCPU.scala 132:31]
  wire [31:0] _addr_cal_io_d_paddr; // @[myCPU.scala 132:31]
  wire  _addr_cal_io_d_cached; // @[myCPU.scala 132:31]
  wire  _muldiv_clock; // @[myCPU.scala 133:26]
  wire  _muldiv_reset; // @[myCPU.scala 133:26]
  wire  _muldiv_io_en; // @[myCPU.scala 133:26]
  wire [23:0] _muldiv_io_ctrl; // @[myCPU.scala 133:26]
  wire [63:0] _muldiv_io_in1; // @[myCPU.scala 133:26]
  wire [63:0] _muldiv_io_in2; // @[myCPU.scala 133:26]
  wire [63:0] _muldiv_io_data_out; // @[myCPU.scala 133:26]
  wire  _muldiv_io_pending; // @[myCPU.scala 133:26]
  wire  _regfile_clock; // @[myCPU.scala 135:26]
  wire  _regfile_reset; // @[myCPU.scala 135:26]
  wire [4:0] _regfile_io_A1; // @[myCPU.scala 135:26]
  wire [4:0] _regfile_io_A2; // @[myCPU.scala 135:26]
  wire  _regfile_io_WE3; // @[myCPU.scala 135:26]
  wire [4:0] _regfile_io_A3; // @[myCPU.scala 135:26]
  wire [63:0] _regfile_io_WD3; // @[myCPU.scala 135:26]
  wire [63:0] _regfile_io_RD1; // @[myCPU.scala 135:26]
  wire [63:0] _regfile_io_RD2; // @[myCPU.scala 135:26]
  wire  fifo_with_bundle_clock; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_reset; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_read_en; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_write_en; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_read_out_0_pc; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_read_out_0_inst; // @[myCPU.scala 157:29]
  wire [1:0] fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_read_out_0_pre_pc_target; // @[myCPU.scala 157:29]
  wire [6:0] fifo_with_bundle_io_read_out_0_pre_lookup_data; // @[myCPU.scala 157:29]
  wire [3:0] fifo_with_bundle_io_read_out_0_pre_hashcode; // @[myCPU.scala 157:29]
  wire [1:0] fifo_with_bundle_io_read_out_0_pre_pht; // @[myCPU.scala 157:29]
  wire [6:0] fifo_with_bundle_io_read_out_0_pre_bht; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_jump; // @[myCPU.scala 157:29]
  wire [5:0] fifo_with_bundle_io_read_out_0_pre_decoder_branchdata; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_jr; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_read_out_0_true_branch_state; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_write_in_0_pc; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_write_in_0_inst; // @[myCPU.scala 157:29]
  wire [31:0] fifo_with_bundle_io_write_in_0_pre_pc_target; // @[myCPU.scala 157:29]
  wire [6:0] fifo_with_bundle_io_write_in_0_pre_lookup_data; // @[myCPU.scala 157:29]
  wire [3:0] fifo_with_bundle_io_write_in_0_pre_hashcode; // @[myCPU.scala 157:29]
  wire [1:0] fifo_with_bundle_io_write_in_0_pre_pht; // @[myCPU.scala 157:29]
  wire [6:0] fifo_with_bundle_io_write_in_0_pre_bht; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_jump; // @[myCPU.scala 157:29]
  wire [5:0] fifo_with_bundle_io_write_in_0_pre_decoder_branchdata; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_jr; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_write_in_0_true_branch_state; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_full; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_empty; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_point_write_en; // @[myCPU.scala 157:29]
  wire  fifo_with_bundle_io_point_flush; // @[myCPU.scala 157:29]
  wire  stage_fec_1_pc_L_clock; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_L_reset; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_L_io_stall; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_L_io_flush; // @[myCPU.scala 423:34]
  wire [31:0] stage_fec_1_pc_L_io_in_pc_value_in; // @[myCPU.scala 423:34]
  wire [31:0] stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 423:34]
  wire  branch_prediction_clock; // @[myCPU.scala 447:21]
  wire  branch_prediction_reset; // @[myCPU.scala 447:21]
  wire [31:0] branch_prediction_io_pc; // @[myCPU.scala 447:21]
  wire [31:0] branch_prediction_io_write_pc; // @[myCPU.scala 447:21]
  wire [3:0] branch_prediction_io_aw_pht_ways_addr; // @[myCPU.scala 447:21]
  wire [6:0] branch_prediction_io_aw_pht_addr; // @[myCPU.scala 447:21]
  wire [6:0] branch_prediction_io_aw_bht_addr; // @[myCPU.scala 447:21]
  wire [31:0] branch_prediction_io_aw_target_addr; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_btb_write; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_bht_write; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_pht_write; // @[myCPU.scala 447:21]
  wire [6:0] branch_prediction_io_bht_in; // @[myCPU.scala 447:21]
  wire [1:0] branch_prediction_io_pht_in; // @[myCPU.scala 447:21]
  wire [1:0] branch_prediction_io_out; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_pre; // @[myCPU.scala 447:21]
  wire [6:0] branch_prediction_io_bht; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_btb_hit; // @[myCPU.scala 447:21]
  wire [31:0] branch_prediction_io_pre_target; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_stage2_stall; // @[myCPU.scala 447:21]
  wire  branch_prediction_io_stage2_flush; // @[myCPU.scala 447:21]
  wire [6:0] branch_prediction_io_lookup_data; // @[myCPU.scala 447:21]
  wire  stage_fec_2_pc_L_clock; // @[myCPU.scala 509:34]
  wire  stage_fec_2_pc_L_reset; // @[myCPU.scala 509:34]
  wire  stage_fec_2_pc_L_io_stall; // @[myCPU.scala 509:34]
  wire  stage_fec_2_pc_L_io_flush; // @[myCPU.scala 509:34]
  wire [31:0] stage_fec_2_pc_L_io_in_pc_value_in; // @[myCPU.scala 509:34]
  wire [31:0] stage_fec_2_pc_L_io_out_pc_value_out; // @[myCPU.scala 509:34]
  wire  id_bru_state_clock; // @[myCPU.scala 666:31]
  wire  id_bru_state_reset; // @[myCPU.scala 666:31]
  wire  id_bru_state_io_stall; // @[myCPU.scala 666:31]
  wire  id_bru_state_io_flush; // @[myCPU.scala 666:31]
  wire [1:0] id_bru_state_io_in_pht; // @[myCPU.scala 666:31]
  wire [6:0] id_bru_state_io_in_bht; // @[myCPU.scala 666:31]
  wire [3:0] id_bru_state_io_in_hashcode; // @[myCPU.scala 666:31]
  wire [63:0] id_bru_state_io_in_target_pc; // @[myCPU.scala 666:31]
  wire [6:0] id_bru_state_io_in_lookup_data; // @[myCPU.scala 666:31]
  wire [1:0] id_bru_state_io_out_pht; // @[myCPU.scala 666:31]
  wire [6:0] id_bru_state_io_out_bht; // @[myCPU.scala 666:31]
  wire [3:0] id_bru_state_io_out_hashcode; // @[myCPU.scala 666:31]
  wire [63:0] id_bru_state_io_out_target_pc; // @[myCPU.scala 666:31]
  wire [6:0] id_bru_state_io_out_lookup_data; // @[myCPU.scala 666:31]
  wire  ex_bru_state_clock; // @[myCPU.scala 670:31]
  wire  ex_bru_state_reset; // @[myCPU.scala 670:31]
  wire  ex_bru_state_io_stall; // @[myCPU.scala 670:31]
  wire  ex_bru_state_io_flush; // @[myCPU.scala 670:31]
  wire [1:0] ex_bru_state_io_in_pht; // @[myCPU.scala 670:31]
  wire [6:0] ex_bru_state_io_in_bht; // @[myCPU.scala 670:31]
  wire [3:0] ex_bru_state_io_in_hashcode; // @[myCPU.scala 670:31]
  wire [63:0] ex_bru_state_io_in_target_pc; // @[myCPU.scala 670:31]
  wire [6:0] ex_bru_state_io_in_lookup_data; // @[myCPU.scala 670:31]
  wire [1:0] ex_bru_state_io_out_pht; // @[myCPU.scala 670:31]
  wire [6:0] ex_bru_state_io_out_bht; // @[myCPU.scala 670:31]
  wire [3:0] ex_bru_state_io_out_hashcode; // @[myCPU.scala 670:31]
  wire [63:0] ex_bru_state_io_out_target_pc; // @[myCPU.scala 670:31]
  wire [6:0] ex_bru_state_io_out_lookup_data; // @[myCPU.scala 670:31]
  wire  mem_bru_state_clock; // @[myCPU.scala 674:32]
  wire  mem_bru_state_reset; // @[myCPU.scala 674:32]
  wire  mem_bru_state_io_stall; // @[myCPU.scala 674:32]
  wire  mem_bru_state_io_flush; // @[myCPU.scala 674:32]
  wire [1:0] mem_bru_state_io_in_pht; // @[myCPU.scala 674:32]
  wire [6:0] mem_bru_state_io_in_bht; // @[myCPU.scala 674:32]
  wire [3:0] mem_bru_state_io_in_hashcode; // @[myCPU.scala 674:32]
  wire [63:0] mem_bru_state_io_in_target_pc; // @[myCPU.scala 674:32]
  wire [6:0] mem_bru_state_io_in_lookup_data; // @[myCPU.scala 674:32]
  wire [1:0] mem_bru_state_io_out_pht; // @[myCPU.scala 674:32]
  wire [6:0] mem_bru_state_io_out_bht; // @[myCPU.scala 674:32]
  wire [3:0] mem_bru_state_io_out_hashcode; // @[myCPU.scala 674:32]
  wire [63:0] mem_bru_state_io_out_target_pc; // @[myCPU.scala 674:32]
  wire [6:0] mem_bru_state_io_out_lookup_data; // @[myCPU.scala 674:32]
  wire  mem2_bru_state_clock; // @[myCPU.scala 678:33]
  wire  mem2_bru_state_reset; // @[myCPU.scala 678:33]
  wire  mem2_bru_state_io_stall; // @[myCPU.scala 678:33]
  wire  mem2_bru_state_io_flush; // @[myCPU.scala 678:33]
  wire [1:0] mem2_bru_state_io_in_pht; // @[myCPU.scala 678:33]
  wire [6:0] mem2_bru_state_io_in_bht; // @[myCPU.scala 678:33]
  wire [3:0] mem2_bru_state_io_in_hashcode; // @[myCPU.scala 678:33]
  wire [63:0] mem2_bru_state_io_in_target_pc; // @[myCPU.scala 678:33]
  wire [6:0] mem2_bru_state_io_in_lookup_data; // @[myCPU.scala 678:33]
  wire [1:0] mem2_bru_state_io_out_pht; // @[myCPU.scala 678:33]
  wire [6:0] mem2_bru_state_io_out_bht; // @[myCPU.scala 678:33]
  wire [3:0] mem2_bru_state_io_out_hashcode; // @[myCPU.scala 678:33]
  wire [63:0] mem2_bru_state_io_out_target_pc; // @[myCPU.scala 678:33]
  wire [6:0] mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 678:33]
  wire  wb_bru_state_clock; // @[myCPU.scala 682:31]
  wire  wb_bru_state_reset; // @[myCPU.scala 682:31]
  wire  wb_bru_state_io_stall; // @[myCPU.scala 682:31]
  wire  wb_bru_state_io_flush; // @[myCPU.scala 682:31]
  wire [1:0] wb_bru_state_io_in_pht; // @[myCPU.scala 682:31]
  wire [6:0] wb_bru_state_io_in_bht; // @[myCPU.scala 682:31]
  wire [3:0] wb_bru_state_io_in_hashcode; // @[myCPU.scala 682:31]
  wire [63:0] wb_bru_state_io_in_target_pc; // @[myCPU.scala 682:31]
  wire [6:0] wb_bru_state_io_in_lookup_data; // @[myCPU.scala 682:31]
  wire [1:0] wb_bru_state_io_out_pht; // @[myCPU.scala 682:31]
  wire [6:0] wb_bru_state_io_out_bht; // @[myCPU.scala 682:31]
  wire [3:0] wb_bru_state_io_out_hashcode; // @[myCPU.scala 682:31]
  wire [63:0] wb_bru_state_io_out_target_pc; // @[myCPU.scala 682:31]
  wire [6:0] wb_bru_state_io_out_lookup_data; // @[myCPU.scala 682:31]
  wire  stage_fec_2_inst_jump = inst_sram_rdata_L[33]; // @[myCPU.scala 177:45]
  wire  stage_fec_2_inst_branch = inst_sram_rdata_L[32]; // @[myCPU.scala 178:47]
  reg  pre_decoder_branchD_flag; // @[myCPU.scala 180:44]
  reg [5:0] pre_decoder_branchdata; // @[myCPU.scala 181:43]
  reg  pre_decoder_jump; // @[myCPU.scala 182:40]
  reg  pre_decoder_jr; // @[myCPU.scala 183:40]
  wire [12:0] _immSB_T_4 = {_if2id_io_InstrD[31],_if2id_io_InstrD[7],_if2id_io_InstrD[30:25],_if2id_io_InstrD[11:8],1'h0
    }; // @[Cat.scala 31:58]
  wire [5:0] immSB_lo_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12]
    }; // @[Cat.scala 31:58]
  wire [11:0] immSB_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [12:0] immSB_lo_hi = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [24:0] immSB_lo_1 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_lo}; // @[Cat.scala 31:58]
  wire [50:0] _immSB_T_56 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_hi,immSB_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] immSB = {_immSB_T_56,_if2id_io_InstrD[31],_if2id_io_InstrD[7],_if2id_io_InstrD[30:25],_if2id_io_InstrD[11:
    8],1'h0}; // @[Cat.scala 31:58]
  wire  _PCSrcD_T_1 = _cfu_io_StallD; // @[myCPU.scala 198:66]
  wire  _PCSrcD_T_3 = _br_io_exe; // @[myCPU.scala 198:85]
  wire [63:0] PCBranchD = immSB + _if2id_io_PCD; // @[myCPU.scala 199:27]
  wire [20:0] _immUJ_T_4 = {_if2id_io_InstrD[31],_if2id_io_InstrD[19:12],_if2id_io_InstrD[20],_if2id_io_InstrD[30:21],1'h0
    }; // @[Cat.scala 31:58]
  wire [4:0] immUJ_lo_lo_lo = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20]}; // @[Cat.scala 31:58]
  wire [9:0] immUJ_lo_lo = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    _immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20]}; // @[Cat.scala 31:58]
  wire [10:0] immUJ_lo_hi = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [20:0] immUJ_lo_1 = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo,immUJ_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] immUJ = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo,immUJ_lo_hi,immUJ_lo_1,_immUJ_T_4}; // @[Cat.scala 31:58]
  wire [5:0] PCJumpD_lo_lo_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31]}; // @[Cat.scala 31:58]
  wire [12:0] PCJumpD_lo_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] PCJumpD_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo,PCJumpD_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _PCJumpD_T_54 = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo,PCJumpD_lo_lo,PCJumpD_lo}; // @[Cat.scala 31:58]
  wire [63:0] _PCJumpD_T_56 = {_PCJumpD_T_54,_if2id_io_InstrD[31:20]}; // @[Cat.scala 31:58]
  reg [63:0] resultE2M_Reg; // @[myCPU.scala 963:32]
  reg [63:0] ResultM2_Reg; // @[myCPU.scala 1016:29]
  wire [63:0] _BranchR1D_T_2 = _cfu_io_Forward1D[1] ? ResultM2_Reg : _regfile_io_RD1; // @[myCPU.scala 751:61]
  wire [63:0] BranchR1D = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 751:20]
  wire [63:0] _PCJumpD_T_58 = BranchR1D + _PCJumpD_T_56; // @[myCPU.scala 202:58]
  wire [63:0] _PCJumpD_T_60 = immUJ + _if2id_io_PCD; // @[myCPU.scala 202:107]
  wire [63:0] PCJumpD = pre_decoder_jr ? _PCJumpD_T_58 : _PCJumpD_T_60; // @[myCPU.scala 202:24]
  reg  fence_i_controlMReg; // @[myCPU.scala 264:34]
  reg [63:0] PCW_Reg; // @[myCPU.scala 299:26]
  wire  _PCW_Reg_T = _mem22wb_io_PCW != 64'h0; // @[myCPU.scala 303:36]
  reg [63:0] pc_next_wait; // @[myCPU.scala 344:33]
  wire  ready_to_branch = fifo_with_bundle_io_point_write_en; // @[myCPU.scala 346:31 580:21]
  reg  stage_fec_2_stall_reg; // @[myCPU.scala 496:40]
  reg  stage_fec_2_valid; // @[myCPU.scala 472:36]
  wire  _stage_fec_2_branch_answer_T_8 = _csr_io_exception; // @[myCPU.scala 499:207]
  wire  _stage_fec_2_branch_answer_T_9 = ~_csr_io_exception; // @[myCPU.scala 499:188]
  wire  stage_fec_2_branch_answer = branch_prediction_io_pre & (stage_fec_2_inst_branch | stage_fec_2_inst_jump) &
    branch_prediction_io_btb_hit & stage_fec_2_stall_reg & stage_fec_2_valid & ~_csr_io_exception; // @[myCPU.scala 499:185]
  wire  _pc_next_wait_T = ready_to_branch | stage_fec_2_branch_answer; // @[myCPU.scala 347:41]
  wire [63:0] _PC_nextD_T_2 = _PCSrcD_T_3 ? PCBranchD : _if2id_io_PCPlus4D; // @[Mux.scala 101:16]
  wire [63:0] PC_nextD = pre_decoder_jump ? PCJumpD : _PC_nextD_T_2; // @[Mux.scala 101:16]
  wire [63:0] stage_fec_2_pre_target_0 = {{32'd0}, branch_prediction_io_pre_target}; // @[myCPU.scala 477:38 490:31]
  wire [63:0] stage_fec_1_pc = {{32'd0}, stage_fec_1_pc_L_io_out_pc_value_out}; // @[myCPU.scala 174:26 444:20]
  wire [63:0] _stage_fec_1_pc_next_T_1 = stage_fec_1_pc + 64'h4; // @[myCPU.scala 418:93]
  wire [63:0] stage_fec_1_pc_next = stage_fec_2_branch_answer ? stage_fec_2_pre_target_0 : _stage_fec_1_pc_next_T_1; // @[myCPU.scala 418:31]
  wire [63:0] Pc_Next_normal = fifo_with_bundle_io_point_write_en ? PC_nextD : stage_fec_1_pc_next; // @[myCPU.scala 743:26]
  reg  pc_req_wait; // @[myCPU.scala 348:30]
  wire  _T_1 = ~inst_sram_en; // @[myCPU.scala 352:10]
  wire  _GEN_0 = pc_req_wait & inst_sram_en | _stage_fec_2_branch_answer_T_8 | ready_to_branch & inst_sram_en ? 1'h0 :
    pc_req_wait; // @[myCPU.scala 354:119 355:21 357:21]
  wire  _GEN_1 = ~inst_sram_en & _pc_next_wait_T & _stage_fec_2_branch_answer_T_9 | _GEN_0; // @[myCPU.scala 352:102 353:21]
  reg [63:0] exception_Pc_reg; // @[myCPU.scala 361:35]
  reg  returnPc_req_wait; // @[myCPU.scala 364:36]
  wire  _GEN_2 = returnPc_req_wait & inst_sram_en ? 1'h0 : returnPc_req_wait; // @[myCPU.scala 369:54 370:27 372:27]
  wire  _GEN_3 = _T_1 & _stage_fec_2_branch_answer_T_8 | _GEN_2; // @[myCPU.scala 367:58 368:27]
  wire [63:0] _inst_sram_addr_T_1 = pc_req_wait ? pc_next_wait : Pc_Next_normal; // @[myCPU.scala 379:142]
  wire [63:0] _inst_sram_addr_T_2 = ready_to_branch ? Pc_Next_normal : _inst_sram_addr_T_1; // @[myCPU.scala 379:107]
  wire [63:0] _inst_sram_addr_T_3 = returnPc_req_wait ? exception_Pc_reg : _inst_sram_addr_T_2; // @[myCPU.scala 379:68]
  wire  _commit_cache_reg_T = _cfu_io_StallE; // @[myCPU.scala 401:40]
  reg  stage_fec_1_valid; // @[myCPU.scala 451:36]
  wire  _stage_fec_1_valid_T_2 = _pc_next_wait_T ? 1'h0 : stage_fec_1_valid; // @[myCPU.scala 455:55]
  wire  stage_fec_2_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 465:42]
  reg [6:0] stage_fec_2_bht_0; // @[myCPU.scala 475:35]
  reg [3:0] stage_fec_2_hascode_0; // @[myCPU.scala 479:39]
  wire  stage_fec_2_hascode_0_num_array_0 = ^branch_prediction_io_pc[7:4]; // @[macros.scala 455:45]
  wire  stage_fec_2_hascode_0_num_array_1 = ^branch_prediction_io_pc[11:8]; // @[macros.scala 455:45]
  wire  stage_fec_2_hascode_0_num_array_2 = ^branch_prediction_io_pc[15:12]; // @[macros.scala 455:45]
  wire  stage_fec_2_hascode_0_num_array_3 = ^branch_prediction_io_pc[19:16]; // @[macros.scala 455:45]
  wire [3:0] _stage_fec_2_hascode_0_T_1 = {stage_fec_2_hascode_0_num_array_3,stage_fec_2_hascode_0_num_array_2,
    stage_fec_2_hascode_0_num_array_1,stage_fec_2_hascode_0_num_array_0}; // @[macros.scala 457:13]
  wire  _stage_fec_2_data_valid_T = ~fifo_with_bundle_io_empty; // @[myCPU.scala 516:88]
  wire [31:0] inst_buffer_write_bundle_inst = inst_sram_rdata_L[31:0]; // @[myCPU.scala 531:60]
  wire [6:0] inst_buffer_write_bundle_pre_decoder_jr_opD = inst_buffer_write_bundle_inst[6:0]; // @[macros.scala 503:24]
  wire [2:0] inst_buffer_write_bundle_pre_decoder_jr_Funct3D = inst_buffer_write_bundle_inst[14:12]; // @[macros.scala 504:28]
  wire  _pre_decoder_branchD_flag_T = _cfu_io_FlushD; // @[myCPU.scala 587:52]
  wire  inst_buffer_read_out_pre_decoder_branchD_flag = fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag; // @[myCPU.scala 583:36 584:26]
  wire  inst_buffer_read_out_pre_decoder_jump = fifo_with_bundle_io_read_out_0_pre_decoder_jump; // @[myCPU.scala 583:36 584:26]
  wire [5:0] inst_buffer_read_out_pre_decoder_branchdata = fifo_with_bundle_io_read_out_0_pre_decoder_branchdata; // @[myCPU.scala 583:36 584:26]
  wire  inst_buffer_read_out_pre_decoder_jr = fifo_with_bundle_io_read_out_0_pre_decoder_jr; // @[myCPU.scala 583:36 584:26]
  wire  __if2id_io_InstrF_T = _cu_io1_BadInstrD; // @[myCPU.scala 602:52]
  wire  __if2id_io_InstrF_T_1 = _cu_io1_SysCallD; // @[myCPU.scala 602:79]
  wire  __if2id_io_InstrF_T_3 = _cu_io1_EretD; // @[myCPU.scala 603:47]
  wire [31:0] inst_buffer_read_out_inst = fifo_with_bundle_io_read_out_0_inst; // @[myCPU.scala 583:36 584:26]
  reg  id_exception; // @[myCPU.scala 606:31]
  wire [1:0] inst_buffer_read_out_exception_type = fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 583:36 584:26]
  reg  ex_exception; // @[myCPU.scala 609:31]
  wire  _ex_exception_T = _cfu_io_FlushE; // @[myCPU.scala 610:40]
  reg  mem_exception; // @[myCPU.scala 612:32]
  wire  _mem_exception_T = _cfu_io_FlushM; // @[myCPU.scala 613:41]
  wire  _mem_exception_T_1 = _cfu_io_StallM; // @[myCPU.scala 613:71]
  reg  mem2_exception; // @[myCPU.scala 615:33]
  wire  _mem2_exception_T = _cfu_io_FlushM2; // @[myCPU.scala 616:43]
  wire  _mem2_exception_T_1 = _cfu_io_StallM2; // @[myCPU.scala 616:74]
  reg  wb_exception; // @[myCPU.scala 618:31]
  wire  _wb_exception_T = _cfu_io_FlushW; // @[myCPU.scala 619:40]
  wire  _wb_exception_T_1 = _cfu_io_StallW; // @[myCPU.scala 619:70]
  reg  id_true_branch_state; // @[myCPU.scala 663:39]
  wire  inst_buffer_read_out_true_branch_state = fifo_with_bundle_io_read_out_0_true_branch_state; // @[myCPU.scala 583:36 584:26]
  reg  inst_tlb_exceptionE; // @[myCPU.scala 693:38]
  wire  target_neq_branchD = id_bru_state_io_out_target_pc != PCBranchD; // @[myCPU.scala 704:62]
  wire  target_neq_jumpD = id_bru_state_io_out_target_pc != PCJumpD; // @[myCPU.scala 705:62]
  wire  target_addr_error = pre_decoder_jump & target_neq_jumpD | _PCSrcD_T_3 & target_neq_branchD; // @[myCPU.scala 707:75]
  wire  _T_28 = pre_decoder_jump | _PCSrcD_T_3; // @[myCPU.scala 710:117]
  wire  _T_34 = ex_exception | mem_exception | mem2_exception | wb_exception; // @[myCPU.scala 710:241]
  wire [63:0] _Pc_targetD_T_2 = pre_decoder_jump ? PCJumpD : 64'h0; // @[Mux.scala 101:16]
  reg  true_branch_stateE; // @[myCPU.scala 721:37]
  wire [1:0] _pht_tobeE_T_1 = true_branch_stateE ? 2'h3 : 2'h2; // @[macros.scala 476:30]
  wire [1:0] _pht_tobeE_T_2 = true_branch_stateE ? 2'h2 : 2'h0; // @[macros.scala 477:32]
  wire [1:0] _pht_tobeE_T_3 = true_branch_stateE ? 2'h3 : 2'h1; // @[macros.scala 478:30]
  wire [1:0] _pht_tobeE_T_5 = 2'h3 == ex_bru_state_io_out_pht ? _pht_tobeE_T_1 : {{1'd0}, true_branch_stateE}; // @[Mux.scala 81:58]
  wire [1:0] _pht_tobeE_T_7 = 2'h1 == ex_bru_state_io_out_pht ? _pht_tobeE_T_2 : _pht_tobeE_T_5; // @[Mux.scala 81:58]
  wire [63:0] _BranchR2D_T_2 = _cfu_io_Forward2D[1] ? ResultM2_Reg : _regfile_io_RD2; // @[myCPU.scala 753:61]
  wire  _ExceptionTypeD_Out_T_1 = _if2id_io_PCD[1:0] != 2'h0; // @[myCPU.scala 755:29]
  wire [20:0] _ExceptionTypeD_Out_T_4 = _ExceptionTypeD_Out_T_1 ? 21'h100000 : 21'h0; // @[Mux.scala 27:73]
  wire [3:0] _ExceptionTypeD_Out_T_5 = _if2id_io_ExceptionTypeD_Out[0] ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _ExceptionTypeD_Out_T_6 = _if2id_io_ExceptionTypeD_Out[1] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [24:0] _ExceptionTypeD_Out_T_7 = _cu_io_fence_i_control ? 25'h1000000 : 25'h0; // @[Mux.scala 27:73]
  wire [20:0] _GEN_12 = {{17'd0}, _ExceptionTypeD_Out_T_5}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_8 = _ExceptionTypeD_Out_T_4 | _GEN_12; // @[Mux.scala 27:73]
  wire [20:0] _GEN_13 = {{18'd0}, _ExceptionTypeD_Out_T_6}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_9 = _ExceptionTypeD_Out_T_8 | _GEN_13; // @[Mux.scala 27:73]
  wire [24:0] _GEN_14 = {{4'd0}, _ExceptionTypeD_Out_T_9}; // @[Mux.scala 27:73]
  wire [24:0] _ExceptionTypeD_Out_T_10 = _GEN_14 | _ExceptionTypeD_Out_T_7; // @[Mux.scala 27:73]
  reg  int_instanceE_timer; // @[myCPU.scala 764:33]
  reg  int_instanceE_out_int; // @[myCPU.scala 764:33]
  reg  int_instanceM_timer; // @[myCPU.scala 765:33]
  reg  int_instanceM_out_int; // @[myCPU.scala 765:33]
  reg  int_instanceM2_timer; // @[myCPU.scala 766:33]
  reg  int_instanceM2_out_int; // @[myCPU.scala 766:33]
  reg  int_instanceW_timer; // @[myCPU.scala 767:33]
  reg  int_instanceW_out_int; // @[myCPU.scala 767:33]
  wire [2:0] _CalCsrDataE_T = _id2ex_io_csr_controlE; // @[myCPU.scala 944:31]
  wire [63:0] _Forward_csr_data_T_1 = 2'h1 == _cfu_io_ForwardcsrE ? _ex2mem_io_WriteDataM : _csr_io_csr_read_data; // @[Mux.scala 81:58]
  wire [63:0] Forward_csr_data = 2'h2 == _cfu_io_ForwardcsrE ? _mem2mem2_io_WriteDataM : _Forward_csr_data_T_1; // @[Mux.scala 81:58]
  wire [4:0] _csr_src1_T = _id2ex_io_R1E; // @[macros.scala 443:38]
  wire [5:0] _csr_src1_T_1 = {1'h0,_csr_src1_T}; // @[Cat.scala 31:58]
  reg  Forward_Lock1E; // @[myCPU.scala 831:34]
  reg [63:0] RD1ForWardE_r; // @[myCPU.scala 829:34]
  wire [63:0] ResultW = _mem22wb_io_ResultW; // @[myCPU.scala 1148:15 296:26]
  wire [63:0] _RD1ForWardE_p_T_1 = 2'h1 == _cfu_io_Forward1E ? ResultW : _id2ex_io_RD1E; // @[Mux.scala 81:58]
  wire [63:0] _RD1ForWardE_p_T_3 = 2'h2 == _cfu_io_Forward1E ? resultE2M_Reg : _RD1ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [63:0] RD1ForWardE_p = 2'h3 == _cfu_io_Forward1E ? ResultM2_Reg : _RD1ForWardE_p_T_3; // @[Mux.scala 81:58]
  wire [63:0] RD1ForWardE = Forward_Lock1E ? RD1ForWardE_r : RD1ForWardE_p; // @[myCPU.scala 837:23]
  wire [63:0] csr_src1 = _id2ex_io_csr_ImmE ? {{58'd0}, _csr_src1_T_1} : RD1ForWardE; // @[myCPU.scala 941:20]
  wire [63:0] _CalCsrDataE_T_2 = Forward_csr_data | csr_src1; // @[myCPU.scala 944:64]
  wire [63:0] _CalCsrDataE_T_9 = _CalCsrDataE_T[0] ? _CalCsrDataE_T_2 : 64'h0; // @[Mux.scala 27:73]
  wire [2:0] _CalCsrDataE_T_3 = {{1'd0}, _id2ex_io_csr_controlE[2:1]}; // @[myCPU.scala 945:31]
  wire [63:0] _CalCsrDataE_T_5 = ~csr_src1; // @[myCPU.scala 945:68]
  wire [63:0] _CalCsrDataE_T_6 = Forward_csr_data & _CalCsrDataE_T_5; // @[myCPU.scala 945:64]
  wire [63:0] _CalCsrDataE_T_10 = _CalCsrDataE_T_3[0] ? _CalCsrDataE_T_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _CalCsrDataE_T_12 = _CalCsrDataE_T_9 | _CalCsrDataE_T_10; // @[Mux.scala 27:73]
  wire [2:0] _CalCsrDataE_T_7 = {{2'd0}, _id2ex_io_csr_controlE[2]}; // @[myCPU.scala 946:31]
  wire [63:0] _CalCsrDataE_T_11 = _CalCsrDataE_T_7[0] ? csr_src1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] CalCsrDataE = _CalCsrDataE_T_12 | _CalCsrDataE_T_11; // @[Mux.scala 27:73]
  wire  _int_disable_T_11 = _ex2mem_io_WritecsrAddrM == 12'h300 & _ex2mem_io_csrWriteM & ~_ex2mem_io_CsrWritedataM[3]; // @[myCPU.scala 772:95]
  wire  _int_disable_T_12 = _id2ex_io2_WritecsrAddrE == 12'h300 & _id2ex_io2_csrWriteE & ~CalCsrDataE[3] |
    _int_disable_T_11; // @[myCPU.scala 771:126]
  wire  _int_disable_T_18 = _mem2mem2_io_WritecsrAddrM == 12'h300 & _mem2mem2_io_csrWriteM & ~_mem2mem2_io_CsrWritedataM
    [3]; // @[myCPU.scala 773:99]
  wire  _int_disable_T_19 = _int_disable_T_12 | _int_disable_T_18; // @[myCPU.scala 772:140]
  wire  _int_disable_T_25 = _csr_io_csr_write_addr == 12'h300 & _csr_io_csr_write_en & ~_csr_io_csr_write_data[3]; // @[myCPU.scala 774:93]
  wire  int_disable = _int_disable_T_19 | _int_disable_T_25; // @[myCPU.scala 773:145]
  wire  _ext_int_with_enable_timer_T = ext_int_timer & _csr_io_int_type_able_timer; // @[myCPU.scala 777:48]
  wire  _ext_int_with_enable_timer_T_2 = ~int_disable; // @[myCPU.scala 777:102]
  wire  ext_int_with_enable_timer = ext_int_timer & _csr_io_int_type_able_timer & _csr_io_Int_able & ~int_disable; // @[myCPU.scala 777:99]
  wire  ext_int_with_enable_out_int = ext_int_out_int & _csr_io_int_type_out_int & _csr_io_Int_able &
    _ext_int_with_enable_timer_T_2; // @[myCPU.scala 778:100]
  wire  __id2ex_io_ExceptionTypeD_T_1 = ext_int_out_int & _csr_io_int_type_able_out_int; // @[myCPU.scala 790:26]
  wire  __id2ex_io_ExceptionTypeD_T_2 = _ext_int_with_enable_timer_T | __id2ex_io_ExceptionTypeD_T_1; // @[myCPU.scala 789:86]
  wire  __id2ex_io_ExceptionTypeD_T_6 = __id2ex_io_ExceptionTypeD_T_2 & _csr_io_Int_able &
    _ext_int_with_enable_timer_T_2; // @[myCPU.scala 790:88]
  wire [31:0] ExceptionTypeD_Out = {{7'd0}, _ExceptionTypeD_Out_T_10}; // @[myCPU.scala 190:34 754:24]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_9 = __if2id_io_InstrF_T ? 11'h400 : 11'h0; // @[myCPU.scala 791:13]
  wire [8:0] __id2ex_io_ExceptionTypeD_T_11 = __if2id_io_InstrF_T_1 ? 9'h100 : 9'h0; // @[myCPU.scala 792:13]
  wire [10:0] _GEN_17 = {{2'd0}, __id2ex_io_ExceptionTypeD_T_11}; // @[myCPU.scala 791:59]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_12 = __id2ex_io_ExceptionTypeD_T_9 | _GEN_17; // @[myCPU.scala 791:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_14 = __if2id_io_InstrF_T_3 ? 32'h80000000 : 32'h0; // @[myCPU.scala 794:13]
  wire [31:0] _GEN_18 = {{21'd0}, __id2ex_io_ExceptionTypeD_T_12}; // @[myCPU.scala 792:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_15 = _GEN_18 | __id2ex_io_ExceptionTypeD_T_14; // @[myCPU.scala 792:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_16 = ExceptionTypeD_Out == 32'h0 ? __id2ex_io_ExceptionTypeD_T_15 :
    ExceptionTypeD_Out; // @[myCPU.scala 790:122]
  reg  inst_tlb_exceptionM; // @[myCPU.scala 824:34]
  wire [63:0] _RD2ForWardE_p_T_1 = 2'h1 == _cfu_io_Forward2E ? ResultW : _id2ex_io_RD2E; // @[Mux.scala 81:58]
  wire [63:0] _RD2ForWardE_p_T_3 = 2'h2 == _cfu_io_Forward2E ? resultE2M_Reg : _RD2ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [63:0] RD2ForWardE_p = 2'h3 == _cfu_io_Forward2E ? ResultM2_Reg : _RD2ForWardE_p_T_3; // @[Mux.scala 81:58]
  reg [63:0] RD2ForWardE_r; // @[myCPU.scala 830:34]
  reg  Forward_Lock2E; // @[myCPU.scala 832:34]
  wire [63:0] RD2ForWardE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 838:23]
  wire  _Forward_Lock1E_T = _ex2mem_io_MemToRegM; // @[myCPU.scala 844:54]
  wire  _Forward_Lock1E_T_1 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 844:87]
  wire  _Forward_Lock1E_T_3 = ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM); // @[myCPU.scala 844:31]
  wire [63:0] Src1E = _id2ex_io2_ALUSrcE_0 ? _id2ex_io2_PCE : RD1ForWardE; // @[myCPU.scala 859:20]
  wire [63:0] Src2E = _id2ex_io2_ALUSrcE_1 ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 866:20]
  wire  csrToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_csrToRegE_Out; // @[myCPU.scala 870:24]
  wire  __muldiv_io_en_T_2 = _ex2mem_io_RegWriteM; // @[myCPU.scala 877:105]
  wire  __muldiv_io_en_T_10 = _id2ex_io_R1E == _ex2mem_io_WriteRegM & __muldiv_io_en_T_2 & _Forward_Lock1E_T; // @[myCPU.scala 878:88]
  wire  __muldiv_io_en_T_11 = _id2ex_io_R2E == _ex2mem_io_WriteRegM & _ex2mem_io_RegWriteM & _Forward_Lock1E_T |
    __muldiv_io_en_T_10; // @[myCPU.scala 877:144]
  wire  __muldiv_io_en_T_13 = _mem2mem2_io_RegWriteM; // @[myCPU.scala 879:85]
  wire  __muldiv_io_en_T_16 = _id2ex_io_R2E == _mem2mem2_io_WriteRegM & _mem2mem2_io_RegWriteM & _Forward_Lock1E_T_1; // @[myCPU.scala 879:92]
  wire  __muldiv_io_en_T_17 = __muldiv_io_en_T_11 | __muldiv_io_en_T_16; // @[myCPU.scala 878:120]
  wire  __muldiv_io_en_T_22 = _id2ex_io_R1E == _mem2mem2_io_WriteRegM & __muldiv_io_en_T_13 & _Forward_Lock1E_T_1; // @[myCPU.scala 880:92]
  wire  __muldiv_io_en_T_23 = __muldiv_io_en_T_17 | __muldiv_io_en_T_22; // @[myCPU.scala 879:126]
  wire [12:0] _temp_exceptionE_T_11 = _alu_io_overflow ? 13'h1000 : 13'h0; // @[myCPU.scala 911:13]
  wire  _resultE_T_1 = _id2ex_io2_LinkE; // @[myCPU.scala 959:25]
  wire [63:0] _resultE_T_2 = _id2ex_io_alu_calE ? _alu_io_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_3 = csrToRegE ? Forward_csr_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_4 = _resultE_T_1 ? _id2ex_io2_PCPlus4E : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_5 = _id2ex_io_muldiv_calE ? _muldiv_io_data_out : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_6 = _resultE_T_2 | _resultE_T_3; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_7 = _resultE_T_6 | _resultE_T_4; // @[Mux.scala 27:73]
  wire [63:0] resultE = _resultE_T_7 | _resultE_T_5; // @[Mux.scala 27:73]
  reg  tlb_exception_csr_writeM2; // @[myCPU.scala 1063:40]
  reg  tlb_exception_co0_writeW; // @[myCPU.scala 1064:40]
  wire [63:0] Mem_withRL_Data = _dmem_io_RD; // @[myCPU.scala 1083:34 1090:21]
  wire  csrWriteW = wb_exception ? 1'h0 : _mem22wb_io_csrWriteW; // @[myCPU.scala 1151:25]
  wire [63:0] __addr_cal_io_d_vaddr_T_1 = _id2ex_io_ImmE + RD1ForWardE; // @[myCPU.scala 1185:44]
  wire [31:0] inst_buffer_read_out_pc = fifo_with_bundle_io_read_out_0_pc; // @[myCPU.scala 583:36 584:26]
  wire [31:0] inst_buffer_read_out_pre_pc_target = fifo_with_bundle_io_read_out_0_pre_pc_target; // @[myCPU.scala 583:36 584:26]
  ysyx_22040886_alu _alu ( // @[myCPU.scala 118:22]
    .io_ctrl(_alu_io_ctrl),
    .io_in1(_alu_io_in1),
    .io_in2(_alu_io_in2),
    .io_result(_alu_io_result),
    .io_overflow(_alu_io_overflow),
    .io_data_w(_alu_io_data_w)
  );
  ysyx_22040886_br _br ( // @[myCPU.scala 119:22]
    .reset(_br_reset),
    .io_r1(_br_io_r1),
    .io_r2(_br_io_r2),
    .io_branch(_br_io_branch),
    .io_exe(_br_io_exe)
  );
  ysyx_22040886_cfu _cfu ( // @[myCPU.scala 120:22]
    .reset(_cfu_reset),
    .io_Inst_Fifo_Empty(_cfu_io_Inst_Fifo_Empty),
    .io_dmem_calD(_cfu_io_dmem_calD),
    .io_BranchD_Flag(_cfu_io_BranchD_Flag),
    .io_JRD(_cfu_io_JRD),
    .io_CanBranchD(_cfu_io_CanBranchD),
    .io_DivPendingE(_cfu_io_DivPendingE),
    .io_DataPendingM(_cfu_io_DataPendingM),
    .io_InException(_cfu_io_InException),
    .io_WriteRegE(_cfu_io_WriteRegE),
    .io_RegWriteE(_cfu_io_RegWriteE),
    .io_csrToRegE(_cfu_io_csrToRegE),
    .io_WriteRegM(_cfu_io_WriteRegM),
    .io_MemToRegM(_cfu_io_MemToRegM),
    .io_RegWriteM(_cfu_io_RegWriteM),
    .io_csrWriteM(_cfu_io_csrWriteM),
    .io_WriteRegM2(_cfu_io_WriteRegM2),
    .io_MemToRegM2(_cfu_io_MemToRegM2),
    .io_RegWriteM2(_cfu_io_RegWriteM2),
    .io_csrWriteM2(_cfu_io_csrWriteM2),
    .io_WriteRegW(_cfu_io_WriteRegW),
    .io_RegWriteW(_cfu_io_RegWriteW),
    .io_ReadcsrAddrE(_cfu_io_ReadcsrAddrE),
    .io_WritecsrAddrM(_cfu_io_WritecsrAddrM),
    .io_WritecsrAddrM2(_cfu_io_WritecsrAddrM2),
    .io_R2D(_cfu_io_R2D),
    .io_R1D(_cfu_io_R1D),
    .io_R2E(_cfu_io_R2E),
    .io_R1E(_cfu_io_R1E),
    .io_StallF(_cfu_io_StallF),
    .io_StallD(_cfu_io_StallD),
    .io_StallE(_cfu_io_StallE),
    .io_StallM(_cfu_io_StallM),
    .io_StallM2(_cfu_io_StallM2),
    .io_StallW(_cfu_io_StallW),
    .io_FlushD(_cfu_io_FlushD),
    .io_FlushE(_cfu_io_FlushE),
    .io_FlushM(_cfu_io_FlushM),
    .io_FlushM2(_cfu_io_FlushM2),
    .io_FlushW(_cfu_io_FlushW),
    .io_Forward1E(_cfu_io_Forward1E),
    .io_Forward2E(_cfu_io_Forward2E),
    .io_Forward1D(_cfu_io_Forward1D),
    .io_Forward2D(_cfu_io_Forward2D),
    .io_ForwardcsrE(_cfu_io_ForwardcsrE)
  );
  ysyx_22040886_csr _csr ( // @[myCPU.scala 121:22]
    .clock(_csr_clock),
    .reset(_csr_reset),
    .io_csr_read_addr(_csr_io_csr_read_addr),
    .io_csr_write_addr(_csr_io_csr_write_addr),
    .io_csr_write_data(_csr_io_csr_write_data),
    .io_csr_write_en(_csr_io_csr_write_en),
    .io_pc(_csr_io_pc),
    .io_exception_type_i(_csr_io_exception_type_i),
    .io_return_pc(_csr_io_return_pc),
    .io_exception(_csr_io_exception),
    .io_csr_read_data(_csr_io_csr_read_data),
    .io_icache_tags_flush(_csr_io_icache_tags_flush),
    .io_int_type_timer(_csr_io_int_type_timer),
    .io_int_type_out_int(_csr_io_int_type_out_int),
    .io_stageW_pc(_csr_io_stageW_pc),
    .io_Int_able(_csr_io_Int_able),
    .io_int_type_able_timer(_csr_io_int_type_able_timer),
    .io_int_type_able_out_int(_csr_io_int_type_able_out_int)
  );
  ysyx_22040886_cu _cu ( // @[myCPU.scala 122:22]
    .io1_InstrD(_cu_io1_InstrD),
    .io1_BadInstrD(_cu_io1_BadInstrD),
    .io1_SysCallD(_cu_io1_SysCallD),
    .io1_EretD(_cu_io1_EretD),
    .io1_dmem_addr_cal(_cu_io1_dmem_addr_cal),
    .io_RegWriteD(_cu_io_RegWriteD),
    .io_MemToRegD(_cu_io_MemToRegD),
    .io_MemWriteD(_cu_io_MemWriteD),
    .io_ALUCtrlD(_cu_io_ALUCtrlD),
    .io_ALUSrcD_0(_cu_io_ALUSrcD_0),
    .io_ALUSrcD_1(_cu_io_ALUSrcD_1),
    .io_RegDstD(_cu_io_RegDstD),
    .io_LinkD(_cu_io_LinkD),
    .io_csrWriteD(_cu_io_csrWriteD),
    .io_csrToRegD(_cu_io_csrToRegD),
    .io_LoadUnsignedD(_cu_io_LoadUnsignedD),
    .io_MemWidthD(_cu_io_MemWidthD),
    .io_ImmD(_cu_io_ImmD),
    .io_data_wD(_cu_io_data_wD),
    .io_muldiv_control(_cu_io_muldiv_control),
    .io_muldiv_cal(_cu_io_muldiv_cal),
    .io_alu_cal(_cu_io_alu_cal),
    .io_csr_control(_cu_io_csr_control),
    .io_csr_Imm(_cu_io_csr_Imm),
    .io_fence_i_control(_cu_io_fence_i_control)
  );
  ysyx_22040886_dmem _dmem ( // @[myCPU.scala 123:23]
    .io_data_ok(_dmem_io_data_ok),
    .io_rdata(_dmem_io_rdata),
    .io_Physisc_Address(_dmem_io_Physisc_Address),
    .io_WIDTH(_dmem_io_WIDTH),
    .io_SIGN(_dmem_io_SIGN),
    .io_RD(_dmem_io_RD),
    .io_data_pending(_dmem_io_data_pending)
  );
  ysyx_22040886_dmemreq _dmemreq ( // @[myCPU.scala 124:26]
    .io_en(_dmemreq_io_en),
    .io_MemWriteE(_dmemreq_io_MemWriteE),
    .io_MemToRegE(_dmemreq_io_MemToRegE),
    .io_MemWidthE(_dmemreq_io_MemWidthE),
    .io_VAddrE(_dmemreq_io_VAddrE),
    .io_WriteDataE(_dmemreq_io_WriteDataE),
    .io_req(_dmemreq_io_req),
    .io_wr(_dmemreq_io_wr),
    .io_size(_dmemreq_io_size),
    .io_addr(_dmemreq_io_addr),
    .io_wdata(_dmemreq_io_wdata),
    .io_wstrb(_dmemreq_io_wstrb)
  );
  ysyx_22040886_ex2mem _ex2mem ( // @[myCPU.scala 125:26]
    .clock(_ex2mem_clock),
    .reset(_ex2mem_reset),
    .io1_RegWriteE(_ex2mem_io1_RegWriteE),
    .io1_MemToRegE(_ex2mem_io1_MemToRegE),
    .io1_LoadUnsignedE(_ex2mem_io1_LoadUnsignedE),
    .io1_MemWidthE(_ex2mem_io1_MemWidthE),
    .io1_csrWriteE(_ex2mem_io1_csrWriteE),
    .io1_WritecsrAddrE(_ex2mem_io1_WritecsrAddrE),
    .io1_PCE(_ex2mem_io1_PCE),
    .io1_BranchJump_JrE(_ex2mem_io1_BranchJump_JrE),
    .io_en(_ex2mem_io_en),
    .io_clr(_ex2mem_io_clr),
    .io_WriteDataE(_ex2mem_io_WriteDataE),
    .io_WriteRegE(_ex2mem_io_WriteRegE),
    .io_PhyAddrE(_ex2mem_io_PhyAddrE),
    .io_CsrWritedataE(_ex2mem_io_CsrWritedataE),
    .io_ExceptionTypeE(_ex2mem_io_ExceptionTypeE),
    .io_RegWriteM(_ex2mem_io_RegWriteM),
    .io_MemToRegM(_ex2mem_io_MemToRegM),
    .io_WriteDataM(_ex2mem_io_WriteDataM),
    .io_WriteRegM(_ex2mem_io_WriteRegM),
    .io_LoadUnsignedM(_ex2mem_io_LoadUnsignedM),
    .io_MemWidthM(_ex2mem_io_MemWidthM),
    .io_PhyAddrM(_ex2mem_io_PhyAddrM),
    .io_csrWriteM(_ex2mem_io_csrWriteM),
    .io_WritecsrAddrM(_ex2mem_io_WritecsrAddrM),
    .io_PCM(_ex2mem_io_PCM),
    .io_ExceptionTypeM_Out(_ex2mem_io_ExceptionTypeM_Out),
    .io_BranchJump_JrM(_ex2mem_io_BranchJump_JrM),
    .io_CsrWritedataM(_ex2mem_io_CsrWritedataM)
  );
  ysyx_22040886_ex2mem _mem2mem2 ( // @[myCPU.scala 126:28]
    .clock(_mem2mem2_clock),
    .reset(_mem2mem2_reset),
    .io1_RegWriteE(_mem2mem2_io1_RegWriteE),
    .io1_MemToRegE(_mem2mem2_io1_MemToRegE),
    .io1_LoadUnsignedE(_mem2mem2_io1_LoadUnsignedE),
    .io1_MemWidthE(_mem2mem2_io1_MemWidthE),
    .io1_csrWriteE(_mem2mem2_io1_csrWriteE),
    .io1_WritecsrAddrE(_mem2mem2_io1_WritecsrAddrE),
    .io1_PCE(_mem2mem2_io1_PCE),
    .io1_BranchJump_JrE(_mem2mem2_io1_BranchJump_JrE),
    .io_en(_mem2mem2_io_en),
    .io_clr(_mem2mem2_io_clr),
    .io_WriteDataE(_mem2mem2_io_WriteDataE),
    .io_WriteRegE(_mem2mem2_io_WriteRegE),
    .io_PhyAddrE(_mem2mem2_io_PhyAddrE),
    .io_CsrWritedataE(_mem2mem2_io_CsrWritedataE),
    .io_ExceptionTypeE(_mem2mem2_io_ExceptionTypeE),
    .io_RegWriteM(_mem2mem2_io_RegWriteM),
    .io_MemToRegM(_mem2mem2_io_MemToRegM),
    .io_WriteDataM(_mem2mem2_io_WriteDataM),
    .io_WriteRegM(_mem2mem2_io_WriteRegM),
    .io_LoadUnsignedM(_mem2mem2_io_LoadUnsignedM),
    .io_MemWidthM(_mem2mem2_io_MemWidthM),
    .io_PhyAddrM(_mem2mem2_io_PhyAddrM),
    .io_csrWriteM(_mem2mem2_io_csrWriteM),
    .io_WritecsrAddrM(_mem2mem2_io_WritecsrAddrM),
    .io_PCM(_mem2mem2_io_PCM),
    .io_ExceptionTypeM_Out(_mem2mem2_io_ExceptionTypeM_Out),
    .io_BranchJump_JrM(_mem2mem2_io_BranchJump_JrM),
    .io_CsrWritedataM(_mem2mem2_io_CsrWritedataM)
  );
  ysyx_22040886_id2ex _id2ex ( // @[myCPU.scala 128:26]
    .clock(_id2ex_clock),
    .reset(_id2ex_reset),
    .io1_RegWriteD(_id2ex_io1_RegWriteD),
    .io1_MemToRegD(_id2ex_io1_MemToRegD),
    .io1_MemWriteD(_id2ex_io1_MemWriteD),
    .io1_ALUCtrlD(_id2ex_io1_ALUCtrlD),
    .io1_ALUSrcD_0(_id2ex_io1_ALUSrcD_0),
    .io1_ALUSrcD_1(_id2ex_io1_ALUSrcD_1),
    .io1_RegDstD(_id2ex_io1_RegDstD),
    .io1_LinkD(_id2ex_io1_LinkD),
    .io1_csrWriteD(_id2ex_io1_csrWriteD),
    .io1_csrToRegD(_id2ex_io1_csrToRegD),
    .io1_LoadUnsignedD(_id2ex_io1_LoadUnsignedD),
    .io1_MemWidthD(_id2ex_io1_MemWidthD),
    .io1_data_wD(_id2ex_io1_data_wD),
    .io1_muldiv_control(_id2ex_io1_muldiv_control),
    .io1_muldiv_cal(_id2ex_io1_muldiv_cal),
    .io1_alu_cal(_id2ex_io1_alu_cal),
    .io1_csr_control(_id2ex_io1_csr_control),
    .io1_csr_Imm(_id2ex_io1_csr_Imm),
    .io1_fence_i_control(_id2ex_io1_fence_i_control),
    .io2_RegWriteE(_id2ex_io2_RegWriteE),
    .io2_MemToRegE(_id2ex_io2_MemToRegE),
    .io2_MemWriteE(_id2ex_io2_MemWriteE),
    .io2_ALUCtrlE(_id2ex_io2_ALUCtrlE),
    .io2_ALUSrcE_0(_id2ex_io2_ALUSrcE_0),
    .io2_ALUSrcE_1(_id2ex_io2_ALUSrcE_1),
    .io2_RegDstE(_id2ex_io2_RegDstE),
    .io2_LinkE(_id2ex_io2_LinkE),
    .io2_PCPlus4E(_id2ex_io2_PCPlus4E),
    .io2_LoadUnsignedE(_id2ex_io2_LoadUnsignedE),
    .io2_MemWidthE(_id2ex_io2_MemWidthE),
    .io2_csrWriteE(_id2ex_io2_csrWriteE),
    .io2_WritecsrAddrE(_id2ex_io2_WritecsrAddrE),
    .io2_ReadcsrAddrE(_id2ex_io2_ReadcsrAddrE),
    .io2_PCE(_id2ex_io2_PCE),
    .io2_BranchJump_JrE(_id2ex_io2_BranchJump_JrE),
    .io_en(_id2ex_io_en),
    .io_clr(_id2ex_io_clr),
    .io_csrToRegE_Out(_id2ex_io_csrToRegE_Out),
    .io_RD1D(_id2ex_io_RD1D),
    .io_RD2D(_id2ex_io_RD2D),
    .io_R2D(_id2ex_io_R2D),
    .io_R1D(_id2ex_io_R1D),
    .io_ImmD(_id2ex_io_ImmD),
    .io_PCPlus4D(_id2ex_io_PCPlus4D),
    .io_WritecsrAddrD(_id2ex_io_WritecsrAddrD),
    .io_ReadcsrAddrD(_id2ex_io_ReadcsrAddrD),
    .io_PCD(_id2ex_io_PCD),
    .io_ExceptionTypeD(_id2ex_io_ExceptionTypeD),
    .io_BranchJump_JrD(_id2ex_io_BranchJump_JrD),
    .io_RD1E(_id2ex_io_RD1E),
    .io_RD2E(_id2ex_io_RD2E),
    .io_R2E(_id2ex_io_R2E),
    .io_R1E(_id2ex_io_R1E),
    .io_ImmE(_id2ex_io_ImmE),
    .io_data_wE(_id2ex_io_data_wE),
    .io_muldiv_control(_id2ex_io_muldiv_control),
    .io_alu_calE(_id2ex_io_alu_calE),
    .io_muldiv_calE(_id2ex_io_muldiv_calE),
    .io_ExceptionTypeE_Out(_id2ex_io_ExceptionTypeE_Out),
    .io_csr_controlE(_id2ex_io_csr_controlE),
    .io_csr_ImmE(_id2ex_io_csr_ImmE),
    .io_fence_i_controlE(_id2ex_io_fence_i_controlE)
  );
  ysyx_22040886_if2id _if2id ( // @[myCPU.scala 129:26]
    .clock(_if2id_clock),
    .reset(_if2id_reset),
    .io_en(_if2id_io_en),
    .io_clr(_if2id_io_clr),
    .io_InstrF(_if2id_io_InstrF),
    .io_PCPlus4F(_if2id_io_PCPlus4F),
    .io_PCF(_if2id_io_PCF),
    .io_ExceptionTypeF(_if2id_io_ExceptionTypeF),
    .io_InstrD(_if2id_io_InstrD),
    .io_PCPlus4D(_if2id_io_PCPlus4D),
    .io_PCD(_if2id_io_PCD),
    .io_ExceptionTypeD_Out(_if2id_io_ExceptionTypeD_Out)
  );
  ysyx_22040886_mem2wb _mem22wb ( // @[myCPU.scala 131:27]
    .clock(_mem22wb_clock),
    .reset(_mem22wb_reset),
    .io_en(_mem22wb_io_en),
    .io_clr(_mem22wb_io_clr),
    .io_RegWriteM(_mem22wb_io_RegWriteM),
    .io_ResultM(_mem22wb_io_ResultM),
    .io_WriteRegM(_mem22wb_io_WriteRegM),
    .io_csrWriteM(_mem22wb_io_csrWriteM),
    .io_WritecsrAddrM(_mem22wb_io_WritecsrAddrM),
    .io_CsrWritedataM(_mem22wb_io_CsrWritedataM),
    .io_PCM(_mem22wb_io_PCM),
    .io_ExceptionTypeM(_mem22wb_io_ExceptionTypeM),
    .io_BranchJump_JrM(_mem22wb_io_BranchJump_JrM),
    .io_RegWriteW_Out(_mem22wb_io_RegWriteW_Out),
    .io_ResultW(_mem22wb_io_ResultW),
    .io_WriteRegW(_mem22wb_io_WriteRegW),
    .io_csrWriteW(_mem22wb_io_csrWriteW),
    .io_WritecsrAddrW(_mem22wb_io_WritecsrAddrW),
    .io_PCW(_mem22wb_io_PCW),
    .io_ExceptionTypeW_Out(_mem22wb_io_ExceptionTypeW_Out),
    .io_BranchJump_JrW(_mem22wb_io_BranchJump_JrW),
    .io_CsrWritedataW(_mem22wb_io_CsrWritedataW)
  );
  ysyx_22040886_addr_cal _addr_cal ( // @[myCPU.scala 132:31]
    .io_d_vaddr(_addr_cal_io_d_vaddr),
    .io_d_paddr(_addr_cal_io_d_paddr),
    .io_d_cached(_addr_cal_io_d_cached)
  );
  ysyx_22040886_muldiv _muldiv ( // @[myCPU.scala 133:26]
    .clock(_muldiv_clock),
    .reset(_muldiv_reset),
    .io_en(_muldiv_io_en),
    .io_ctrl(_muldiv_io_ctrl),
    .io_in1(_muldiv_io_in1),
    .io_in2(_muldiv_io_in2),
    .io_data_out(_muldiv_io_data_out),
    .io_pending(_muldiv_io_pending)
  );
  ysyx_22040886_regfile _regfile ( // @[myCPU.scala 135:26]
    .clock(_regfile_clock),
    .reset(_regfile_reset),
    .io_A1(_regfile_io_A1),
    .io_A2(_regfile_io_A2),
    .io_WE3(_regfile_io_WE3),
    .io_A3(_regfile_io_A3),
    .io_WD3(_regfile_io_WD3),
    .io_RD1(_regfile_io_RD1),
    .io_RD2(_regfile_io_RD2)
  );
  ysyx_22040886_fifo_with_bundle fifo_with_bundle ( // @[myCPU.scala 157:29]
    .clock(fifo_with_bundle_clock),
    .reset(fifo_with_bundle_reset),
    .io_read_en(fifo_with_bundle_io_read_en),
    .io_write_en(fifo_with_bundle_io_write_en),
    .io_read_out_0_pc(fifo_with_bundle_io_read_out_0_pc),
    .io_read_out_0_inst(fifo_with_bundle_io_read_out_0_inst),
    .io_read_out_0_exception_type(fifo_with_bundle_io_read_out_0_exception_type),
    .io_read_out_0_pre_pc_target(fifo_with_bundle_io_read_out_0_pre_pc_target),
    .io_read_out_0_pre_lookup_data(fifo_with_bundle_io_read_out_0_pre_lookup_data),
    .io_read_out_0_pre_hashcode(fifo_with_bundle_io_read_out_0_pre_hashcode),
    .io_read_out_0_pre_pht(fifo_with_bundle_io_read_out_0_pre_pht),
    .io_read_out_0_pre_bht(fifo_with_bundle_io_read_out_0_pre_bht),
    .io_read_out_0_pre_decoder_branchD_flag(fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag),
    .io_read_out_0_pre_decoder_jump(fifo_with_bundle_io_read_out_0_pre_decoder_jump),
    .io_read_out_0_pre_decoder_branchdata(fifo_with_bundle_io_read_out_0_pre_decoder_branchdata),
    .io_read_out_0_pre_decoder_jr(fifo_with_bundle_io_read_out_0_pre_decoder_jr),
    .io_read_out_0_true_branch_state(fifo_with_bundle_io_read_out_0_true_branch_state),
    .io_write_in_0_pc(fifo_with_bundle_io_write_in_0_pc),
    .io_write_in_0_inst(fifo_with_bundle_io_write_in_0_inst),
    .io_write_in_0_pre_pc_target(fifo_with_bundle_io_write_in_0_pre_pc_target),
    .io_write_in_0_pre_lookup_data(fifo_with_bundle_io_write_in_0_pre_lookup_data),
    .io_write_in_0_pre_hashcode(fifo_with_bundle_io_write_in_0_pre_hashcode),
    .io_write_in_0_pre_pht(fifo_with_bundle_io_write_in_0_pre_pht),
    .io_write_in_0_pre_bht(fifo_with_bundle_io_write_in_0_pre_bht),
    .io_write_in_0_pre_decoder_branchD_flag(fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag),
    .io_write_in_0_pre_decoder_jump(fifo_with_bundle_io_write_in_0_pre_decoder_jump),
    .io_write_in_0_pre_decoder_branchdata(fifo_with_bundle_io_write_in_0_pre_decoder_branchdata),
    .io_write_in_0_pre_decoder_jr(fifo_with_bundle_io_write_in_0_pre_decoder_jr),
    .io_write_in_0_true_branch_state(fifo_with_bundle_io_write_in_0_true_branch_state),
    .io_full(fifo_with_bundle_io_full),
    .io_empty(fifo_with_bundle_io_empty),
    .io_point_write_en(fifo_with_bundle_io_point_write_en),
    .io_point_flush(fifo_with_bundle_io_point_flush)
  );
  ysyx_22040886_pc_detail stage_fec_1_pc_L ( // @[myCPU.scala 423:34]
    .clock(stage_fec_1_pc_L_clock),
    .reset(stage_fec_1_pc_L_reset),
    .io_stall(stage_fec_1_pc_L_io_stall),
    .io_flush(stage_fec_1_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_L_io_out_pc_value_out)
  );
  ysyx_22040886_branch_prediction branch_prediction ( // @[myCPU.scala 447:21]
    .clock(branch_prediction_clock),
    .reset(branch_prediction_reset),
    .io_pc(branch_prediction_io_pc),
    .io_write_pc(branch_prediction_io_write_pc),
    .io_aw_pht_ways_addr(branch_prediction_io_aw_pht_ways_addr),
    .io_aw_pht_addr(branch_prediction_io_aw_pht_addr),
    .io_aw_bht_addr(branch_prediction_io_aw_bht_addr),
    .io_aw_target_addr(branch_prediction_io_aw_target_addr),
    .io_btb_write(branch_prediction_io_btb_write),
    .io_bht_write(branch_prediction_io_bht_write),
    .io_pht_write(branch_prediction_io_pht_write),
    .io_bht_in(branch_prediction_io_bht_in),
    .io_pht_in(branch_prediction_io_pht_in),
    .io_out(branch_prediction_io_out),
    .io_pre(branch_prediction_io_pre),
    .io_bht(branch_prediction_io_bht),
    .io_btb_hit(branch_prediction_io_btb_hit),
    .io_pre_target(branch_prediction_io_pre_target),
    .io_stage2_stall(branch_prediction_io_stage2_stall),
    .io_stage2_flush(branch_prediction_io_stage2_flush),
    .io_lookup_data(branch_prediction_io_lookup_data)
  );
  ysyx_22040886_pc_detail stage_fec_2_pc_L ( // @[myCPU.scala 509:34]
    .clock(stage_fec_2_pc_L_clock),
    .reset(stage_fec_2_pc_L_reset),
    .io_stall(stage_fec_2_pc_L_io_stall),
    .io_flush(stage_fec_2_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_L_io_out_pc_value_out)
  );
  ysyx_22040886_bru_detail id_bru_state ( // @[myCPU.scala 666:31]
    .clock(id_bru_state_clock),
    .reset(id_bru_state_reset),
    .io_stall(id_bru_state_io_stall),
    .io_flush(id_bru_state_io_flush),
    .io_in_pht(id_bru_state_io_in_pht),
    .io_in_bht(id_bru_state_io_in_bht),
    .io_in_hashcode(id_bru_state_io_in_hashcode),
    .io_in_target_pc(id_bru_state_io_in_target_pc),
    .io_in_lookup_data(id_bru_state_io_in_lookup_data),
    .io_out_pht(id_bru_state_io_out_pht),
    .io_out_bht(id_bru_state_io_out_bht),
    .io_out_hashcode(id_bru_state_io_out_hashcode),
    .io_out_target_pc(id_bru_state_io_out_target_pc),
    .io_out_lookup_data(id_bru_state_io_out_lookup_data)
  );
  ysyx_22040886_bru_detail ex_bru_state ( // @[myCPU.scala 670:31]
    .clock(ex_bru_state_clock),
    .reset(ex_bru_state_reset),
    .io_stall(ex_bru_state_io_stall),
    .io_flush(ex_bru_state_io_flush),
    .io_in_pht(ex_bru_state_io_in_pht),
    .io_in_bht(ex_bru_state_io_in_bht),
    .io_in_hashcode(ex_bru_state_io_in_hashcode),
    .io_in_target_pc(ex_bru_state_io_in_target_pc),
    .io_in_lookup_data(ex_bru_state_io_in_lookup_data),
    .io_out_pht(ex_bru_state_io_out_pht),
    .io_out_bht(ex_bru_state_io_out_bht),
    .io_out_hashcode(ex_bru_state_io_out_hashcode),
    .io_out_target_pc(ex_bru_state_io_out_target_pc),
    .io_out_lookup_data(ex_bru_state_io_out_lookup_data)
  );
  ysyx_22040886_bru_detail mem_bru_state ( // @[myCPU.scala 674:32]
    .clock(mem_bru_state_clock),
    .reset(mem_bru_state_reset),
    .io_stall(mem_bru_state_io_stall),
    .io_flush(mem_bru_state_io_flush),
    .io_in_pht(mem_bru_state_io_in_pht),
    .io_in_bht(mem_bru_state_io_in_bht),
    .io_in_hashcode(mem_bru_state_io_in_hashcode),
    .io_in_target_pc(mem_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem_bru_state_io_in_lookup_data),
    .io_out_pht(mem_bru_state_io_out_pht),
    .io_out_bht(mem_bru_state_io_out_bht),
    .io_out_hashcode(mem_bru_state_io_out_hashcode),
    .io_out_target_pc(mem_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem_bru_state_io_out_lookup_data)
  );
  ysyx_22040886_bru_detail mem2_bru_state ( // @[myCPU.scala 678:33]
    .clock(mem2_bru_state_clock),
    .reset(mem2_bru_state_reset),
    .io_stall(mem2_bru_state_io_stall),
    .io_flush(mem2_bru_state_io_flush),
    .io_in_pht(mem2_bru_state_io_in_pht),
    .io_in_bht(mem2_bru_state_io_in_bht),
    .io_in_hashcode(mem2_bru_state_io_in_hashcode),
    .io_in_target_pc(mem2_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem2_bru_state_io_in_lookup_data),
    .io_out_pht(mem2_bru_state_io_out_pht),
    .io_out_bht(mem2_bru_state_io_out_bht),
    .io_out_hashcode(mem2_bru_state_io_out_hashcode),
    .io_out_target_pc(mem2_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem2_bru_state_io_out_lookup_data)
  );
  ysyx_22040886_bru_detail wb_bru_state ( // @[myCPU.scala 682:31]
    .clock(wb_bru_state_clock),
    .reset(wb_bru_state_reset),
    .io_stall(wb_bru_state_io_stall),
    .io_flush(wb_bru_state_io_flush),
    .io_in_pht(wb_bru_state_io_in_pht),
    .io_in_bht(wb_bru_state_io_in_bht),
    .io_in_hashcode(wb_bru_state_io_in_hashcode),
    .io_in_target_pc(wb_bru_state_io_in_target_pc),
    .io_in_lookup_data(wb_bru_state_io_in_lookup_data),
    .io_out_pht(wb_bru_state_io_out_pht),
    .io_out_bht(wb_bru_state_io_out_bht),
    .io_out_hashcode(wb_bru_state_io_out_hashcode),
    .io_out_target_pc(wb_bru_state_io_out_target_pc),
    .io_out_lookup_data(wb_bru_state_io_out_lookup_data)
  );
  assign inst_cache = inst_sram_addr[31:29] == 3'h4; // @[macros.scala 487:55]
  assign inst_sram_en = stage2_stall; // @[myCPU.scala 386:17]
  assign inst_sram_addr = _stage_fec_2_branch_answer_T_8 ? _csr_io_return_pc : _inst_sram_addr_T_3; // @[myCPU.scala 379:21]
  assign stage2_flush = fifo_with_bundle_io_point_write_en & _stage_fec_2_data_valid_T | _stage_fec_2_branch_answer_T_8; // @[myCPU.scala 562:72]
  assign stage1_valid_flush = _pc_next_wait_T | _stage_fec_2_branch_answer_T_8; // @[myCPU.scala 572:85]
  assign inst_ready_to_use = inst_sram_addr[1:0] == 2'h0; // @[myCPU.scala 387:41]
  assign inst_buffer_full = fifo_with_bundle_io_full; // @[myCPU.scala 581:22]
  assign data_sram_en = _dmemreq_io_req & ~_dmem_io_data_pending; // @[myCPU.scala 244:44]
  assign data_sram_wen = _dmemreq_io_wr; // @[myCPU.scala 250:13]
  assign data_size = _dmemreq_io_size; // @[myCPU.scala 1192:15]
  assign data_sram_addr = _dmemreq_io_addr; // @[myCPU.scala 246:15]
  assign data_sram_wdata = _dmemreq_io_wdata; // @[myCPU.scala 247:16]
  assign data_cache = _addr_cal_io_d_cached; // @[myCPU.scala 1191:63]
  assign data_wstrb = _dmemreq_io_wstrb; // @[myCPU.scala 248:16]
  assign data_fence_i_control = fence_i_controlMReg; // @[myCPU.scala 936:26]
  assign icache_tag_flush = _csr_io_icache_tags_flush; // @[myCPU.scala 1202:22]
  assign _alu_io_ctrl = _id2ex_io2_ALUCtrlE; // @[myCPU.scala 874:18]
  assign _alu_io_in1 = {Src1E[63:32],Src1E[31:0]}; // @[Cat.scala 31:58]
  assign _alu_io_in2 = {Src2E[63:32],Src2E[31:0]}; // @[Cat.scala 31:58]
  assign _alu_io_data_w = _id2ex_io_data_wE; // @[myCPU.scala 875:20]
  assign _br_reset = reset;
  assign _br_io_r1 = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 751:20]
  assign _br_io_r2 = _cfu_io_Forward2D[0] ? resultE2M_Reg : _BranchR2D_T_2; // @[myCPU.scala 753:20]
  assign _br_io_branch = pre_decoder_branchdata; // @[myCPU.scala 761:19]
  assign _cfu_reset = reset;
  assign _cfu_io_Inst_Fifo_Empty = fifo_with_bundle_io_empty; // @[myCPU.scala 565:29]
  assign _cfu_io_dmem_calD = _cu_io1_dmem_addr_cal; // @[myCPU.scala 818:23]
  assign _cfu_io_BranchD_Flag = pre_decoder_branchD_flag; // @[myCPU.scala 1224:26]
  assign _cfu_io_JRD = pre_decoder_jr; // @[myCPU.scala 1221:25]
  assign _cfu_io_CanBranchD = ~(id_exception | ex_exception | mem_exception | mem2_exception | wb_exception); // @[myCPU.scala 1222:111]
  assign _cfu_io_DivPendingE = _muldiv_io_pending; // @[myCPU.scala 1225:33]
  assign _cfu_io_DataPendingM = _dmem_io_data_pending; // @[myCPU.scala 1227:33]
  assign _cfu_io_InException = _csr_io_exception; // @[myCPU.scala 1215:25]
  assign _cfu_io_WriteRegE = _id2ex_io2_RegDstE; // @[myCPU.scala 1231:33]
  assign _cfu_io_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 1233:33]
  assign _cfu_io_csrToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_csrToRegE_Out; // @[myCPU.scala 870:24]
  assign _cfu_io_WriteRegM = _ex2mem_io_WriteRegM; // @[myCPU.scala 1237:33]
  assign _cfu_io_MemToRegM = _ex2mem_io_MemToRegM; // @[myCPU.scala 1238:33]
  assign _cfu_io_RegWriteM = _ex2mem_io_RegWriteM; // @[myCPU.scala 1239:33]
  assign _cfu_io_csrWriteM = _ex2mem_io_csrWriteM; // @[myCPU.scala 1240:33]
  assign _cfu_io_WriteRegM2 = _mem2mem2_io_WriteRegM; // @[myCPU.scala 1261:25]
  assign _cfu_io_MemToRegM2 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 1262:25]
  assign _cfu_io_RegWriteM2 = _mem2mem2_io_RegWriteM; // @[myCPU.scala 1263:25]
  assign _cfu_io_csrWriteM2 = _mem2mem2_io_csrWriteM; // @[myCPU.scala 1259:24]
  assign _cfu_io_WriteRegW = _mem22wb_io_WriteRegW; // @[myCPU.scala 1250:33]
  assign _cfu_io_RegWriteW = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1149:21]
  assign _cfu_io_ReadcsrAddrE = _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 1242:34]
  assign _cfu_io_WritecsrAddrM = _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 1245:34]
  assign _cfu_io_WritecsrAddrM2 = _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 1260:28]
  assign _cfu_io_R2D = _if2id_io_InstrD[24:20]; // @[myCPU.scala 203:27]
  assign _cfu_io_R1D = _if2id_io_InstrD[19:15]; // @[myCPU.scala 204:27]
  assign _cfu_io_R2E = _id2ex_io_R2E; // @[myCPU.scala 1256:33]
  assign _cfu_io_R1E = _id2ex_io_R1E; // @[myCPU.scala 1255:33]
  assign _csr_clock = clock;
  assign _csr_reset = reset;
  assign _csr_io_csr_read_addr = _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 952:27]
  assign _csr_io_csr_write_addr = _mem22wb_io_WritecsrAddrW; // @[myCPU.scala 953:28]
  assign _csr_io_csr_write_data = _mem22wb_io_CsrWritedataW; // @[myCPU.scala 1209:30]
  assign _csr_io_csr_write_en = csrWriteW | tlb_exception_co0_writeW; // @[myCPU.scala 1199:47]
  assign _csr_io_pc = _PCW_Reg_T ? _mem22wb_io_PCW : PCW_Reg; // @[myCPU.scala 1197:25]
  assign _csr_io_exception_type_i = _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 1200:30]
  assign _csr_io_int_type_timer = int_instanceW_timer; // @[myCPU.scala 1196:22]
  assign _csr_io_int_type_out_int = int_instanceW_out_int; // @[myCPU.scala 1196:22]
  assign _csr_io_stageW_pc = _mem22wb_io_PCW; // @[myCPU.scala 1210:30]
  assign _cu_io1_InstrD = _if2id_io_InstrD; // @[myCPU.scala 749:20]
  assign _dmem_io_data_ok = data_stage2_stall; // @[myCPU.scala 273:25]
  assign _dmem_io_rdata = data_sram_rdata; // @[myCPU.scala 274:25]
  assign _dmem_io_Physisc_Address = _mem2mem2_io_PhyAddrM[2:0]; // @[myCPU.scala 278:54]
  assign _dmem_io_WIDTH = _mem2mem2_io_MemWidthM; // @[myCPU.scala 276:25]
  assign _dmem_io_SIGN = ~_mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 277:22]
  assign _dmemreq_io_en = _T_34 ? 1'h0 : _commit_cache_reg_T; // @[myCPU.scala 892:26]
  assign _dmemreq_io_MemWriteE = _id2ex_io2_MemWriteE; // @[myCPU.scala 898:27]
  assign _dmemreq_io_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 895:27]
  assign _dmemreq_io_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 896:27]
  assign _dmemreq_io_VAddrE = _addr_cal_io_d_paddr; // @[myCPU.scala 1187:23]
  assign _dmemreq_io_WriteDataE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 838:23]
  assign _ex2mem_clock = clock;
  assign _ex2mem_reset = reset;
  assign _ex2mem_io1_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_LoadUnsignedE = _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_csrWriteE = _id2ex_io2_csrWriteE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_WritecsrAddrE = _id2ex_io2_WritecsrAddrE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_PCE = _id2ex_io2_PCE; // @[myCPU.scala 163:15]
  assign _ex2mem_io1_BranchJump_JrE = _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 163:15]
  assign _ex2mem_io_en = _cfu_io_StallE; // @[myCPU.scala 210:30]
  assign _ex2mem_io_clr = _cfu_io_FlushM; // @[myCPU.scala 211:30]
  assign _ex2mem_io_WriteDataE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 838:23]
  assign _ex2mem_io_WriteRegE = _id2ex_io2_RegDstE; // @[myCPU.scala 924:26]
  assign _ex2mem_io_PhyAddrE = {{32'd0}, _addr_cal_io_d_paddr}; // @[myCPU.scala 927:27]
  assign _ex2mem_io_CsrWritedataE = _CalCsrDataE_T_12 | _CalCsrDataE_T_11; // @[Mux.scala 27:73]
  assign _ex2mem_io_ExceptionTypeE = _id2ex_io_ExceptionTypeE_Out != 32'h0 ? _id2ex_io_ExceptionTypeE_Out : {{19'd0},
    _temp_exceptionE_T_11}; // @[myCPU.scala 908:30]
  assign _mem2mem2_clock = clock;
  assign _mem2mem2_reset = reset;
  assign _mem2mem2_io1_RegWriteE = _ex2mem_io_RegWriteM; // @[myCPU.scala 1037:30]
  assign _mem2mem2_io1_MemToRegE = _ex2mem_io_MemToRegM; // @[myCPU.scala 1038:30]
  assign _mem2mem2_io1_LoadUnsignedE = _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 1042:30]
  assign _mem2mem2_io1_MemWidthE = _ex2mem_io_MemWidthM; // @[myCPU.scala 1043:30]
  assign _mem2mem2_io1_csrWriteE = _ex2mem_io_csrWriteM; // @[myCPU.scala 1046:54]
  assign _mem2mem2_io1_WritecsrAddrE = inst_tlb_exceptionM ? 12'ha : _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 1047:36]
  assign _mem2mem2_io1_PCE = _ex2mem_io_PCM; // @[myCPU.scala 1048:30]
  assign _mem2mem2_io1_BranchJump_JrE = _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 1051:30]
  assign _mem2mem2_io_en = _cfu_io_StallM2; // @[myCPU.scala 1079:20]
  assign _mem2mem2_io_clr = _cfu_io_FlushM2; // @[myCPU.scala 1078:20]
  assign _mem2mem2_io_WriteDataE = _ex2mem_io_WriteDataM; // @[myCPU.scala 1075:30]
  assign _mem2mem2_io_WriteRegE = _ex2mem_io_WriteRegM; // @[myCPU.scala 1027:24]
  assign _mem2mem2_io_PhyAddrE = _ex2mem_io_PhyAddrM; // @[myCPU.scala 1028:23]
  assign _mem2mem2_io_CsrWritedataE = _ex2mem_io_CsrWritedataM; // @[myCPU.scala 1061:29]
  assign _mem2mem2_io_ExceptionTypeE = mem_exception ? _ex2mem_io_ExceptionTypeM_Out : 32'h0; // @[myCPU.scala 1020:21]
  assign _id2ex_clock = clock;
  assign _id2ex_reset = reset;
  assign _id2ex_io1_RegWriteD = _cu_io_RegWriteD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_MemToRegD = _cu_io_MemToRegD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_MemWriteD = _cu_io_MemWriteD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_ALUCtrlD = _cu_io_ALUCtrlD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_ALUSrcD_0 = _cu_io_ALUSrcD_0; // @[myCPU.scala 162:15]
  assign _id2ex_io1_ALUSrcD_1 = _cu_io_ALUSrcD_1; // @[myCPU.scala 162:15]
  assign _id2ex_io1_RegDstD = _cu_io_RegDstD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_LinkD = _cu_io_LinkD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_csrWriteD = _cu_io_csrWriteD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_csrToRegD = _cu_io_csrToRegD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_LoadUnsignedD = _cu_io_LoadUnsignedD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_MemWidthD = _cu_io_MemWidthD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_data_wD = _cu_io_data_wD; // @[myCPU.scala 162:15]
  assign _id2ex_io1_muldiv_control = _cu_io_muldiv_control; // @[myCPU.scala 162:15]
  assign _id2ex_io1_muldiv_cal = _cu_io_muldiv_cal; // @[myCPU.scala 162:15]
  assign _id2ex_io1_alu_cal = _cu_io_alu_cal; // @[myCPU.scala 162:15]
  assign _id2ex_io1_csr_control = _cu_io_csr_control; // @[myCPU.scala 162:15]
  assign _id2ex_io1_csr_Imm = _cu_io_csr_Imm; // @[myCPU.scala 162:15]
  assign _id2ex_io1_fence_i_control = _cu_io_fence_i_control; // @[myCPU.scala 162:15]
  assign _id2ex_io_en = _cfu_io_StallD; // @[myCPU.scala 191:29]
  assign _id2ex_io_clr = _cfu_io_FlushE; // @[myCPU.scala 192:29]
  assign _id2ex_io_RD1D = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 801:25]
  assign _id2ex_io_RD2D = _cfu_io_Forward2D[0] ? resultE2M_Reg : _BranchR2D_T_2; // @[myCPU.scala 802:25]
  assign _id2ex_io_R2D = _if2id_io_InstrD[24:20]; // @[myCPU.scala 203:27]
  assign _id2ex_io_R1D = _if2id_io_InstrD[19:15]; // @[myCPU.scala 204:27]
  assign _id2ex_io_ImmD = _cu_io_ImmD; // @[myCPU.scala 800:19]
  assign _id2ex_io_PCPlus4D = _if2id_io_PCPlus4D; // @[myCPU.scala 808:29]
  assign _id2ex_io_WritecsrAddrD = _if2id_io_InstrD[31:20]; // @[myCPU.scala 803:38]
  assign _id2ex_io_ReadcsrAddrD = _if2id_io_InstrD[31:20]; // @[myCPU.scala 805:38]
  assign _id2ex_io_PCD = _if2id_io_PCD; // @[myCPU.scala 809:28]
  assign _id2ex_io_ExceptionTypeD = __id2ex_io_ExceptionTypeD_T_6 ? 32'h1 : __id2ex_io_ExceptionTypeD_T_16; // @[myCPU.scala 789:37]
  assign _id2ex_io_BranchJump_JrD = pre_decoder_branchD_flag | pre_decoder_jump; // @[myCPU.scala 811:66]
  assign _if2id_clock = clock;
  assign _if2id_reset = reset;
  assign _if2id_io_en = _cfu_io_StallD; // @[myCPU.scala 598:30]
  assign _if2id_io_clr = _cfu_io_FlushD; // @[myCPU.scala 599:30]
  assign _if2id_io_InstrF = _cu_io1_BadInstrD | _cu_io1_SysCallD | __if2id_io_InstrF_T_3 ? 32'h0 :
    inst_buffer_read_out_inst; // @[myCPU.scala 602:33]
  assign _if2id_io_PCPlus4F = _if2id_io_PCF + 64'h4; // @[myCPU.scala 596:48]
  assign _if2id_io_PCF = {{32'd0}, inst_buffer_read_out_pc}; // @[myCPU.scala 595:30]
  assign _if2id_io_ExceptionTypeF = fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 583:36 584:26]
  assign _mem22wb_clock = clock;
  assign _mem22wb_reset = reset;
  assign _mem22wb_io_en = _cfu_io_StallW; // @[myCPU.scala 282:31]
  assign _mem22wb_io_clr = _cfu_io_FlushW; // @[myCPU.scala 283:31]
  assign _mem22wb_io_RegWriteM = _mem2mem2_io_RegWriteM; // @[myCPU.scala 285:38]
  assign _mem22wb_io_ResultM = _Forward_Lock1E_T_1 ? Mem_withRL_Data : ResultM2_Reg; // @[myCPU.scala 1086:25]
  assign _mem22wb_io_WriteRegM = _mem2mem2_io_WriteRegM; // @[myCPU.scala 287:38]
  assign _mem22wb_io_csrWriteM = _mem2mem2_io_csrWriteM; // @[myCPU.scala 289:38]
  assign _mem22wb_io_WritecsrAddrM = _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 290:38]
  assign _mem22wb_io_CsrWritedataM = _mem2mem2_io_CsrWritedataM; // @[myCPU.scala 1097:33]
  assign _mem22wb_io_PCM = _mem2mem2_io_PCM; // @[myCPU.scala 288:38]
  assign _mem22wb_io_ExceptionTypeM = _mem2mem2_io_ExceptionTypeM_Out[31:1]; // @[myCPU.scala 1092:67]
  assign _mem22wb_io_BranchJump_JrM = _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 1096:33]
  assign _addr_cal_io_d_vaddr = __addr_cal_io_d_vaddr_T_1[31:0]; // @[myCPU.scala 1185:26]
  assign _muldiv_clock = clock;
  assign _muldiv_reset = reset;
  assign _muldiv_io_en = ~ex_exception & ~__muldiv_io_en_T_23; // @[myCPU.scala 877:36]
  assign _muldiv_io_ctrl = _id2ex_io_muldiv_control; // @[myCPU.scala 884:21]
  assign _muldiv_io_in1 = _id2ex_io2_ALUSrcE_0 ? _id2ex_io2_PCE : RD1ForWardE; // @[myCPU.scala 859:20]
  assign _muldiv_io_in2 = _id2ex_io2_ALUSrcE_1 ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 866:20]
  assign _regfile_clock = clock;
  assign _regfile_reset = reset;
  assign _regfile_io_A1 = _if2id_io_InstrD[19:15]; // @[myCPU.scala 747:29]
  assign _regfile_io_A2 = _if2id_io_InstrD[24:20]; // @[myCPU.scala 748:29]
  assign _regfile_io_WE3 = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1149:21]
  assign _regfile_io_A3 = _mem22wb_io_WriteRegW; // @[myCPU.scala 1155:21]
  assign _regfile_io_WD3 = _mem22wb_io_ResultW; // @[myCPU.scala 1148:15 296:26]
  assign fifo_with_bundle_clock = clock;
  assign fifo_with_bundle_reset = reset;
  assign fifo_with_bundle_io_read_en = _cfu_io_StallF; // @[myCPU.scala 558:51]
  assign fifo_with_bundle_io_write_en = inst_write_en[0]; // @[myCPU.scala 550:29]
  assign fifo_with_bundle_io_write_in_0_pc = stage_fec_2_pc_L_io_out_pc_value_out; // @[myCPU.scala 529:40 532:45]
  assign fifo_with_bundle_io_write_in_0_inst = inst_sram_rdata_L[31:0]; // @[myCPU.scala 531:60]
  assign fifo_with_bundle_io_write_in_0_pre_pc_target = stage_fec_2_pre_target_0[31:0]; // @[myCPU.scala 529:40 544:55]
  assign fifo_with_bundle_io_write_in_0_pre_lookup_data = branch_prediction_io_lookup_data; // @[myCPU.scala 480:40 482:32]
  assign fifo_with_bundle_io_write_in_0_pre_hashcode = stage_fec_2_hascode_0; // @[myCPU.scala 529:40 543:55]
  assign fifo_with_bundle_io_write_in_0_pre_pht = branch_prediction_io_out; // @[myCPU.scala 476:32 488:24]
  assign fifo_with_bundle_io_write_in_0_pre_bht = stage_fec_2_bht_0; // @[myCPU.scala 529:40 534:45]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag = inst_sram_rdata_L[32]; // @[myCPU.scala 538:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_jump = inst_sram_rdata_L[33]; // @[myCPU.scala 539:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_branchdata = inst_sram_rdata_L[39:34]; // @[myCPU.scala 541:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_jr = inst_buffer_write_bundle_pre_decoder_jr_opD == 7'h67 &
    inst_buffer_write_bundle_pre_decoder_jr_Funct3D == 3'h0; // @[macros.scala 505:30]
  assign fifo_with_bundle_io_write_in_0_true_branch_state = branch_prediction_io_pre & (stage_fec_2_inst_branch |
    stage_fec_2_inst_jump) & branch_prediction_io_btb_hit & stage_fec_2_stall_reg & stage_fec_2_valid & ~
    _csr_io_exception; // @[myCPU.scala 499:185]
  assign fifo_with_bundle_io_point_write_en = _stage_fec_2_branch_answer_T_8 | _PCSrcD_T_1 & ((pre_decoder_jump |
    _PCSrcD_T_3) != id_true_branch_state | target_addr_error) & ~(ex_exception | mem_exception | mem2_exception |
    wb_exception); // @[myCPU.scala 710:60]
  assign fifo_with_bundle_io_point_flush = _csr_io_exception; // @[myCPU.scala 559:29]
  assign stage_fec_1_pc_L_clock = clock;
  assign stage_fec_1_pc_L_reset = reset;
  assign stage_fec_1_pc_L_io_stall = stage2_stall; // @[myCPU.scala 439:31]
  assign stage_fec_1_pc_L_io_flush = _stage_fec_2_branch_answer_T_8 & ~stage2_stall; // @[myCPU.scala 404:54]
  assign stage_fec_1_pc_L_io_in_pc_value_in = inst_sram_addr[31:0]; // @[myCPU.scala 430:40]
  assign branch_prediction_clock = clock;
  assign branch_prediction_reset = reset;
  assign branch_prediction_io_pc = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 448:12]
  assign branch_prediction_io_write_pc = _mem22wb_io_PCW[31:0]; // @[myCPU.scala 1173:17]
  assign branch_prediction_io_aw_pht_ways_addr = wb_bru_state_io_out_hashcode; // @[myCPU.scala 1172:25]
  assign branch_prediction_io_aw_pht_addr = wb_bru_state_io_out_lookup_data; // @[myCPU.scala 1170:20]
  assign branch_prediction_io_aw_bht_addr = _mem22wb_io_PCW[10:4]; // @[myCPU.scala 1169:38]
  assign branch_prediction_io_aw_target_addr = wb_bru_state_io_out_target_pc[31:0]; // @[myCPU.scala 1171:23]
  assign branch_prediction_io_btb_write = branch_prediction_io_bht_write; // @[myCPU.scala 1168:18]
  assign branch_prediction_io_bht_write = _mem22wb_io_BranchJump_JrW; // @[myCPU.scala 1166:47]
  assign branch_prediction_io_pht_write = branch_prediction_io_bht_write; // @[myCPU.scala 1167:18]
  assign branch_prediction_io_bht_in = wb_bru_state_io_out_bht; // @[myCPU.scala 1164:15]
  assign branch_prediction_io_pht_in = wb_bru_state_io_out_pht; // @[myCPU.scala 1165:15]
  assign branch_prediction_io_stage2_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 465:42]
  assign branch_prediction_io_stage2_flush = stage2_flush; // @[myCPU.scala 468:22]
  assign stage_fec_2_pc_L_clock = clock;
  assign stage_fec_2_pc_L_reset = reset;
  assign stage_fec_2_pc_L_io_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 465:42]
  assign stage_fec_2_pc_L_io_flush = stage2_flush; // @[myCPU.scala 523:31]
  assign stage_fec_2_pc_L_io_in_pc_value_in = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 519:40]
  assign id_bru_state_clock = clock;
  assign id_bru_state_reset = reset;
  assign id_bru_state_io_stall = _cfu_io_StallD; // @[myCPU.scala 668:27]
  assign id_bru_state_io_flush = _cfu_io_FlushD; // @[myCPU.scala 667:27]
  assign id_bru_state_io_in_pht = fifo_with_bundle_io_read_out_0_pre_pht; // @[myCPU.scala 583:36 584:26]
  assign id_bru_state_io_in_bht = fifo_with_bundle_io_read_out_0_pre_bht; // @[myCPU.scala 583:36 584:26]
  assign id_bru_state_io_in_hashcode = fifo_with_bundle_io_read_out_0_pre_hashcode; // @[myCPU.scala 583:36 584:26]
  assign id_bru_state_io_in_target_pc = {{32'd0}, inst_buffer_read_out_pre_pc_target}; // @[myCPU.scala 698:34]
  assign id_bru_state_io_in_lookup_data = fifo_with_bundle_io_read_out_0_pre_lookup_data; // @[myCPU.scala 583:36 584:26]
  assign ex_bru_state_clock = clock;
  assign ex_bru_state_reset = reset;
  assign ex_bru_state_io_stall = _cfu_io_StallE; // @[myCPU.scala 672:27]
  assign ex_bru_state_io_flush = _cfu_io_FlushE; // @[myCPU.scala 671:27]
  assign ex_bru_state_io_in_pht = id_bru_state_io_out_pht; // @[myCPU.scala 727:28]
  assign ex_bru_state_io_in_bht = id_bru_state_io_out_bht; // @[myCPU.scala 726:28]
  assign ex_bru_state_io_in_hashcode = id_bru_state_io_out_hashcode; // @[myCPU.scala 728:33]
  assign ex_bru_state_io_in_target_pc = pre_decoder_branchD_flag ? PCBranchD : _Pc_targetD_T_2; // @[Mux.scala 101:16]
  assign ex_bru_state_io_in_lookup_data = id_bru_state_io_out_lookup_data; // @[myCPU.scala 729:36]
  assign mem_bru_state_clock = clock;
  assign mem_bru_state_reset = reset;
  assign mem_bru_state_io_stall = _cfu_io_StallM; // @[myCPU.scala 676:28]
  assign mem_bru_state_io_flush = _cfu_io_FlushM; // @[myCPU.scala 675:28]
  assign mem_bru_state_io_in_pht = 2'h2 == ex_bru_state_io_out_pht ? _pht_tobeE_T_3 : _pht_tobeE_T_7; // @[Mux.scala 81:58]
  assign mem_bru_state_io_in_bht = {ex_bru_state_io_out_bht[5:0],true_branch_stateE}; // @[Cat.scala 31:58]
  assign mem_bru_state_io_in_hashcode = ex_bru_state_io_out_hashcode; // @[myCPU.scala 687:26]
  assign mem_bru_state_io_in_target_pc = ex_bru_state_io_out_target_pc; // @[myCPU.scala 687:26]
  assign mem_bru_state_io_in_lookup_data = ex_bru_state_io_out_lookup_data; // @[myCPU.scala 687:26]
  assign mem2_bru_state_clock = clock;
  assign mem2_bru_state_reset = reset;
  assign mem2_bru_state_io_stall = _cfu_io_StallM2; // @[myCPU.scala 680:29]
  assign mem2_bru_state_io_flush = _cfu_io_FlushM2; // @[myCPU.scala 679:29]
  assign mem2_bru_state_io_in_pht = mem_bru_state_io_out_pht; // @[myCPU.scala 688:26]
  assign mem2_bru_state_io_in_bht = mem_bru_state_io_out_bht; // @[myCPU.scala 688:26]
  assign mem2_bru_state_io_in_hashcode = mem_bru_state_io_out_hashcode; // @[myCPU.scala 688:26]
  assign mem2_bru_state_io_in_target_pc = mem_bru_state_io_out_target_pc; // @[myCPU.scala 688:26]
  assign mem2_bru_state_io_in_lookup_data = mem_bru_state_io_out_lookup_data; // @[myCPU.scala 688:26]
  assign wb_bru_state_clock = clock;
  assign wb_bru_state_reset = reset;
  assign wb_bru_state_io_stall = _cfu_io_StallW; // @[myCPU.scala 684:27]
  assign wb_bru_state_io_flush = _cfu_io_FlushW; // @[myCPU.scala 683:27]
  assign wb_bru_state_io_in_pht = mem2_bru_state_io_out_pht; // @[myCPU.scala 689:26]
  assign wb_bru_state_io_in_bht = mem2_bru_state_io_out_bht; // @[myCPU.scala 689:26]
  assign wb_bru_state_io_in_hashcode = mem2_bru_state_io_out_hashcode; // @[myCPU.scala 689:26]
  assign wb_bru_state_io_in_target_pc = mem2_bru_state_io_out_target_pc; // @[myCPU.scala 689:26]
  assign wb_bru_state_io_in_lookup_data = mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 689:26]
  always @(posedge clock) begin
    if (reset) begin // @[myCPU.scala 180:44]
      pre_decoder_branchD_flag <= 1'h0; // @[myCPU.scala 180:44]
    end else if (_cfu_io_FlushD) begin // @[myCPU.scala 587:36]
      pre_decoder_branchD_flag <= 1'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 587:66]
      pre_decoder_branchD_flag <= inst_buffer_read_out_pre_decoder_branchD_flag;
    end
    if (reset) begin // @[myCPU.scala 181:43]
      pre_decoder_branchdata <= 6'h0; // @[myCPU.scala 181:43]
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 589:34]
      pre_decoder_branchdata <= 6'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 589:64]
      pre_decoder_branchdata <= inst_buffer_read_out_pre_decoder_branchdata;
    end
    if (reset) begin // @[myCPU.scala 182:40]
      pre_decoder_jump <= 1'h0; // @[myCPU.scala 182:40]
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 588:28]
      pre_decoder_jump <= 1'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 588:58]
      pre_decoder_jump <= inst_buffer_read_out_pre_decoder_jump;
    end
    if (reset) begin // @[myCPU.scala 183:40]
      pre_decoder_jr <= 1'h0; // @[myCPU.scala 183:40]
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 590:26]
      pre_decoder_jr <= 1'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 590:56]
      pre_decoder_jr <= inst_buffer_read_out_pre_decoder_jr;
    end
    if (reset) begin // @[myCPU.scala 963:32]
      resultE2M_Reg <= 64'h0; // @[myCPU.scala 963:32]
    end else if (_mem_exception_T) begin // @[myCPU.scala 968:25]
      resultE2M_Reg <= 64'h0;
    end else if (_mem_exception_T_1) begin // @[myCPU.scala 968:55]
      resultE2M_Reg <= resultE;
    end
    if (reset) begin // @[myCPU.scala 1016:29]
      ResultM2_Reg <= 64'h0; // @[myCPU.scala 1016:29]
    end else if (_mem2_exception_T) begin // @[myCPU.scala 1018:24]
      ResultM2_Reg <= 64'h0;
    end else if (_mem2_exception_T_1) begin // @[myCPU.scala 1018:55]
      ResultM2_Reg <= resultE2M_Reg;
    end
    if (reset) begin // @[myCPU.scala 264:34]
      fence_i_controlMReg <= 1'h0; // @[myCPU.scala 264:34]
    end else if (_ex2mem_io_clr) begin // @[myCPU.scala 265:27]
      fence_i_controlMReg <= 1'h0;
    end else if (_ex2mem_io_en) begin // @[myCPU.scala 266:12]
      fence_i_controlMReg <= _id2ex_io_fence_i_controlE;
    end
    if (reset) begin // @[myCPU.scala 299:26]
      PCW_Reg <= 64'h0; // @[myCPU.scala 299:26]
    end else if (_mem22wb_io_PCW != 64'h0) begin // @[myCPU.scala 303:19]
      PCW_Reg <= _mem22wb_io_PCW;
    end
    if (reset) begin // @[myCPU.scala 344:33]
      pc_next_wait <= 64'h0; // @[myCPU.scala 344:33]
    end else if (ready_to_branch | stage_fec_2_branch_answer) begin // @[myCPU.scala 347:24]
      if (fifo_with_bundle_io_point_write_en) begin // @[myCPU.scala 743:26]
        if (pre_decoder_jump) begin // @[Mux.scala 101:16]
          pc_next_wait <= PCJumpD;
        end else begin
          pc_next_wait <= _PC_nextD_T_2;
        end
      end else if (stage_fec_2_branch_answer) begin // @[myCPU.scala 418:31]
        pc_next_wait <= stage_fec_2_pre_target_0;
      end else begin
        pc_next_wait <= _stage_fec_1_pc_next_T_1;
      end
    end
    if (reset) begin // @[myCPU.scala 496:40]
      stage_fec_2_stall_reg <= 1'h0; // @[myCPU.scala 496:40]
    end else begin
      stage_fec_2_stall_reg <= stage_fec_2_stall; // @[myCPU.scala 497:27]
    end
    if (reset) begin // @[myCPU.scala 472:36]
      stage_fec_2_valid <= 1'h0; // @[myCPU.scala 472:36]
    end else if (stage_fec_2_stall) begin // @[myCPU.scala 473:29]
      if (fifo_with_bundle_io_point_write_en) begin // @[myCPU.scala 473:51]
        stage_fec_2_valid <= 1'h0;
      end else begin
        stage_fec_2_valid <= stage_fec_1_valid;
      end
    end
    if (reset) begin // @[myCPU.scala 348:30]
      pc_req_wait <= 1'h0; // @[myCPU.scala 348:30]
    end else begin
      pc_req_wait <= _GEN_1;
    end
    if (reset) begin // @[myCPU.scala 361:35]
      exception_Pc_reg <= 64'h0; // @[myCPU.scala 361:35]
    end else if (_stage_fec_2_branch_answer_T_8) begin // @[myCPU.scala 362:28]
      exception_Pc_reg <= _csr_io_return_pc;
    end
    if (reset) begin // @[myCPU.scala 364:36]
      returnPc_req_wait <= 1'h0; // @[myCPU.scala 364:36]
    end else begin
      returnPc_req_wait <= _GEN_3;
    end
    if (reset) begin // @[myCPU.scala 451:36]
      stage_fec_1_valid <= 1'h0; // @[myCPU.scala 451:36]
    end else begin
      stage_fec_1_valid <= stage2_stall | _stage_fec_1_valid_T_2; // @[myCPU.scala 455:23]
    end
    if (reset) begin // @[myCPU.scala 475:35]
      stage_fec_2_bht_0 <= 7'h0; // @[myCPU.scala 475:35]
    end else if (stage2_flush) begin // @[myCPU.scala 485:30]
      stage_fec_2_bht_0 <= 7'h0;
    end else if (stage2_stall) begin // @[myCPU.scala 485:51]
      stage_fec_2_bht_0 <= branch_prediction_io_bht;
    end
    if (reset) begin // @[myCPU.scala 479:39]
      stage_fec_2_hascode_0 <= 4'h0; // @[myCPU.scala 479:39]
    end else if (stage2_flush) begin // @[myCPU.scala 493:36]
      stage_fec_2_hascode_0 <= 4'h0;
    end else if (stage2_stall) begin // @[myCPU.scala 493:57]
      stage_fec_2_hascode_0 <= _stage_fec_2_hascode_0_T_1;
    end
    if (reset) begin // @[myCPU.scala 606:31]
      id_exception <= 1'h0; // @[myCPU.scala 606:31]
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 607:24]
      id_exception <= 1'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 607:54]
      id_exception <= _if2id_io_PCF[1:0] != 2'h0 | inst_buffer_read_out_exception_type != 2'h0;
    end
    if (reset) begin // @[myCPU.scala 609:31]
      ex_exception <= 1'h0; // @[myCPU.scala 609:31]
    end else if (_cfu_io_FlushE) begin // @[myCPU.scala 610:24]
      ex_exception <= 1'h0;
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 610:54]
      ex_exception <= _id2ex_io_ExceptionTypeD != 32'h0;
    end
    if (reset) begin // @[myCPU.scala 612:32]
      mem_exception <= 1'h0; // @[myCPU.scala 612:32]
    end else if (_cfu_io_FlushM) begin // @[myCPU.scala 613:25]
      mem_exception <= 1'h0;
    end else if (_cfu_io_StallM) begin // @[myCPU.scala 613:55]
      mem_exception <= _ex2mem_io_ExceptionTypeE != 32'h0;
    end
    if (reset) begin // @[myCPU.scala 615:33]
      mem2_exception <= 1'h0; // @[myCPU.scala 615:33]
    end else if (_cfu_io_FlushM2) begin // @[myCPU.scala 616:26]
      mem2_exception <= 1'h0;
    end else if (_cfu_io_StallM2) begin // @[myCPU.scala 616:57]
      mem2_exception <= _mem2mem2_io_ExceptionTypeE != 32'h0;
    end
    if (reset) begin // @[myCPU.scala 618:31]
      wb_exception <= 1'h0; // @[myCPU.scala 618:31]
    end else if (_cfu_io_FlushW) begin // @[myCPU.scala 619:24]
      wb_exception <= 1'h0;
    end else if (_cfu_io_StallW) begin // @[myCPU.scala 619:54]
      wb_exception <= mem2_exception;
    end
    if (reset) begin // @[myCPU.scala 663:39]
      id_true_branch_state <= 1'h0; // @[myCPU.scala 663:39]
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 664:32]
      id_true_branch_state <= 1'h0;
    end else if (_PCSrcD_T_1) begin // @[myCPU.scala 664:62]
      id_true_branch_state <= inst_buffer_read_out_true_branch_state;
    end
    if (reset) begin // @[myCPU.scala 693:38]
      inst_tlb_exceptionE <= 1'h0; // @[myCPU.scala 693:38]
    end else if (_ex_exception_T) begin // @[myCPU.scala 694:31]
      inst_tlb_exceptionE <= 1'h0;
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 694:61]
      inst_tlb_exceptionE <= _if2id_io_ExceptionTypeD_Out != 2'h0;
    end
    if (reset) begin // @[myCPU.scala 721:37]
      true_branch_stateE <= 1'h0; // @[myCPU.scala 721:37]
    end else if (_ex_exception_T) begin // @[myCPU.scala 723:30]
      true_branch_stateE <= 1'h0;
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 723:61]
      true_branch_stateE <= _T_28;
    end
    if (reset) begin // @[myCPU.scala 764:33]
      int_instanceE_timer <= 1'h0; // @[myCPU.scala 764:33]
    end else if (_ex_exception_T) begin // @[myCPU.scala 780:25]
      int_instanceE_timer <= 1'h0;
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 780:82]
      int_instanceE_timer <= ext_int_with_enable_timer;
    end
    if (reset) begin // @[myCPU.scala 764:33]
      int_instanceE_out_int <= 1'h0; // @[myCPU.scala 764:33]
    end else if (_ex_exception_T) begin // @[myCPU.scala 780:25]
      int_instanceE_out_int <= 1'h0;
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 780:82]
      int_instanceE_out_int <= ext_int_with_enable_out_int;
    end
    if (reset) begin // @[myCPU.scala 765:33]
      int_instanceM_timer <= 1'h0; // @[myCPU.scala 765:33]
    end else if (_mem_exception_T) begin // @[myCPU.scala 781:25]
      int_instanceM_timer <= 1'h0;
    end else if (_mem_exception_T_1) begin // @[myCPU.scala 781:82]
      int_instanceM_timer <= int_instanceE_timer;
    end
    if (reset) begin // @[myCPU.scala 765:33]
      int_instanceM_out_int <= 1'h0; // @[myCPU.scala 765:33]
    end else if (_mem_exception_T) begin // @[myCPU.scala 781:25]
      int_instanceM_out_int <= 1'h0;
    end else if (_mem_exception_T_1) begin // @[myCPU.scala 781:82]
      int_instanceM_out_int <= int_instanceE_out_int;
    end
    if (reset) begin // @[myCPU.scala 766:33]
      int_instanceM2_timer <= 1'h0; // @[myCPU.scala 766:33]
    end else if (_mem2_exception_T) begin // @[myCPU.scala 782:26]
      int_instanceM2_timer <= 1'h0;
    end else if (_mem2_exception_T_1) begin // @[myCPU.scala 782:82]
      int_instanceM2_timer <= int_instanceM_timer;
    end
    if (reset) begin // @[myCPU.scala 766:33]
      int_instanceM2_out_int <= 1'h0; // @[myCPU.scala 766:33]
    end else if (_mem2_exception_T) begin // @[myCPU.scala 782:26]
      int_instanceM2_out_int <= 1'h0;
    end else if (_mem2_exception_T_1) begin // @[myCPU.scala 782:82]
      int_instanceM2_out_int <= int_instanceM_out_int;
    end
    if (reset) begin // @[myCPU.scala 767:33]
      int_instanceW_timer <= 1'h0; // @[myCPU.scala 767:33]
    end else if (_wb_exception_T) begin // @[myCPU.scala 783:25]
      int_instanceW_timer <= 1'h0;
    end else if (_wb_exception_T_1) begin // @[myCPU.scala 783:82]
      int_instanceW_timer <= int_instanceM2_timer;
    end
    if (reset) begin // @[myCPU.scala 767:33]
      int_instanceW_out_int <= 1'h0; // @[myCPU.scala 767:33]
    end else if (_wb_exception_T) begin // @[myCPU.scala 783:25]
      int_instanceW_out_int <= 1'h0;
    end else if (_wb_exception_T_1) begin // @[myCPU.scala 783:82]
      int_instanceW_out_int <= int_instanceM2_out_int;
    end
    if (reset) begin // @[myCPU.scala 831:34]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 831:34]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 839:33]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 840:24]
    end else if ((_cfu_io_Forward1E[0] | _cfu_io_Forward1E[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 843:88]
      Forward_Lock1E <= ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM); // @[myCPU.scala 844:28]
    end
    if (reset) begin // @[myCPU.scala 829:34]
      RD1ForWardE_r <= 64'h0; // @[myCPU.scala 829:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 839:33]
      if ((_cfu_io_Forward1E[0] | _cfu_io_Forward1E[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 843:88]
        if (2'h3 == _cfu_io_Forward1E) begin // @[Mux.scala 81:58]
          RD1ForWardE_r <= ResultM2_Reg;
        end else begin
          RD1ForWardE_r <= _RD1ForWardE_p_T_3;
        end
      end
    end
    if (reset) begin // @[myCPU.scala 824:34]
      inst_tlb_exceptionM <= 1'h0; // @[myCPU.scala 824:34]
    end else if (_mem_exception_T) begin // @[myCPU.scala 825:27]
      inst_tlb_exceptionM <= 1'h0;
    end else if (_mem_exception_T_1) begin // @[myCPU.scala 825:57]
      inst_tlb_exceptionM <= inst_tlb_exceptionE;
    end
    if (reset) begin // @[myCPU.scala 830:34]
      RD2ForWardE_r <= 64'h0; // @[myCPU.scala 830:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 839:33]
      if ((_cfu_io_Forward2E[0] | _cfu_io_Forward2E[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 847:87]
        if (2'h3 == _cfu_io_Forward2E) begin // @[Mux.scala 81:58]
          RD2ForWardE_r <= ResultM2_Reg;
        end else begin
          RD2ForWardE_r <= _RD2ForWardE_p_T_3;
        end
      end
    end
    if (reset) begin // @[myCPU.scala 832:34]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 832:34]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 839:33]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 841:24]
    end else if ((_cfu_io_Forward2E[0] | _cfu_io_Forward2E[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 847:87]
      Forward_Lock2E <= _Forward_Lock1E_T_3; // @[myCPU.scala 848:28]
    end
    if (reset) begin // @[myCPU.scala 1063:40]
      tlb_exception_csr_writeM2 <= 1'h0; // @[myCPU.scala 1063:40]
    end else if (_mem2_exception_T) begin // @[myCPU.scala 1065:33]
      tlb_exception_csr_writeM2 <= 1'h0;
    end else if (_mem2_exception_T_1) begin // @[myCPU.scala 1065:64]
      tlb_exception_csr_writeM2 <= inst_tlb_exceptionM;
    end
    if (reset) begin // @[myCPU.scala 1064:40]
      tlb_exception_co0_writeW <= 1'h0; // @[myCPU.scala 1064:40]
    end else if (_wb_exception_T) begin // @[myCPU.scala 1066:33]
      tlb_exception_co0_writeW <= 1'h0;
    end else if (_wb_exception_T_1) begin // @[myCPU.scala 1066:63]
      tlb_exception_co0_writeW <= tlb_exception_csr_writeM2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_decoder_branchD_flag = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pre_decoder_branchdata = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  pre_decoder_jump = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pre_decoder_jr = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  resultE2M_Reg = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ResultM2_Reg = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  fence_i_controlMReg = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  PCW_Reg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  pc_next_wait = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  stage_fec_2_stall_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  stage_fec_2_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pc_req_wait = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  exception_Pc_reg = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  returnPc_req_wait = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  stage_fec_1_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  stage_fec_2_bht_0 = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  stage_fec_2_hascode_0 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  id_exception = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ex_exception = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  mem_exception = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mem2_exception = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  wb_exception = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  id_true_branch_state = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inst_tlb_exceptionE = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  true_branch_stateE = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  int_instanceE_timer = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  int_instanceE_out_int = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  int_instanceM_timer = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  int_instanceM_out_int = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  int_instanceM2_timer = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  int_instanceM2_out_int = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  int_instanceW_timer = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  int_instanceW_out_int = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  Forward_Lock1E = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  RD1ForWardE_r = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  inst_tlb_exceptionM = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  RD2ForWardE_r = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  Forward_Lock2E = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tlb_exception_csr_writeM2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tlb_exception_co0_writeW = _RAND_39[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_icache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [21:0] io_wdata,
  input  [31:0] io_addr,
  output        io_hit,
  output        io_valid,
  input         io_tag_all_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] tag_regs_0; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_1; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_2; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_3; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_4; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_5; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_6; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_7; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_8; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_9; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_10; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_11; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_12; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_13; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_14; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_15; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_16; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_17; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_18; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_19; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_20; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_21; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_22; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_23; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_24; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_25; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_26; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_27; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_28; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_29; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_30; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_31; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_32; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_33; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_34; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_35; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_36; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_37; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_38; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_39; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_40; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_41; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_42; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_43; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_44; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_45; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_46; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_47; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_48; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_49; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_50; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_51; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_52; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_53; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_54; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_55; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_56; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_57; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_58; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_59; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_60; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_61; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_62; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_63; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_64; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_65; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_66; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_67; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_68; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_69; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_70; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_71; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_72; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_73; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_74; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_75; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_76; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_77; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_78; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_79; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_80; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_81; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_82; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_83; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_84; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_85; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_86; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_87; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_88; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_89; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_90; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_91; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_92; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_93; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_94; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_95; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_96; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_97; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_98; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_99; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_100; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_101; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_102; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_103; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_104; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_105; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_106; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_107; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_108; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_109; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_110; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_111; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_112; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_113; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_114; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_115; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_116; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_117; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_118; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_119; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_120; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_121; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_122; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_123; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_124; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_125; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_126; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_127; // @[icache_tag.scala 21:27]
  wire  _valid_to_be_T_5 = io_wen & io_addr[10:4] == 7'h0; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_8 = io_wen & io_addr[10:4] == 7'h0 ? io_wdata[21] : tag_regs_0[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be = io_tag_all_flush ? 1'h0 : _valid_to_be_T_8; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be = _valid_to_be_T_5 ? io_wdata[20:0] : tag_regs_0[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_0_T = {valid_to_be,tag_to_be}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_14 = io_wen & io_addr[10:4] == 7'h1; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_17 = io_wen & io_addr[10:4] == 7'h1 ? io_wdata[21] : tag_regs_1[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_1 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_17; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_1 = _valid_to_be_T_14 ? io_wdata[20:0] : tag_regs_1[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_1_T = {valid_to_be_1,tag_to_be_1}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_23 = io_wen & io_addr[10:4] == 7'h2; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_26 = io_wen & io_addr[10:4] == 7'h2 ? io_wdata[21] : tag_regs_2[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_2 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_26; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_2 = _valid_to_be_T_23 ? io_wdata[20:0] : tag_regs_2[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_2_T = {valid_to_be_2,tag_to_be_2}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_32 = io_wen & io_addr[10:4] == 7'h3; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_35 = io_wen & io_addr[10:4] == 7'h3 ? io_wdata[21] : tag_regs_3[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_3 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_35; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_3 = _valid_to_be_T_32 ? io_wdata[20:0] : tag_regs_3[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_3_T = {valid_to_be_3,tag_to_be_3}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_41 = io_wen & io_addr[10:4] == 7'h4; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_44 = io_wen & io_addr[10:4] == 7'h4 ? io_wdata[21] : tag_regs_4[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_4 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_44; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_4 = _valid_to_be_T_41 ? io_wdata[20:0] : tag_regs_4[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_4_T = {valid_to_be_4,tag_to_be_4}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_50 = io_wen & io_addr[10:4] == 7'h5; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_53 = io_wen & io_addr[10:4] == 7'h5 ? io_wdata[21] : tag_regs_5[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_5 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_53; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_5 = _valid_to_be_T_50 ? io_wdata[20:0] : tag_regs_5[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_5_T = {valid_to_be_5,tag_to_be_5}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_59 = io_wen & io_addr[10:4] == 7'h6; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_62 = io_wen & io_addr[10:4] == 7'h6 ? io_wdata[21] : tag_regs_6[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_6 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_62; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_6 = _valid_to_be_T_59 ? io_wdata[20:0] : tag_regs_6[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_6_T = {valid_to_be_6,tag_to_be_6}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_68 = io_wen & io_addr[10:4] == 7'h7; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_71 = io_wen & io_addr[10:4] == 7'h7 ? io_wdata[21] : tag_regs_7[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_7 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_71; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_7 = _valid_to_be_T_68 ? io_wdata[20:0] : tag_regs_7[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_7_T = {valid_to_be_7,tag_to_be_7}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_77 = io_wen & io_addr[10:4] == 7'h8; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_80 = io_wen & io_addr[10:4] == 7'h8 ? io_wdata[21] : tag_regs_8[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_8 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_80; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_8 = _valid_to_be_T_77 ? io_wdata[20:0] : tag_regs_8[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_8_T = {valid_to_be_8,tag_to_be_8}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_86 = io_wen & io_addr[10:4] == 7'h9; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_89 = io_wen & io_addr[10:4] == 7'h9 ? io_wdata[21] : tag_regs_9[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_9 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_89; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_9 = _valid_to_be_T_86 ? io_wdata[20:0] : tag_regs_9[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_9_T = {valid_to_be_9,tag_to_be_9}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_95 = io_wen & io_addr[10:4] == 7'ha; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_98 = io_wen & io_addr[10:4] == 7'ha ? io_wdata[21] : tag_regs_10[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_10 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_98; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_10 = _valid_to_be_T_95 ? io_wdata[20:0] : tag_regs_10[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_10_T = {valid_to_be_10,tag_to_be_10}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_104 = io_wen & io_addr[10:4] == 7'hb; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_107 = io_wen & io_addr[10:4] == 7'hb ? io_wdata[21] : tag_regs_11[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_11 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_107; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_11 = _valid_to_be_T_104 ? io_wdata[20:0] : tag_regs_11[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_11_T = {valid_to_be_11,tag_to_be_11}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_113 = io_wen & io_addr[10:4] == 7'hc; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_116 = io_wen & io_addr[10:4] == 7'hc ? io_wdata[21] : tag_regs_12[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_12 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_116; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_12 = _valid_to_be_T_113 ? io_wdata[20:0] : tag_regs_12[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_12_T = {valid_to_be_12,tag_to_be_12}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_122 = io_wen & io_addr[10:4] == 7'hd; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_125 = io_wen & io_addr[10:4] == 7'hd ? io_wdata[21] : tag_regs_13[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_13 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_125; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_13 = _valid_to_be_T_122 ? io_wdata[20:0] : tag_regs_13[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_13_T = {valid_to_be_13,tag_to_be_13}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_131 = io_wen & io_addr[10:4] == 7'he; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_134 = io_wen & io_addr[10:4] == 7'he ? io_wdata[21] : tag_regs_14[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_14 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_134; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_14 = _valid_to_be_T_131 ? io_wdata[20:0] : tag_regs_14[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_14_T = {valid_to_be_14,tag_to_be_14}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_140 = io_wen & io_addr[10:4] == 7'hf; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_143 = io_wen & io_addr[10:4] == 7'hf ? io_wdata[21] : tag_regs_15[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_15 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_143; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_15 = _valid_to_be_T_140 ? io_wdata[20:0] : tag_regs_15[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_15_T = {valid_to_be_15,tag_to_be_15}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_149 = io_wen & io_addr[10:4] == 7'h10; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_152 = io_wen & io_addr[10:4] == 7'h10 ? io_wdata[21] : tag_regs_16[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_16 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_152; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_16 = _valid_to_be_T_149 ? io_wdata[20:0] : tag_regs_16[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_16_T = {valid_to_be_16,tag_to_be_16}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_158 = io_wen & io_addr[10:4] == 7'h11; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_161 = io_wen & io_addr[10:4] == 7'h11 ? io_wdata[21] : tag_regs_17[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_17 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_161; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_17 = _valid_to_be_T_158 ? io_wdata[20:0] : tag_regs_17[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_17_T = {valid_to_be_17,tag_to_be_17}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_167 = io_wen & io_addr[10:4] == 7'h12; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_170 = io_wen & io_addr[10:4] == 7'h12 ? io_wdata[21] : tag_regs_18[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_18 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_170; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_18 = _valid_to_be_T_167 ? io_wdata[20:0] : tag_regs_18[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_18_T = {valid_to_be_18,tag_to_be_18}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_176 = io_wen & io_addr[10:4] == 7'h13; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_179 = io_wen & io_addr[10:4] == 7'h13 ? io_wdata[21] : tag_regs_19[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_19 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_179; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_19 = _valid_to_be_T_176 ? io_wdata[20:0] : tag_regs_19[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_19_T = {valid_to_be_19,tag_to_be_19}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_185 = io_wen & io_addr[10:4] == 7'h14; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_188 = io_wen & io_addr[10:4] == 7'h14 ? io_wdata[21] : tag_regs_20[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_20 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_188; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_20 = _valid_to_be_T_185 ? io_wdata[20:0] : tag_regs_20[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_20_T = {valid_to_be_20,tag_to_be_20}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_194 = io_wen & io_addr[10:4] == 7'h15; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_197 = io_wen & io_addr[10:4] == 7'h15 ? io_wdata[21] : tag_regs_21[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_21 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_197; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_21 = _valid_to_be_T_194 ? io_wdata[20:0] : tag_regs_21[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_21_T = {valid_to_be_21,tag_to_be_21}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_203 = io_wen & io_addr[10:4] == 7'h16; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_206 = io_wen & io_addr[10:4] == 7'h16 ? io_wdata[21] : tag_regs_22[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_22 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_206; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_22 = _valid_to_be_T_203 ? io_wdata[20:0] : tag_regs_22[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_22_T = {valid_to_be_22,tag_to_be_22}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_212 = io_wen & io_addr[10:4] == 7'h17; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_215 = io_wen & io_addr[10:4] == 7'h17 ? io_wdata[21] : tag_regs_23[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_23 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_215; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_23 = _valid_to_be_T_212 ? io_wdata[20:0] : tag_regs_23[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_23_T = {valid_to_be_23,tag_to_be_23}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_221 = io_wen & io_addr[10:4] == 7'h18; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_224 = io_wen & io_addr[10:4] == 7'h18 ? io_wdata[21] : tag_regs_24[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_24 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_224; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_24 = _valid_to_be_T_221 ? io_wdata[20:0] : tag_regs_24[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_24_T = {valid_to_be_24,tag_to_be_24}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_230 = io_wen & io_addr[10:4] == 7'h19; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_233 = io_wen & io_addr[10:4] == 7'h19 ? io_wdata[21] : tag_regs_25[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_25 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_233; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_25 = _valid_to_be_T_230 ? io_wdata[20:0] : tag_regs_25[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_25_T = {valid_to_be_25,tag_to_be_25}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_239 = io_wen & io_addr[10:4] == 7'h1a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_242 = io_wen & io_addr[10:4] == 7'h1a ? io_wdata[21] : tag_regs_26[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_26 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_242; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_26 = _valid_to_be_T_239 ? io_wdata[20:0] : tag_regs_26[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_26_T = {valid_to_be_26,tag_to_be_26}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_248 = io_wen & io_addr[10:4] == 7'h1b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_251 = io_wen & io_addr[10:4] == 7'h1b ? io_wdata[21] : tag_regs_27[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_27 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_251; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_27 = _valid_to_be_T_248 ? io_wdata[20:0] : tag_regs_27[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_27_T = {valid_to_be_27,tag_to_be_27}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_257 = io_wen & io_addr[10:4] == 7'h1c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_260 = io_wen & io_addr[10:4] == 7'h1c ? io_wdata[21] : tag_regs_28[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_28 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_260; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_28 = _valid_to_be_T_257 ? io_wdata[20:0] : tag_regs_28[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_28_T = {valid_to_be_28,tag_to_be_28}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_266 = io_wen & io_addr[10:4] == 7'h1d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_269 = io_wen & io_addr[10:4] == 7'h1d ? io_wdata[21] : tag_regs_29[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_29 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_269; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_29 = _valid_to_be_T_266 ? io_wdata[20:0] : tag_regs_29[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_29_T = {valid_to_be_29,tag_to_be_29}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_275 = io_wen & io_addr[10:4] == 7'h1e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_278 = io_wen & io_addr[10:4] == 7'h1e ? io_wdata[21] : tag_regs_30[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_30 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_278; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_30 = _valid_to_be_T_275 ? io_wdata[20:0] : tag_regs_30[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_30_T = {valid_to_be_30,tag_to_be_30}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_284 = io_wen & io_addr[10:4] == 7'h1f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_287 = io_wen & io_addr[10:4] == 7'h1f ? io_wdata[21] : tag_regs_31[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_31 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_287; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_31 = _valid_to_be_T_284 ? io_wdata[20:0] : tag_regs_31[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_31_T = {valid_to_be_31,tag_to_be_31}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_293 = io_wen & io_addr[10:4] == 7'h20; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_296 = io_wen & io_addr[10:4] == 7'h20 ? io_wdata[21] : tag_regs_32[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_32 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_296; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_32 = _valid_to_be_T_293 ? io_wdata[20:0] : tag_regs_32[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_32_T = {valid_to_be_32,tag_to_be_32}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_302 = io_wen & io_addr[10:4] == 7'h21; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_305 = io_wen & io_addr[10:4] == 7'h21 ? io_wdata[21] : tag_regs_33[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_33 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_305; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_33 = _valid_to_be_T_302 ? io_wdata[20:0] : tag_regs_33[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_33_T = {valid_to_be_33,tag_to_be_33}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_311 = io_wen & io_addr[10:4] == 7'h22; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_314 = io_wen & io_addr[10:4] == 7'h22 ? io_wdata[21] : tag_regs_34[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_34 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_314; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_34 = _valid_to_be_T_311 ? io_wdata[20:0] : tag_regs_34[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_34_T = {valid_to_be_34,tag_to_be_34}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_320 = io_wen & io_addr[10:4] == 7'h23; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_323 = io_wen & io_addr[10:4] == 7'h23 ? io_wdata[21] : tag_regs_35[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_35 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_323; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_35 = _valid_to_be_T_320 ? io_wdata[20:0] : tag_regs_35[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_35_T = {valid_to_be_35,tag_to_be_35}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_329 = io_wen & io_addr[10:4] == 7'h24; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_332 = io_wen & io_addr[10:4] == 7'h24 ? io_wdata[21] : tag_regs_36[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_36 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_332; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_36 = _valid_to_be_T_329 ? io_wdata[20:0] : tag_regs_36[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_36_T = {valid_to_be_36,tag_to_be_36}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_338 = io_wen & io_addr[10:4] == 7'h25; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_341 = io_wen & io_addr[10:4] == 7'h25 ? io_wdata[21] : tag_regs_37[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_37 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_341; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_37 = _valid_to_be_T_338 ? io_wdata[20:0] : tag_regs_37[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_37_T = {valid_to_be_37,tag_to_be_37}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_347 = io_wen & io_addr[10:4] == 7'h26; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_350 = io_wen & io_addr[10:4] == 7'h26 ? io_wdata[21] : tag_regs_38[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_38 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_350; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_38 = _valid_to_be_T_347 ? io_wdata[20:0] : tag_regs_38[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_38_T = {valid_to_be_38,tag_to_be_38}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_356 = io_wen & io_addr[10:4] == 7'h27; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_359 = io_wen & io_addr[10:4] == 7'h27 ? io_wdata[21] : tag_regs_39[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_39 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_359; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_39 = _valid_to_be_T_356 ? io_wdata[20:0] : tag_regs_39[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_39_T = {valid_to_be_39,tag_to_be_39}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_365 = io_wen & io_addr[10:4] == 7'h28; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_368 = io_wen & io_addr[10:4] == 7'h28 ? io_wdata[21] : tag_regs_40[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_40 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_368; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_40 = _valid_to_be_T_365 ? io_wdata[20:0] : tag_regs_40[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_40_T = {valid_to_be_40,tag_to_be_40}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_374 = io_wen & io_addr[10:4] == 7'h29; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_377 = io_wen & io_addr[10:4] == 7'h29 ? io_wdata[21] : tag_regs_41[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_41 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_377; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_41 = _valid_to_be_T_374 ? io_wdata[20:0] : tag_regs_41[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_41_T = {valid_to_be_41,tag_to_be_41}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_383 = io_wen & io_addr[10:4] == 7'h2a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_386 = io_wen & io_addr[10:4] == 7'h2a ? io_wdata[21] : tag_regs_42[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_42 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_386; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_42 = _valid_to_be_T_383 ? io_wdata[20:0] : tag_regs_42[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_42_T = {valid_to_be_42,tag_to_be_42}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_392 = io_wen & io_addr[10:4] == 7'h2b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_395 = io_wen & io_addr[10:4] == 7'h2b ? io_wdata[21] : tag_regs_43[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_43 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_395; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_43 = _valid_to_be_T_392 ? io_wdata[20:0] : tag_regs_43[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_43_T = {valid_to_be_43,tag_to_be_43}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_401 = io_wen & io_addr[10:4] == 7'h2c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_404 = io_wen & io_addr[10:4] == 7'h2c ? io_wdata[21] : tag_regs_44[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_44 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_404; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_44 = _valid_to_be_T_401 ? io_wdata[20:0] : tag_regs_44[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_44_T = {valid_to_be_44,tag_to_be_44}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_410 = io_wen & io_addr[10:4] == 7'h2d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_413 = io_wen & io_addr[10:4] == 7'h2d ? io_wdata[21] : tag_regs_45[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_45 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_413; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_45 = _valid_to_be_T_410 ? io_wdata[20:0] : tag_regs_45[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_45_T = {valid_to_be_45,tag_to_be_45}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_419 = io_wen & io_addr[10:4] == 7'h2e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_422 = io_wen & io_addr[10:4] == 7'h2e ? io_wdata[21] : tag_regs_46[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_46 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_422; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_46 = _valid_to_be_T_419 ? io_wdata[20:0] : tag_regs_46[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_46_T = {valid_to_be_46,tag_to_be_46}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_428 = io_wen & io_addr[10:4] == 7'h2f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_431 = io_wen & io_addr[10:4] == 7'h2f ? io_wdata[21] : tag_regs_47[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_47 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_431; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_47 = _valid_to_be_T_428 ? io_wdata[20:0] : tag_regs_47[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_47_T = {valid_to_be_47,tag_to_be_47}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_437 = io_wen & io_addr[10:4] == 7'h30; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_440 = io_wen & io_addr[10:4] == 7'h30 ? io_wdata[21] : tag_regs_48[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_48 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_440; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_48 = _valid_to_be_T_437 ? io_wdata[20:0] : tag_regs_48[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_48_T = {valid_to_be_48,tag_to_be_48}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_446 = io_wen & io_addr[10:4] == 7'h31; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_449 = io_wen & io_addr[10:4] == 7'h31 ? io_wdata[21] : tag_regs_49[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_49 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_449; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_49 = _valid_to_be_T_446 ? io_wdata[20:0] : tag_regs_49[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_49_T = {valid_to_be_49,tag_to_be_49}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_455 = io_wen & io_addr[10:4] == 7'h32; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_458 = io_wen & io_addr[10:4] == 7'h32 ? io_wdata[21] : tag_regs_50[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_50 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_458; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_50 = _valid_to_be_T_455 ? io_wdata[20:0] : tag_regs_50[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_50_T = {valid_to_be_50,tag_to_be_50}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_464 = io_wen & io_addr[10:4] == 7'h33; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_467 = io_wen & io_addr[10:4] == 7'h33 ? io_wdata[21] : tag_regs_51[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_51 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_467; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_51 = _valid_to_be_T_464 ? io_wdata[20:0] : tag_regs_51[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_51_T = {valid_to_be_51,tag_to_be_51}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_473 = io_wen & io_addr[10:4] == 7'h34; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_476 = io_wen & io_addr[10:4] == 7'h34 ? io_wdata[21] : tag_regs_52[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_52 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_476; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_52 = _valid_to_be_T_473 ? io_wdata[20:0] : tag_regs_52[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_52_T = {valid_to_be_52,tag_to_be_52}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_482 = io_wen & io_addr[10:4] == 7'h35; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_485 = io_wen & io_addr[10:4] == 7'h35 ? io_wdata[21] : tag_regs_53[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_53 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_485; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_53 = _valid_to_be_T_482 ? io_wdata[20:0] : tag_regs_53[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_53_T = {valid_to_be_53,tag_to_be_53}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_491 = io_wen & io_addr[10:4] == 7'h36; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_494 = io_wen & io_addr[10:4] == 7'h36 ? io_wdata[21] : tag_regs_54[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_54 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_494; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_54 = _valid_to_be_T_491 ? io_wdata[20:0] : tag_regs_54[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_54_T = {valid_to_be_54,tag_to_be_54}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_500 = io_wen & io_addr[10:4] == 7'h37; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_503 = io_wen & io_addr[10:4] == 7'h37 ? io_wdata[21] : tag_regs_55[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_55 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_503; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_55 = _valid_to_be_T_500 ? io_wdata[20:0] : tag_regs_55[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_55_T = {valid_to_be_55,tag_to_be_55}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_509 = io_wen & io_addr[10:4] == 7'h38; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_512 = io_wen & io_addr[10:4] == 7'h38 ? io_wdata[21] : tag_regs_56[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_56 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_512; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_56 = _valid_to_be_T_509 ? io_wdata[20:0] : tag_regs_56[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_56_T = {valid_to_be_56,tag_to_be_56}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_518 = io_wen & io_addr[10:4] == 7'h39; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_521 = io_wen & io_addr[10:4] == 7'h39 ? io_wdata[21] : tag_regs_57[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_57 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_521; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_57 = _valid_to_be_T_518 ? io_wdata[20:0] : tag_regs_57[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_57_T = {valid_to_be_57,tag_to_be_57}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_527 = io_wen & io_addr[10:4] == 7'h3a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_530 = io_wen & io_addr[10:4] == 7'h3a ? io_wdata[21] : tag_regs_58[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_58 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_530; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_58 = _valid_to_be_T_527 ? io_wdata[20:0] : tag_regs_58[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_58_T = {valid_to_be_58,tag_to_be_58}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_536 = io_wen & io_addr[10:4] == 7'h3b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_539 = io_wen & io_addr[10:4] == 7'h3b ? io_wdata[21] : tag_regs_59[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_59 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_539; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_59 = _valid_to_be_T_536 ? io_wdata[20:0] : tag_regs_59[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_59_T = {valid_to_be_59,tag_to_be_59}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_545 = io_wen & io_addr[10:4] == 7'h3c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_548 = io_wen & io_addr[10:4] == 7'h3c ? io_wdata[21] : tag_regs_60[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_60 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_548; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_60 = _valid_to_be_T_545 ? io_wdata[20:0] : tag_regs_60[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_60_T = {valid_to_be_60,tag_to_be_60}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_554 = io_wen & io_addr[10:4] == 7'h3d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_557 = io_wen & io_addr[10:4] == 7'h3d ? io_wdata[21] : tag_regs_61[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_61 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_557; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_61 = _valid_to_be_T_554 ? io_wdata[20:0] : tag_regs_61[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_61_T = {valid_to_be_61,tag_to_be_61}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_563 = io_wen & io_addr[10:4] == 7'h3e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_566 = io_wen & io_addr[10:4] == 7'h3e ? io_wdata[21] : tag_regs_62[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_62 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_566; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_62 = _valid_to_be_T_563 ? io_wdata[20:0] : tag_regs_62[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_62_T = {valid_to_be_62,tag_to_be_62}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_572 = io_wen & io_addr[10:4] == 7'h3f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_575 = io_wen & io_addr[10:4] == 7'h3f ? io_wdata[21] : tag_regs_63[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_63 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_575; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_63 = _valid_to_be_T_572 ? io_wdata[20:0] : tag_regs_63[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_63_T = {valid_to_be_63,tag_to_be_63}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_581 = io_wen & io_addr[10:4] == 7'h40; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_584 = io_wen & io_addr[10:4] == 7'h40 ? io_wdata[21] : tag_regs_64[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_64 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_584; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_64 = _valid_to_be_T_581 ? io_wdata[20:0] : tag_regs_64[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_64_T = {valid_to_be_64,tag_to_be_64}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_590 = io_wen & io_addr[10:4] == 7'h41; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_593 = io_wen & io_addr[10:4] == 7'h41 ? io_wdata[21] : tag_regs_65[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_65 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_593; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_65 = _valid_to_be_T_590 ? io_wdata[20:0] : tag_regs_65[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_65_T = {valid_to_be_65,tag_to_be_65}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_599 = io_wen & io_addr[10:4] == 7'h42; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_602 = io_wen & io_addr[10:4] == 7'h42 ? io_wdata[21] : tag_regs_66[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_66 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_602; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_66 = _valid_to_be_T_599 ? io_wdata[20:0] : tag_regs_66[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_66_T = {valid_to_be_66,tag_to_be_66}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_608 = io_wen & io_addr[10:4] == 7'h43; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_611 = io_wen & io_addr[10:4] == 7'h43 ? io_wdata[21] : tag_regs_67[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_67 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_611; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_67 = _valid_to_be_T_608 ? io_wdata[20:0] : tag_regs_67[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_67_T = {valid_to_be_67,tag_to_be_67}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_617 = io_wen & io_addr[10:4] == 7'h44; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_620 = io_wen & io_addr[10:4] == 7'h44 ? io_wdata[21] : tag_regs_68[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_68 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_620; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_68 = _valid_to_be_T_617 ? io_wdata[20:0] : tag_regs_68[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_68_T = {valid_to_be_68,tag_to_be_68}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_626 = io_wen & io_addr[10:4] == 7'h45; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_629 = io_wen & io_addr[10:4] == 7'h45 ? io_wdata[21] : tag_regs_69[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_69 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_629; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_69 = _valid_to_be_T_626 ? io_wdata[20:0] : tag_regs_69[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_69_T = {valid_to_be_69,tag_to_be_69}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_635 = io_wen & io_addr[10:4] == 7'h46; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_638 = io_wen & io_addr[10:4] == 7'h46 ? io_wdata[21] : tag_regs_70[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_70 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_638; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_70 = _valid_to_be_T_635 ? io_wdata[20:0] : tag_regs_70[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_70_T = {valid_to_be_70,tag_to_be_70}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_644 = io_wen & io_addr[10:4] == 7'h47; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_647 = io_wen & io_addr[10:4] == 7'h47 ? io_wdata[21] : tag_regs_71[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_71 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_647; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_71 = _valid_to_be_T_644 ? io_wdata[20:0] : tag_regs_71[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_71_T = {valid_to_be_71,tag_to_be_71}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_653 = io_wen & io_addr[10:4] == 7'h48; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_656 = io_wen & io_addr[10:4] == 7'h48 ? io_wdata[21] : tag_regs_72[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_72 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_656; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_72 = _valid_to_be_T_653 ? io_wdata[20:0] : tag_regs_72[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_72_T = {valid_to_be_72,tag_to_be_72}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_662 = io_wen & io_addr[10:4] == 7'h49; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_665 = io_wen & io_addr[10:4] == 7'h49 ? io_wdata[21] : tag_regs_73[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_73 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_665; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_73 = _valid_to_be_T_662 ? io_wdata[20:0] : tag_regs_73[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_73_T = {valid_to_be_73,tag_to_be_73}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_671 = io_wen & io_addr[10:4] == 7'h4a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_674 = io_wen & io_addr[10:4] == 7'h4a ? io_wdata[21] : tag_regs_74[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_74 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_674; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_74 = _valid_to_be_T_671 ? io_wdata[20:0] : tag_regs_74[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_74_T = {valid_to_be_74,tag_to_be_74}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_680 = io_wen & io_addr[10:4] == 7'h4b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_683 = io_wen & io_addr[10:4] == 7'h4b ? io_wdata[21] : tag_regs_75[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_75 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_683; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_75 = _valid_to_be_T_680 ? io_wdata[20:0] : tag_regs_75[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_75_T = {valid_to_be_75,tag_to_be_75}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_689 = io_wen & io_addr[10:4] == 7'h4c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_692 = io_wen & io_addr[10:4] == 7'h4c ? io_wdata[21] : tag_regs_76[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_76 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_692; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_76 = _valid_to_be_T_689 ? io_wdata[20:0] : tag_regs_76[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_76_T = {valid_to_be_76,tag_to_be_76}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_698 = io_wen & io_addr[10:4] == 7'h4d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_701 = io_wen & io_addr[10:4] == 7'h4d ? io_wdata[21] : tag_regs_77[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_77 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_701; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_77 = _valid_to_be_T_698 ? io_wdata[20:0] : tag_regs_77[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_77_T = {valid_to_be_77,tag_to_be_77}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_707 = io_wen & io_addr[10:4] == 7'h4e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_710 = io_wen & io_addr[10:4] == 7'h4e ? io_wdata[21] : tag_regs_78[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_78 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_710; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_78 = _valid_to_be_T_707 ? io_wdata[20:0] : tag_regs_78[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_78_T = {valid_to_be_78,tag_to_be_78}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_716 = io_wen & io_addr[10:4] == 7'h4f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_719 = io_wen & io_addr[10:4] == 7'h4f ? io_wdata[21] : tag_regs_79[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_79 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_719; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_79 = _valid_to_be_T_716 ? io_wdata[20:0] : tag_regs_79[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_79_T = {valid_to_be_79,tag_to_be_79}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_725 = io_wen & io_addr[10:4] == 7'h50; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_728 = io_wen & io_addr[10:4] == 7'h50 ? io_wdata[21] : tag_regs_80[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_80 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_728; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_80 = _valid_to_be_T_725 ? io_wdata[20:0] : tag_regs_80[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_80_T = {valid_to_be_80,tag_to_be_80}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_734 = io_wen & io_addr[10:4] == 7'h51; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_737 = io_wen & io_addr[10:4] == 7'h51 ? io_wdata[21] : tag_regs_81[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_81 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_737; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_81 = _valid_to_be_T_734 ? io_wdata[20:0] : tag_regs_81[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_81_T = {valid_to_be_81,tag_to_be_81}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_743 = io_wen & io_addr[10:4] == 7'h52; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_746 = io_wen & io_addr[10:4] == 7'h52 ? io_wdata[21] : tag_regs_82[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_82 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_746; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_82 = _valid_to_be_T_743 ? io_wdata[20:0] : tag_regs_82[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_82_T = {valid_to_be_82,tag_to_be_82}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_752 = io_wen & io_addr[10:4] == 7'h53; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_755 = io_wen & io_addr[10:4] == 7'h53 ? io_wdata[21] : tag_regs_83[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_83 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_755; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_83 = _valid_to_be_T_752 ? io_wdata[20:0] : tag_regs_83[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_83_T = {valid_to_be_83,tag_to_be_83}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_761 = io_wen & io_addr[10:4] == 7'h54; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_764 = io_wen & io_addr[10:4] == 7'h54 ? io_wdata[21] : tag_regs_84[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_84 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_764; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_84 = _valid_to_be_T_761 ? io_wdata[20:0] : tag_regs_84[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_84_T = {valid_to_be_84,tag_to_be_84}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_770 = io_wen & io_addr[10:4] == 7'h55; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_773 = io_wen & io_addr[10:4] == 7'h55 ? io_wdata[21] : tag_regs_85[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_85 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_773; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_85 = _valid_to_be_T_770 ? io_wdata[20:0] : tag_regs_85[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_85_T = {valid_to_be_85,tag_to_be_85}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_779 = io_wen & io_addr[10:4] == 7'h56; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_782 = io_wen & io_addr[10:4] == 7'h56 ? io_wdata[21] : tag_regs_86[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_86 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_782; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_86 = _valid_to_be_T_779 ? io_wdata[20:0] : tag_regs_86[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_86_T = {valid_to_be_86,tag_to_be_86}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_788 = io_wen & io_addr[10:4] == 7'h57; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_791 = io_wen & io_addr[10:4] == 7'h57 ? io_wdata[21] : tag_regs_87[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_87 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_791; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_87 = _valid_to_be_T_788 ? io_wdata[20:0] : tag_regs_87[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_87_T = {valid_to_be_87,tag_to_be_87}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_797 = io_wen & io_addr[10:4] == 7'h58; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_800 = io_wen & io_addr[10:4] == 7'h58 ? io_wdata[21] : tag_regs_88[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_88 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_800; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_88 = _valid_to_be_T_797 ? io_wdata[20:0] : tag_regs_88[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_88_T = {valid_to_be_88,tag_to_be_88}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_806 = io_wen & io_addr[10:4] == 7'h59; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_809 = io_wen & io_addr[10:4] == 7'h59 ? io_wdata[21] : tag_regs_89[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_89 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_809; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_89 = _valid_to_be_T_806 ? io_wdata[20:0] : tag_regs_89[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_89_T = {valid_to_be_89,tag_to_be_89}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_815 = io_wen & io_addr[10:4] == 7'h5a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_818 = io_wen & io_addr[10:4] == 7'h5a ? io_wdata[21] : tag_regs_90[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_90 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_818; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_90 = _valid_to_be_T_815 ? io_wdata[20:0] : tag_regs_90[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_90_T = {valid_to_be_90,tag_to_be_90}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_824 = io_wen & io_addr[10:4] == 7'h5b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_827 = io_wen & io_addr[10:4] == 7'h5b ? io_wdata[21] : tag_regs_91[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_91 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_827; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_91 = _valid_to_be_T_824 ? io_wdata[20:0] : tag_regs_91[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_91_T = {valid_to_be_91,tag_to_be_91}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_833 = io_wen & io_addr[10:4] == 7'h5c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_836 = io_wen & io_addr[10:4] == 7'h5c ? io_wdata[21] : tag_regs_92[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_92 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_836; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_92 = _valid_to_be_T_833 ? io_wdata[20:0] : tag_regs_92[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_92_T = {valid_to_be_92,tag_to_be_92}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_842 = io_wen & io_addr[10:4] == 7'h5d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_845 = io_wen & io_addr[10:4] == 7'h5d ? io_wdata[21] : tag_regs_93[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_93 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_845; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_93 = _valid_to_be_T_842 ? io_wdata[20:0] : tag_regs_93[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_93_T = {valid_to_be_93,tag_to_be_93}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_851 = io_wen & io_addr[10:4] == 7'h5e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_854 = io_wen & io_addr[10:4] == 7'h5e ? io_wdata[21] : tag_regs_94[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_94 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_854; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_94 = _valid_to_be_T_851 ? io_wdata[20:0] : tag_regs_94[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_94_T = {valid_to_be_94,tag_to_be_94}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_860 = io_wen & io_addr[10:4] == 7'h5f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_863 = io_wen & io_addr[10:4] == 7'h5f ? io_wdata[21] : tag_regs_95[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_95 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_863; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_95 = _valid_to_be_T_860 ? io_wdata[20:0] : tag_regs_95[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_95_T = {valid_to_be_95,tag_to_be_95}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_869 = io_wen & io_addr[10:4] == 7'h60; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_872 = io_wen & io_addr[10:4] == 7'h60 ? io_wdata[21] : tag_regs_96[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_96 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_872; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_96 = _valid_to_be_T_869 ? io_wdata[20:0] : tag_regs_96[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_96_T = {valid_to_be_96,tag_to_be_96}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_878 = io_wen & io_addr[10:4] == 7'h61; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_881 = io_wen & io_addr[10:4] == 7'h61 ? io_wdata[21] : tag_regs_97[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_97 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_881; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_97 = _valid_to_be_T_878 ? io_wdata[20:0] : tag_regs_97[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_97_T = {valid_to_be_97,tag_to_be_97}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_887 = io_wen & io_addr[10:4] == 7'h62; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_890 = io_wen & io_addr[10:4] == 7'h62 ? io_wdata[21] : tag_regs_98[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_98 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_890; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_98 = _valid_to_be_T_887 ? io_wdata[20:0] : tag_regs_98[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_98_T = {valid_to_be_98,tag_to_be_98}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_896 = io_wen & io_addr[10:4] == 7'h63; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_899 = io_wen & io_addr[10:4] == 7'h63 ? io_wdata[21] : tag_regs_99[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_99 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_899; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_99 = _valid_to_be_T_896 ? io_wdata[20:0] : tag_regs_99[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_99_T = {valid_to_be_99,tag_to_be_99}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_905 = io_wen & io_addr[10:4] == 7'h64; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_908 = io_wen & io_addr[10:4] == 7'h64 ? io_wdata[21] : tag_regs_100[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_100 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_908; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_100 = _valid_to_be_T_905 ? io_wdata[20:0] : tag_regs_100[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_100_T = {valid_to_be_100,tag_to_be_100}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_914 = io_wen & io_addr[10:4] == 7'h65; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_917 = io_wen & io_addr[10:4] == 7'h65 ? io_wdata[21] : tag_regs_101[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_101 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_917; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_101 = _valid_to_be_T_914 ? io_wdata[20:0] : tag_regs_101[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_101_T = {valid_to_be_101,tag_to_be_101}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_923 = io_wen & io_addr[10:4] == 7'h66; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_926 = io_wen & io_addr[10:4] == 7'h66 ? io_wdata[21] : tag_regs_102[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_102 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_926; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_102 = _valid_to_be_T_923 ? io_wdata[20:0] : tag_regs_102[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_102_T = {valid_to_be_102,tag_to_be_102}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_932 = io_wen & io_addr[10:4] == 7'h67; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_935 = io_wen & io_addr[10:4] == 7'h67 ? io_wdata[21] : tag_regs_103[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_103 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_935; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_103 = _valid_to_be_T_932 ? io_wdata[20:0] : tag_regs_103[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_103_T = {valid_to_be_103,tag_to_be_103}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_941 = io_wen & io_addr[10:4] == 7'h68; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_944 = io_wen & io_addr[10:4] == 7'h68 ? io_wdata[21] : tag_regs_104[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_104 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_944; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_104 = _valid_to_be_T_941 ? io_wdata[20:0] : tag_regs_104[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_104_T = {valid_to_be_104,tag_to_be_104}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_950 = io_wen & io_addr[10:4] == 7'h69; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_953 = io_wen & io_addr[10:4] == 7'h69 ? io_wdata[21] : tag_regs_105[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_105 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_953; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_105 = _valid_to_be_T_950 ? io_wdata[20:0] : tag_regs_105[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_105_T = {valid_to_be_105,tag_to_be_105}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_959 = io_wen & io_addr[10:4] == 7'h6a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_962 = io_wen & io_addr[10:4] == 7'h6a ? io_wdata[21] : tag_regs_106[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_106 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_962; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_106 = _valid_to_be_T_959 ? io_wdata[20:0] : tag_regs_106[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_106_T = {valid_to_be_106,tag_to_be_106}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_968 = io_wen & io_addr[10:4] == 7'h6b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_971 = io_wen & io_addr[10:4] == 7'h6b ? io_wdata[21] : tag_regs_107[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_107 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_971; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_107 = _valid_to_be_T_968 ? io_wdata[20:0] : tag_regs_107[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_107_T = {valid_to_be_107,tag_to_be_107}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_977 = io_wen & io_addr[10:4] == 7'h6c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_980 = io_wen & io_addr[10:4] == 7'h6c ? io_wdata[21] : tag_regs_108[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_108 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_980; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_108 = _valid_to_be_T_977 ? io_wdata[20:0] : tag_regs_108[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_108_T = {valid_to_be_108,tag_to_be_108}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_986 = io_wen & io_addr[10:4] == 7'h6d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_989 = io_wen & io_addr[10:4] == 7'h6d ? io_wdata[21] : tag_regs_109[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_109 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_989; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_109 = _valid_to_be_T_986 ? io_wdata[20:0] : tag_regs_109[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_109_T = {valid_to_be_109,tag_to_be_109}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_995 = io_wen & io_addr[10:4] == 7'h6e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_998 = io_wen & io_addr[10:4] == 7'h6e ? io_wdata[21] : tag_regs_110[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_110 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_998; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_110 = _valid_to_be_T_995 ? io_wdata[20:0] : tag_regs_110[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_110_T = {valid_to_be_110,tag_to_be_110}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1004 = io_wen & io_addr[10:4] == 7'h6f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1007 = io_wen & io_addr[10:4] == 7'h6f ? io_wdata[21] : tag_regs_111[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_111 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1007; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_111 = _valid_to_be_T_1004 ? io_wdata[20:0] : tag_regs_111[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_111_T = {valid_to_be_111,tag_to_be_111}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1013 = io_wen & io_addr[10:4] == 7'h70; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1016 = io_wen & io_addr[10:4] == 7'h70 ? io_wdata[21] : tag_regs_112[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_112 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1016; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_112 = _valid_to_be_T_1013 ? io_wdata[20:0] : tag_regs_112[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_112_T = {valid_to_be_112,tag_to_be_112}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1022 = io_wen & io_addr[10:4] == 7'h71; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1025 = io_wen & io_addr[10:4] == 7'h71 ? io_wdata[21] : tag_regs_113[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_113 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1025; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_113 = _valid_to_be_T_1022 ? io_wdata[20:0] : tag_regs_113[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_113_T = {valid_to_be_113,tag_to_be_113}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1031 = io_wen & io_addr[10:4] == 7'h72; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1034 = io_wen & io_addr[10:4] == 7'h72 ? io_wdata[21] : tag_regs_114[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_114 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1034; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_114 = _valid_to_be_T_1031 ? io_wdata[20:0] : tag_regs_114[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_114_T = {valid_to_be_114,tag_to_be_114}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1040 = io_wen & io_addr[10:4] == 7'h73; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1043 = io_wen & io_addr[10:4] == 7'h73 ? io_wdata[21] : tag_regs_115[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_115 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1043; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_115 = _valid_to_be_T_1040 ? io_wdata[20:0] : tag_regs_115[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_115_T = {valid_to_be_115,tag_to_be_115}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1049 = io_wen & io_addr[10:4] == 7'h74; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1052 = io_wen & io_addr[10:4] == 7'h74 ? io_wdata[21] : tag_regs_116[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_116 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1052; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_116 = _valid_to_be_T_1049 ? io_wdata[20:0] : tag_regs_116[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_116_T = {valid_to_be_116,tag_to_be_116}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1058 = io_wen & io_addr[10:4] == 7'h75; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1061 = io_wen & io_addr[10:4] == 7'h75 ? io_wdata[21] : tag_regs_117[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_117 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1061; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_117 = _valid_to_be_T_1058 ? io_wdata[20:0] : tag_regs_117[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_117_T = {valid_to_be_117,tag_to_be_117}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1067 = io_wen & io_addr[10:4] == 7'h76; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1070 = io_wen & io_addr[10:4] == 7'h76 ? io_wdata[21] : tag_regs_118[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_118 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1070; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_118 = _valid_to_be_T_1067 ? io_wdata[20:0] : tag_regs_118[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_118_T = {valid_to_be_118,tag_to_be_118}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1076 = io_wen & io_addr[10:4] == 7'h77; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1079 = io_wen & io_addr[10:4] == 7'h77 ? io_wdata[21] : tag_regs_119[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_119 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1079; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_119 = _valid_to_be_T_1076 ? io_wdata[20:0] : tag_regs_119[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_119_T = {valid_to_be_119,tag_to_be_119}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1085 = io_wen & io_addr[10:4] == 7'h78; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1088 = io_wen & io_addr[10:4] == 7'h78 ? io_wdata[21] : tag_regs_120[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_120 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1088; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_120 = _valid_to_be_T_1085 ? io_wdata[20:0] : tag_regs_120[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_120_T = {valid_to_be_120,tag_to_be_120}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1094 = io_wen & io_addr[10:4] == 7'h79; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1097 = io_wen & io_addr[10:4] == 7'h79 ? io_wdata[21] : tag_regs_121[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_121 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1097; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_121 = _valid_to_be_T_1094 ? io_wdata[20:0] : tag_regs_121[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_121_T = {valid_to_be_121,tag_to_be_121}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1103 = io_wen & io_addr[10:4] == 7'h7a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1106 = io_wen & io_addr[10:4] == 7'h7a ? io_wdata[21] : tag_regs_122[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_122 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1106; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_122 = _valid_to_be_T_1103 ? io_wdata[20:0] : tag_regs_122[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_122_T = {valid_to_be_122,tag_to_be_122}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1112 = io_wen & io_addr[10:4] == 7'h7b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1115 = io_wen & io_addr[10:4] == 7'h7b ? io_wdata[21] : tag_regs_123[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_123 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1115; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_123 = _valid_to_be_T_1112 ? io_wdata[20:0] : tag_regs_123[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_123_T = {valid_to_be_123,tag_to_be_123}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1121 = io_wen & io_addr[10:4] == 7'h7c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1124 = io_wen & io_addr[10:4] == 7'h7c ? io_wdata[21] : tag_regs_124[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_124 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1124; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_124 = _valid_to_be_T_1121 ? io_wdata[20:0] : tag_regs_124[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_124_T = {valid_to_be_124,tag_to_be_124}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1130 = io_wen & io_addr[10:4] == 7'h7d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1133 = io_wen & io_addr[10:4] == 7'h7d ? io_wdata[21] : tag_regs_125[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_125 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1133; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_125 = _valid_to_be_T_1130 ? io_wdata[20:0] : tag_regs_125[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_125_T = {valid_to_be_125,tag_to_be_125}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1139 = io_wen & io_addr[10:4] == 7'h7e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1142 = io_wen & io_addr[10:4] == 7'h7e ? io_wdata[21] : tag_regs_126[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_126 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1142; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_126 = _valid_to_be_T_1139 ? io_wdata[20:0] : tag_regs_126[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_126_T = {valid_to_be_126,tag_to_be_126}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1148 = io_wen & io_addr[10:4] == 7'h7f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1151 = io_wen & io_addr[10:4] == 7'h7f ? io_wdata[21] : tag_regs_127[21]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_127 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1151; // @[icache_tag.scala 27:30]
  wire [20:0] tag_to_be_127 = _valid_to_be_T_1148 ? io_wdata[20:0] : tag_regs_127[20:0]; // @[icache_tag.scala 30:28]
  wire [21:0] _tag_regs_127_T = {valid_to_be_127,tag_to_be_127}; // @[Cat.scala 31:58]
  wire [21:0] _GEN_1 = 7'h1 == io_addr[10:4] ? tag_regs_1 : tag_regs_0; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_2 = 7'h2 == io_addr[10:4] ? tag_regs_2 : _GEN_1; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_3 = 7'h3 == io_addr[10:4] ? tag_regs_3 : _GEN_2; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_4 = 7'h4 == io_addr[10:4] ? tag_regs_4 : _GEN_3; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_5 = 7'h5 == io_addr[10:4] ? tag_regs_5 : _GEN_4; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_6 = 7'h6 == io_addr[10:4] ? tag_regs_6 : _GEN_5; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_7 = 7'h7 == io_addr[10:4] ? tag_regs_7 : _GEN_6; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_8 = 7'h8 == io_addr[10:4] ? tag_regs_8 : _GEN_7; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_9 = 7'h9 == io_addr[10:4] ? tag_regs_9 : _GEN_8; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_10 = 7'ha == io_addr[10:4] ? tag_regs_10 : _GEN_9; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_11 = 7'hb == io_addr[10:4] ? tag_regs_11 : _GEN_10; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_12 = 7'hc == io_addr[10:4] ? tag_regs_12 : _GEN_11; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_13 = 7'hd == io_addr[10:4] ? tag_regs_13 : _GEN_12; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_14 = 7'he == io_addr[10:4] ? tag_regs_14 : _GEN_13; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_15 = 7'hf == io_addr[10:4] ? tag_regs_15 : _GEN_14; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_16 = 7'h10 == io_addr[10:4] ? tag_regs_16 : _GEN_15; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_17 = 7'h11 == io_addr[10:4] ? tag_regs_17 : _GEN_16; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_18 = 7'h12 == io_addr[10:4] ? tag_regs_18 : _GEN_17; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_19 = 7'h13 == io_addr[10:4] ? tag_regs_19 : _GEN_18; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_20 = 7'h14 == io_addr[10:4] ? tag_regs_20 : _GEN_19; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_21 = 7'h15 == io_addr[10:4] ? tag_regs_21 : _GEN_20; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_22 = 7'h16 == io_addr[10:4] ? tag_regs_22 : _GEN_21; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_23 = 7'h17 == io_addr[10:4] ? tag_regs_23 : _GEN_22; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_24 = 7'h18 == io_addr[10:4] ? tag_regs_24 : _GEN_23; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_25 = 7'h19 == io_addr[10:4] ? tag_regs_25 : _GEN_24; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_26 = 7'h1a == io_addr[10:4] ? tag_regs_26 : _GEN_25; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_27 = 7'h1b == io_addr[10:4] ? tag_regs_27 : _GEN_26; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_28 = 7'h1c == io_addr[10:4] ? tag_regs_28 : _GEN_27; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_29 = 7'h1d == io_addr[10:4] ? tag_regs_29 : _GEN_28; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_30 = 7'h1e == io_addr[10:4] ? tag_regs_30 : _GEN_29; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_31 = 7'h1f == io_addr[10:4] ? tag_regs_31 : _GEN_30; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_32 = 7'h20 == io_addr[10:4] ? tag_regs_32 : _GEN_31; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_33 = 7'h21 == io_addr[10:4] ? tag_regs_33 : _GEN_32; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_34 = 7'h22 == io_addr[10:4] ? tag_regs_34 : _GEN_33; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_35 = 7'h23 == io_addr[10:4] ? tag_regs_35 : _GEN_34; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_36 = 7'h24 == io_addr[10:4] ? tag_regs_36 : _GEN_35; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_37 = 7'h25 == io_addr[10:4] ? tag_regs_37 : _GEN_36; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_38 = 7'h26 == io_addr[10:4] ? tag_regs_38 : _GEN_37; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_39 = 7'h27 == io_addr[10:4] ? tag_regs_39 : _GEN_38; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_40 = 7'h28 == io_addr[10:4] ? tag_regs_40 : _GEN_39; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_41 = 7'h29 == io_addr[10:4] ? tag_regs_41 : _GEN_40; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_42 = 7'h2a == io_addr[10:4] ? tag_regs_42 : _GEN_41; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_43 = 7'h2b == io_addr[10:4] ? tag_regs_43 : _GEN_42; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_44 = 7'h2c == io_addr[10:4] ? tag_regs_44 : _GEN_43; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_45 = 7'h2d == io_addr[10:4] ? tag_regs_45 : _GEN_44; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_46 = 7'h2e == io_addr[10:4] ? tag_regs_46 : _GEN_45; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_47 = 7'h2f == io_addr[10:4] ? tag_regs_47 : _GEN_46; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_48 = 7'h30 == io_addr[10:4] ? tag_regs_48 : _GEN_47; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_49 = 7'h31 == io_addr[10:4] ? tag_regs_49 : _GEN_48; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_50 = 7'h32 == io_addr[10:4] ? tag_regs_50 : _GEN_49; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_51 = 7'h33 == io_addr[10:4] ? tag_regs_51 : _GEN_50; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_52 = 7'h34 == io_addr[10:4] ? tag_regs_52 : _GEN_51; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_53 = 7'h35 == io_addr[10:4] ? tag_regs_53 : _GEN_52; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_54 = 7'h36 == io_addr[10:4] ? tag_regs_54 : _GEN_53; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_55 = 7'h37 == io_addr[10:4] ? tag_regs_55 : _GEN_54; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_56 = 7'h38 == io_addr[10:4] ? tag_regs_56 : _GEN_55; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_57 = 7'h39 == io_addr[10:4] ? tag_regs_57 : _GEN_56; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_58 = 7'h3a == io_addr[10:4] ? tag_regs_58 : _GEN_57; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_59 = 7'h3b == io_addr[10:4] ? tag_regs_59 : _GEN_58; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_60 = 7'h3c == io_addr[10:4] ? tag_regs_60 : _GEN_59; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_61 = 7'h3d == io_addr[10:4] ? tag_regs_61 : _GEN_60; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_62 = 7'h3e == io_addr[10:4] ? tag_regs_62 : _GEN_61; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_63 = 7'h3f == io_addr[10:4] ? tag_regs_63 : _GEN_62; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_64 = 7'h40 == io_addr[10:4] ? tag_regs_64 : _GEN_63; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_65 = 7'h41 == io_addr[10:4] ? tag_regs_65 : _GEN_64; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_66 = 7'h42 == io_addr[10:4] ? tag_regs_66 : _GEN_65; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_67 = 7'h43 == io_addr[10:4] ? tag_regs_67 : _GEN_66; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_68 = 7'h44 == io_addr[10:4] ? tag_regs_68 : _GEN_67; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_69 = 7'h45 == io_addr[10:4] ? tag_regs_69 : _GEN_68; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_70 = 7'h46 == io_addr[10:4] ? tag_regs_70 : _GEN_69; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_71 = 7'h47 == io_addr[10:4] ? tag_regs_71 : _GEN_70; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_72 = 7'h48 == io_addr[10:4] ? tag_regs_72 : _GEN_71; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_73 = 7'h49 == io_addr[10:4] ? tag_regs_73 : _GEN_72; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_74 = 7'h4a == io_addr[10:4] ? tag_regs_74 : _GEN_73; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_75 = 7'h4b == io_addr[10:4] ? tag_regs_75 : _GEN_74; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_76 = 7'h4c == io_addr[10:4] ? tag_regs_76 : _GEN_75; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_77 = 7'h4d == io_addr[10:4] ? tag_regs_77 : _GEN_76; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_78 = 7'h4e == io_addr[10:4] ? tag_regs_78 : _GEN_77; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_79 = 7'h4f == io_addr[10:4] ? tag_regs_79 : _GEN_78; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_80 = 7'h50 == io_addr[10:4] ? tag_regs_80 : _GEN_79; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_81 = 7'h51 == io_addr[10:4] ? tag_regs_81 : _GEN_80; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_82 = 7'h52 == io_addr[10:4] ? tag_regs_82 : _GEN_81; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_83 = 7'h53 == io_addr[10:4] ? tag_regs_83 : _GEN_82; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_84 = 7'h54 == io_addr[10:4] ? tag_regs_84 : _GEN_83; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_85 = 7'h55 == io_addr[10:4] ? tag_regs_85 : _GEN_84; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_86 = 7'h56 == io_addr[10:4] ? tag_regs_86 : _GEN_85; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_87 = 7'h57 == io_addr[10:4] ? tag_regs_87 : _GEN_86; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_88 = 7'h58 == io_addr[10:4] ? tag_regs_88 : _GEN_87; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_89 = 7'h59 == io_addr[10:4] ? tag_regs_89 : _GEN_88; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_90 = 7'h5a == io_addr[10:4] ? tag_regs_90 : _GEN_89; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_91 = 7'h5b == io_addr[10:4] ? tag_regs_91 : _GEN_90; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_92 = 7'h5c == io_addr[10:4] ? tag_regs_92 : _GEN_91; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_93 = 7'h5d == io_addr[10:4] ? tag_regs_93 : _GEN_92; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_94 = 7'h5e == io_addr[10:4] ? tag_regs_94 : _GEN_93; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_95 = 7'h5f == io_addr[10:4] ? tag_regs_95 : _GEN_94; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_96 = 7'h60 == io_addr[10:4] ? tag_regs_96 : _GEN_95; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_97 = 7'h61 == io_addr[10:4] ? tag_regs_97 : _GEN_96; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_98 = 7'h62 == io_addr[10:4] ? tag_regs_98 : _GEN_97; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_99 = 7'h63 == io_addr[10:4] ? tag_regs_99 : _GEN_98; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_100 = 7'h64 == io_addr[10:4] ? tag_regs_100 : _GEN_99; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_101 = 7'h65 == io_addr[10:4] ? tag_regs_101 : _GEN_100; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_102 = 7'h66 == io_addr[10:4] ? tag_regs_102 : _GEN_101; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_103 = 7'h67 == io_addr[10:4] ? tag_regs_103 : _GEN_102; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_104 = 7'h68 == io_addr[10:4] ? tag_regs_104 : _GEN_103; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_105 = 7'h69 == io_addr[10:4] ? tag_regs_105 : _GEN_104; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_106 = 7'h6a == io_addr[10:4] ? tag_regs_106 : _GEN_105; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_107 = 7'h6b == io_addr[10:4] ? tag_regs_107 : _GEN_106; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_108 = 7'h6c == io_addr[10:4] ? tag_regs_108 : _GEN_107; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_109 = 7'h6d == io_addr[10:4] ? tag_regs_109 : _GEN_108; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_110 = 7'h6e == io_addr[10:4] ? tag_regs_110 : _GEN_109; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_111 = 7'h6f == io_addr[10:4] ? tag_regs_111 : _GEN_110; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_112 = 7'h70 == io_addr[10:4] ? tag_regs_112 : _GEN_111; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_113 = 7'h71 == io_addr[10:4] ? tag_regs_113 : _GEN_112; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_114 = 7'h72 == io_addr[10:4] ? tag_regs_114 : _GEN_113; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_115 = 7'h73 == io_addr[10:4] ? tag_regs_115 : _GEN_114; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_116 = 7'h74 == io_addr[10:4] ? tag_regs_116 : _GEN_115; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_117 = 7'h75 == io_addr[10:4] ? tag_regs_117 : _GEN_116; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_118 = 7'h76 == io_addr[10:4] ? tag_regs_118 : _GEN_117; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_119 = 7'h77 == io_addr[10:4] ? tag_regs_119 : _GEN_118; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_120 = 7'h78 == io_addr[10:4] ? tag_regs_120 : _GEN_119; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_121 = 7'h79 == io_addr[10:4] ? tag_regs_121 : _GEN_120; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_122 = 7'h7a == io_addr[10:4] ? tag_regs_122 : _GEN_121; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_123 = 7'h7b == io_addr[10:4] ? tag_regs_123 : _GEN_122; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_124 = 7'h7c == io_addr[10:4] ? tag_regs_124 : _GEN_123; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_125 = 7'h7d == io_addr[10:4] ? tag_regs_125 : _GEN_124; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_126 = 7'h7e == io_addr[10:4] ? tag_regs_126 : _GEN_125; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_127 = 7'h7f == io_addr[10:4] ? tag_regs_127 : _GEN_126; // @[icache_tag.scala 36:{22,22}]
  assign io_hit = _GEN_127[20:0] == io_addr[31:11]; // @[icache_tag.scala 37:31]
  assign io_valid = _GEN_127[21]; // @[icache_tag.scala 36:22]
  always @(posedge clock) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_0 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_0 <= _tag_regs_0_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_1 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_1 <= _tag_regs_1_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_2 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_2 <= _tag_regs_2_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_3 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_3 <= _tag_regs_3_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_4 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_4 <= _tag_regs_4_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_5 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_5 <= _tag_regs_5_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_6 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_6 <= _tag_regs_6_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_7 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_7 <= _tag_regs_7_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_8 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_8 <= _tag_regs_8_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_9 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_9 <= _tag_regs_9_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_10 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_10 <= _tag_regs_10_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_11 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_11 <= _tag_regs_11_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_12 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_12 <= _tag_regs_12_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_13 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_13 <= _tag_regs_13_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_14 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_14 <= _tag_regs_14_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_15 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_15 <= _tag_regs_15_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_16 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_16 <= _tag_regs_16_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_17 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_17 <= _tag_regs_17_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_18 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_18 <= _tag_regs_18_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_19 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_19 <= _tag_regs_19_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_20 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_20 <= _tag_regs_20_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_21 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_21 <= _tag_regs_21_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_22 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_22 <= _tag_regs_22_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_23 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_23 <= _tag_regs_23_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_24 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_24 <= _tag_regs_24_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_25 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_25 <= _tag_regs_25_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_26 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_26 <= _tag_regs_26_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_27 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_27 <= _tag_regs_27_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_28 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_28 <= _tag_regs_28_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_29 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_29 <= _tag_regs_29_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_30 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_30 <= _tag_regs_30_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_31 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_31 <= _tag_regs_31_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_32 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_32 <= _tag_regs_32_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_33 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_33 <= _tag_regs_33_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_34 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_34 <= _tag_regs_34_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_35 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_35 <= _tag_regs_35_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_36 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_36 <= _tag_regs_36_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_37 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_37 <= _tag_regs_37_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_38 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_38 <= _tag_regs_38_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_39 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_39 <= _tag_regs_39_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_40 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_40 <= _tag_regs_40_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_41 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_41 <= _tag_regs_41_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_42 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_42 <= _tag_regs_42_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_43 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_43 <= _tag_regs_43_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_44 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_44 <= _tag_regs_44_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_45 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_45 <= _tag_regs_45_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_46 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_46 <= _tag_regs_46_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_47 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_47 <= _tag_regs_47_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_48 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_48 <= _tag_regs_48_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_49 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_49 <= _tag_regs_49_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_50 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_50 <= _tag_regs_50_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_51 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_51 <= _tag_regs_51_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_52 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_52 <= _tag_regs_52_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_53 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_53 <= _tag_regs_53_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_54 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_54 <= _tag_regs_54_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_55 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_55 <= _tag_regs_55_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_56 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_56 <= _tag_regs_56_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_57 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_57 <= _tag_regs_57_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_58 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_58 <= _tag_regs_58_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_59 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_59 <= _tag_regs_59_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_60 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_60 <= _tag_regs_60_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_61 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_61 <= _tag_regs_61_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_62 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_62 <= _tag_regs_62_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_63 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_63 <= _tag_regs_63_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_64 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_64 <= _tag_regs_64_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_65 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_65 <= _tag_regs_65_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_66 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_66 <= _tag_regs_66_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_67 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_67 <= _tag_regs_67_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_68 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_68 <= _tag_regs_68_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_69 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_69 <= _tag_regs_69_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_70 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_70 <= _tag_regs_70_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_71 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_71 <= _tag_regs_71_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_72 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_72 <= _tag_regs_72_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_73 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_73 <= _tag_regs_73_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_74 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_74 <= _tag_regs_74_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_75 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_75 <= _tag_regs_75_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_76 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_76 <= _tag_regs_76_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_77 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_77 <= _tag_regs_77_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_78 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_78 <= _tag_regs_78_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_79 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_79 <= _tag_regs_79_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_80 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_80 <= _tag_regs_80_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_81 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_81 <= _tag_regs_81_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_82 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_82 <= _tag_regs_82_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_83 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_83 <= _tag_regs_83_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_84 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_84 <= _tag_regs_84_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_85 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_85 <= _tag_regs_85_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_86 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_86 <= _tag_regs_86_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_87 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_87 <= _tag_regs_87_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_88 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_88 <= _tag_regs_88_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_89 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_89 <= _tag_regs_89_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_90 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_90 <= _tag_regs_90_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_91 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_91 <= _tag_regs_91_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_92 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_92 <= _tag_regs_92_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_93 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_93 <= _tag_regs_93_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_94 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_94 <= _tag_regs_94_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_95 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_95 <= _tag_regs_95_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_96 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_96 <= _tag_regs_96_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_97 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_97 <= _tag_regs_97_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_98 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_98 <= _tag_regs_98_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_99 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_99 <= _tag_regs_99_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_100 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_100 <= _tag_regs_100_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_101 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_101 <= _tag_regs_101_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_102 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_102 <= _tag_regs_102_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_103 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_103 <= _tag_regs_103_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_104 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_104 <= _tag_regs_104_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_105 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_105 <= _tag_regs_105_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_106 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_106 <= _tag_regs_106_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_107 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_107 <= _tag_regs_107_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_108 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_108 <= _tag_regs_108_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_109 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_109 <= _tag_regs_109_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_110 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_110 <= _tag_regs_110_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_111 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_111 <= _tag_regs_111_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_112 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_112 <= _tag_regs_112_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_113 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_113 <= _tag_regs_113_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_114 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_114 <= _tag_regs_114_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_115 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_115 <= _tag_regs_115_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_116 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_116 <= _tag_regs_116_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_117 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_117 <= _tag_regs_117_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_118 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_118 <= _tag_regs_118_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_119 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_119 <= _tag_regs_119_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_120 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_120 <= _tag_regs_120_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_121 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_121 <= _tag_regs_121_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_122 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_122 <= _tag_regs_122_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_123 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_123 <= _tag_regs_123_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_124 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_124 <= _tag_regs_124_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_125 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_125 <= _tag_regs_125_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_126 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_126 <= _tag_regs_126_T; // @[icache_tag.scala 31:25]
    end
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_127 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_127 <= _tag_regs_127_T; // @[icache_tag.scala 31:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_regs_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_regs_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_regs_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_regs_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_regs_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_regs_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_regs_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_regs_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_regs_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_regs_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_regs_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_regs_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_regs_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_regs_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_regs_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_regs_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_regs_16 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_regs_17 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_regs_18 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_regs_19 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_regs_20 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_regs_21 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_regs_22 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_regs_23 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_regs_24 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_regs_25 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_regs_26 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_regs_27 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_regs_28 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_regs_29 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_regs_30 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_regs_31 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_regs_32 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_regs_33 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_regs_34 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_regs_35 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_regs_36 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_regs_37 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_regs_38 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_regs_39 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_regs_40 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_regs_41 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_regs_42 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_regs_43 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_regs_44 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_regs_45 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_regs_46 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_regs_47 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_regs_48 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_regs_49 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_regs_50 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_regs_51 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_regs_52 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_regs_53 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_regs_54 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_regs_55 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_regs_56 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_regs_57 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_regs_58 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_regs_59 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_regs_60 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_regs_61 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_regs_62 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_regs_63 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  tag_regs_64 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  tag_regs_65 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tag_regs_66 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tag_regs_67 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tag_regs_68 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tag_regs_69 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tag_regs_70 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tag_regs_71 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tag_regs_72 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tag_regs_73 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tag_regs_74 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tag_regs_75 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tag_regs_76 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tag_regs_77 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tag_regs_78 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tag_regs_79 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tag_regs_80 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tag_regs_81 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tag_regs_82 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tag_regs_83 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tag_regs_84 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tag_regs_85 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tag_regs_86 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tag_regs_87 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tag_regs_88 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tag_regs_89 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tag_regs_90 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tag_regs_91 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tag_regs_92 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tag_regs_93 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tag_regs_94 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tag_regs_95 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tag_regs_96 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tag_regs_97 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tag_regs_98 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tag_regs_99 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tag_regs_100 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tag_regs_101 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tag_regs_102 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tag_regs_103 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tag_regs_104 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tag_regs_105 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tag_regs_106 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tag_regs_107 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tag_regs_108 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tag_regs_109 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tag_regs_110 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tag_regs_111 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tag_regs_112 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tag_regs_113 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tag_regs_114 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tag_regs_115 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tag_regs_116 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tag_regs_117 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tag_regs_118 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tag_regs_119 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tag_regs_120 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tag_regs_121 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tag_regs_122 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tag_regs_123 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tag_regs_124 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tag_regs_125 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tag_regs_126 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tag_regs_127 = _RAND_127[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_ysyx_sram_with_mask(
  input          clock,
  input  [7:0]   io_wea,
  input  [6:0]   io_addra,
  input  [63:0]  io_dina,
  output [63:0]  io_douta,
  output [5:0]   io_sram_port_addr,
  output         io_sram_port_wen,
  output [127:0] io_sram_port_wmask,
  output [127:0] io_sram_port_wdata,
  input  [127:0] io_sram_port_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] final_write_data_1 = {io_dina, 64'h0}; // @[ip_user.scala 163:44]
  wire [7:0] ena_budle__0 = io_wea[0] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__1 = io_wea[1] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__2 = io_wea[2] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__3 = io_wea[3] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__4 = io_wea[4] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__5 = io_wea[5] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__6 = io_wea[6] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [7:0] ena_budle__7 = io_wea[7] ? 8'h0 : 8'hff; // @[ip_user.scala 168:35]
  wire [63:0] _final_ena_data_0_T_2 = {ena_budle__7,ena_budle__6,ena_budle__5,ena_budle__4,ena_budle__3,ena_budle__2,
    ena_budle__1,ena_budle__0}; // @[ip_user.scala 170:96]
  wire [63:0] final_ena_data_0 = ~io_addra[0] ? _final_ena_data_0_T_2 : 64'hffffffffffffffff; // @[ip_user.scala 170:38]
  wire [63:0] final_ena_data_1 = io_addra[0] ? _final_ena_data_0_T_2 : 64'hffffffffffffffff; // @[ip_user.scala 170:38]
  wire [127:0] final_write_data_0 = {{64'd0}, io_dina}; // @[ip_user.scala 160:32 163:33]
  reg [6:0] addr_reg; // @[ip_user.scala 178:28]
  wire  shift_num = addr_reg[0]; // @[ip_user.scala 179:30]
  wire [63:0] sram_data_bundle_0 = io_sram_port_rdata[63:0]; // @[ip_user.scala 182:54]
  wire [63:0] sram_data_bundle_1 = io_sram_port_rdata[127:64]; // @[ip_user.scala 182:54]
  assign io_douta = shift_num ? sram_data_bundle_1 : sram_data_bundle_0; // @[ip_user.scala 184:{14,14}]
  assign io_sram_port_addr = io_addra[6:1]; // @[ip_user.scala 177:34]
  assign io_sram_port_wen = io_wea == 8'h0; // @[ip_user.scala 157:32]
  assign io_sram_port_wmask = {final_ena_data_1,final_ena_data_0}; // @[ip_user.scala 176:42]
  assign io_sram_port_wdata = io_addra[0] ? final_write_data_1 : final_write_data_0; // @[ip_user.scala 175:{24,24}]
  always @(posedge clock) begin
    addr_reg <= io_addra; // @[ip_user.scala 178:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_icache_data(
  input          clock,
  input  [7:0]   io_wen,
  input  [31:0]  io_addr,
  input  [63:0]  io_wdata,
  output [39:0]  io_rdata,
  output [5:0]   io_sram_addr,
  output         io_sram_wen,
  output [127:0] io_sram_wmask,
  output [127:0] io_sram_wdata,
  input  [127:0] io_sram_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  icache_data_ram_0_clock; // @[icache_data.scala 32:35]
  wire [7:0] icache_data_ram_0_io_wea; // @[icache_data.scala 32:35]
  wire [6:0] icache_data_ram_0_io_addra; // @[icache_data.scala 32:35]
  wire [63:0] icache_data_ram_0_io_dina; // @[icache_data.scala 32:35]
  wire [63:0] icache_data_ram_0_io_douta; // @[icache_data.scala 32:35]
  wire [5:0] icache_data_ram_0_io_sram_port_addr; // @[icache_data.scala 32:35]
  wire  icache_data_ram_0_io_sram_port_wen; // @[icache_data.scala 32:35]
  wire [127:0] icache_data_ram_0_io_sram_port_wmask; // @[icache_data.scala 32:35]
  wire [127:0] icache_data_ram_0_io_sram_port_wdata; // @[icache_data.scala 32:35]
  wire [127:0] icache_data_ram_0_io_sram_port_rdata; // @[icache_data.scala 32:35]
  reg [31:0] addr_reg; // @[icache_data.scala 38:27]
  wire [31:0] get_data = addr_reg[2] ? icache_data_ram_0_io_douta[63:32] : icache_data_ram_0_io_douta[31:0]; // @[icache_data.scala 40:26]
  wire [6:0] io_rdata_opD = get_data[6:0]; // @[macros.scala 532:24]
  wire [2:0] io_rdata_Funct3D = get_data[14:12]; // @[macros.scala 533:28]
  wire [1:0] _io_rdata_T_3 = 3'h1 == io_rdata_Funct3D ? 2'h2 : {{1'd0}, 3'h0 == io_rdata_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _io_rdata_T_5 = 3'h4 == io_rdata_Funct3D ? 3'h4 : {{1'd0}, _io_rdata_T_3}; // @[Mux.scala 81:58]
  wire [3:0] _io_rdata_T_7 = 3'h5 == io_rdata_Funct3D ? 4'h8 : {{1'd0}, _io_rdata_T_5}; // @[Mux.scala 81:58]
  wire [4:0] _io_rdata_T_9 = 3'h6 == io_rdata_Funct3D ? 5'h10 : {{1'd0}, _io_rdata_T_7}; // @[Mux.scala 81:58]
  wire [5:0] _io_rdata_T_11 = 3'h7 == io_rdata_Funct3D ? 6'h20 : {{1'd0}, _io_rdata_T_9}; // @[Mux.scala 81:58]
  wire [5:0] _io_rdata_T_13 = 7'h63 == io_rdata_opD ? _io_rdata_T_11 : 6'h0; // @[Mux.scala 81:58]
  wire  _io_rdata_T_16 = io_rdata_opD == 7'h67 & io_rdata_Funct3D == 3'h0; // @[macros.scala 505:30]
  wire  _io_rdata_T_18 = _io_rdata_T_16 | io_rdata_opD == 7'h6f; // @[macros.scala 510:27]
  wire  _io_rdata_T_19 = io_rdata_opD == 7'h63; // @[macros.scala 528:13]
  wire [32:0] io_rdata_lo = {_io_rdata_T_19,get_data}; // @[Cat.scala 31:58]
  wire [6:0] io_rdata_hi = {_io_rdata_T_13,_io_rdata_T_18}; // @[Cat.scala 31:58]
  ysyx_22040886_ysyx_sram_with_mask icache_data_ram_0 ( // @[icache_data.scala 32:35]
    .clock(icache_data_ram_0_clock),
    .io_wea(icache_data_ram_0_io_wea),
    .io_addra(icache_data_ram_0_io_addra),
    .io_dina(icache_data_ram_0_io_dina),
    .io_douta(icache_data_ram_0_io_douta),
    .io_sram_port_addr(icache_data_ram_0_io_sram_port_addr),
    .io_sram_port_wen(icache_data_ram_0_io_sram_port_wen),
    .io_sram_port_wmask(icache_data_ram_0_io_sram_port_wmask),
    .io_sram_port_wdata(icache_data_ram_0_io_sram_port_wdata),
    .io_sram_port_rdata(icache_data_ram_0_io_sram_port_rdata)
  );
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[Cat.scala 31:58]
  assign io_sram_addr = icache_data_ram_0_io_sram_port_addr; // @[icache_data.scala 37:13]
  assign io_sram_wen = icache_data_ram_0_io_sram_port_wen; // @[icache_data.scala 37:13]
  assign io_sram_wmask = icache_data_ram_0_io_sram_port_wmask; // @[icache_data.scala 37:13]
  assign io_sram_wdata = icache_data_ram_0_io_sram_port_wdata; // @[icache_data.scala 37:13]
  assign icache_data_ram_0_clock = clock;
  assign icache_data_ram_0_io_wea = io_wen; // @[icache_data.scala 34:31]
  assign icache_data_ram_0_io_addra = io_addr[10:4]; // @[icache_data.scala 35:42]
  assign icache_data_ram_0_io_dina = io_wdata; // @[icache_data.scala 36:31]
  assign icache_data_ram_0_io_sram_port_rdata = io_sram_rdata; // @[icache_data.scala 37:13]
  always @(posedge clock) begin
    addr_reg <= io_addr; // @[icache_data.scala 38:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_inst_cache(
  input          clock,
  input          reset,
  output [31:0]  io_port_araddr,
  output [7:0]   io_port_arlen,
  output [2:0]   io_port_arsize,
  output [1:0]   io_port_arburst,
  output         io_port_arvalid,
  input          io_port_arready,
  input  [63:0]  io_port_rdata,
  input          io_port_rlast,
  input          io_port_rvalid,
  input          io_stage2_flush,
  output         io_stage2_stall,
  input          io_stage1_valid_flush,
  input          io_inst_ready_to_use,
  input          io_inst_buffer_full,
  output [63:0]  io_v_addr_for_tlb,
  input  [63:0]  io_p_addr_for_tlb,
  input          io_sram_req,
  input  [63:0]  io_sram_addr,
  output [1:0]   io_sram_write_en,
  output [39:0]  io_sram_rdata_L,
  input          io_sram_cache,
  input          io_tag_valid_flush,
  output [5:0]   io_sram_0_addr,
  output         io_sram_0_wen,
  output [127:0] io_sram_0_wmask,
  output [127:0] io_sram_0_wdata,
  input  [127:0] io_sram_0_rdata,
  output [5:0]   io_sram_1_addr,
  output         io_sram_1_wen,
  output [127:0] io_sram_1_wmask,
  output [127:0] io_sram_1_wdata,
  input  [127:0] io_sram_1_rdata,
  output [5:0]   io_sram_2_addr,
  output         io_sram_2_wen,
  output [127:0] io_sram_2_wmask,
  output [127:0] io_sram_2_wdata,
  input  [127:0] io_sram_2_rdata,
  output [5:0]   io_sram_3_addr,
  output         io_sram_3_wen,
  output [127:0] io_sram_3_wmask,
  output [127:0] io_sram_3_wdata,
  input  [127:0] io_sram_3_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [63:0] _RAND_142;
`endif // RANDOMIZE_REG_INIT
  wire  icache_tag_clock; // @[inst_cache.scala 83:34]
  wire  icache_tag_reset; // @[inst_cache.scala 83:34]
  wire  icache_tag_io_wen; // @[inst_cache.scala 83:34]
  wire [21:0] icache_tag_io_wdata; // @[inst_cache.scala 83:34]
  wire [31:0] icache_tag_io_addr; // @[inst_cache.scala 83:34]
  wire  icache_tag_io_hit; // @[inst_cache.scala 83:34]
  wire  icache_tag_io_valid; // @[inst_cache.scala 83:34]
  wire  icache_tag_io_tag_all_flush; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_clock; // @[inst_cache.scala 85:34]
  wire  icache_tag_1_reset; // @[inst_cache.scala 85:34]
  wire  icache_tag_1_io_wen; // @[inst_cache.scala 85:34]
  wire [21:0] icache_tag_1_io_wdata; // @[inst_cache.scala 85:34]
  wire [31:0] icache_tag_1_io_addr; // @[inst_cache.scala 85:34]
  wire  icache_tag_1_io_hit; // @[inst_cache.scala 85:34]
  wire  icache_tag_1_io_valid; // @[inst_cache.scala 85:34]
  wire  icache_tag_1_io_tag_all_flush; // @[inst_cache.scala 85:34]
  wire  icache_data_clock; // @[inst_cache.scala 91:55]
  wire [7:0] icache_data_io_wen; // @[inst_cache.scala 91:55]
  wire [31:0] icache_data_io_addr; // @[inst_cache.scala 91:55]
  wire [63:0] icache_data_io_wdata; // @[inst_cache.scala 91:55]
  wire [39:0] icache_data_io_rdata; // @[inst_cache.scala 91:55]
  wire [5:0] icache_data_io_sram_addr; // @[inst_cache.scala 91:55]
  wire  icache_data_io_sram_wen; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_io_sram_wmask; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_io_sram_wdata; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_io_sram_rdata; // @[inst_cache.scala 91:55]
  wire  icache_data_1_clock; // @[inst_cache.scala 91:55]
  wire [7:0] icache_data_1_io_wen; // @[inst_cache.scala 91:55]
  wire [31:0] icache_data_1_io_addr; // @[inst_cache.scala 91:55]
  wire [63:0] icache_data_1_io_wdata; // @[inst_cache.scala 91:55]
  wire [39:0] icache_data_1_io_rdata; // @[inst_cache.scala 91:55]
  wire [5:0] icache_data_1_io_sram_addr; // @[inst_cache.scala 91:55]
  wire  icache_data_1_io_sram_wen; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_1_io_sram_wmask; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_1_io_sram_wdata; // @[inst_cache.scala 91:55]
  wire [127:0] icache_data_1_io_sram_rdata; // @[inst_cache.scala 91:55]
  wire  icache_data_2_clock; // @[inst_cache.scala 92:55]
  wire [7:0] icache_data_2_io_wen; // @[inst_cache.scala 92:55]
  wire [31:0] icache_data_2_io_addr; // @[inst_cache.scala 92:55]
  wire [63:0] icache_data_2_io_wdata; // @[inst_cache.scala 92:55]
  wire [39:0] icache_data_2_io_rdata; // @[inst_cache.scala 92:55]
  wire [5:0] icache_data_2_io_sram_addr; // @[inst_cache.scala 92:55]
  wire  icache_data_2_io_sram_wen; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_2_io_sram_wmask; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_2_io_sram_wdata; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_2_io_sram_rdata; // @[inst_cache.scala 92:55]
  wire  icache_data_3_clock; // @[inst_cache.scala 92:55]
  wire [7:0] icache_data_3_io_wen; // @[inst_cache.scala 92:55]
  wire [31:0] icache_data_3_io_addr; // @[inst_cache.scala 92:55]
  wire [63:0] icache_data_3_io_wdata; // @[inst_cache.scala 92:55]
  wire [39:0] icache_data_3_io_rdata; // @[inst_cache.scala 92:55]
  wire [5:0] icache_data_3_io_sram_addr; // @[inst_cache.scala 92:55]
  wire  icache_data_3_io_sram_wen; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_3_io_sram_wmask; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_3_io_sram_wdata; // @[inst_cache.scala 92:55]
  wire [127:0] icache_data_3_io_sram_rdata; // @[inst_cache.scala 92:55]
  reg  lru_0; // @[inst_cache.scala 76:22]
  reg  lru_1; // @[inst_cache.scala 76:22]
  reg  lru_2; // @[inst_cache.scala 76:22]
  reg  lru_3; // @[inst_cache.scala 76:22]
  reg  lru_4; // @[inst_cache.scala 76:22]
  reg  lru_5; // @[inst_cache.scala 76:22]
  reg  lru_6; // @[inst_cache.scala 76:22]
  reg  lru_7; // @[inst_cache.scala 76:22]
  reg  lru_8; // @[inst_cache.scala 76:22]
  reg  lru_9; // @[inst_cache.scala 76:22]
  reg  lru_10; // @[inst_cache.scala 76:22]
  reg  lru_11; // @[inst_cache.scala 76:22]
  reg  lru_12; // @[inst_cache.scala 76:22]
  reg  lru_13; // @[inst_cache.scala 76:22]
  reg  lru_14; // @[inst_cache.scala 76:22]
  reg  lru_15; // @[inst_cache.scala 76:22]
  reg  lru_16; // @[inst_cache.scala 76:22]
  reg  lru_17; // @[inst_cache.scala 76:22]
  reg  lru_18; // @[inst_cache.scala 76:22]
  reg  lru_19; // @[inst_cache.scala 76:22]
  reg  lru_20; // @[inst_cache.scala 76:22]
  reg  lru_21; // @[inst_cache.scala 76:22]
  reg  lru_22; // @[inst_cache.scala 76:22]
  reg  lru_23; // @[inst_cache.scala 76:22]
  reg  lru_24; // @[inst_cache.scala 76:22]
  reg  lru_25; // @[inst_cache.scala 76:22]
  reg  lru_26; // @[inst_cache.scala 76:22]
  reg  lru_27; // @[inst_cache.scala 76:22]
  reg  lru_28; // @[inst_cache.scala 76:22]
  reg  lru_29; // @[inst_cache.scala 76:22]
  reg  lru_30; // @[inst_cache.scala 76:22]
  reg  lru_31; // @[inst_cache.scala 76:22]
  reg  lru_32; // @[inst_cache.scala 76:22]
  reg  lru_33; // @[inst_cache.scala 76:22]
  reg  lru_34; // @[inst_cache.scala 76:22]
  reg  lru_35; // @[inst_cache.scala 76:22]
  reg  lru_36; // @[inst_cache.scala 76:22]
  reg  lru_37; // @[inst_cache.scala 76:22]
  reg  lru_38; // @[inst_cache.scala 76:22]
  reg  lru_39; // @[inst_cache.scala 76:22]
  reg  lru_40; // @[inst_cache.scala 76:22]
  reg  lru_41; // @[inst_cache.scala 76:22]
  reg  lru_42; // @[inst_cache.scala 76:22]
  reg  lru_43; // @[inst_cache.scala 76:22]
  reg  lru_44; // @[inst_cache.scala 76:22]
  reg  lru_45; // @[inst_cache.scala 76:22]
  reg  lru_46; // @[inst_cache.scala 76:22]
  reg  lru_47; // @[inst_cache.scala 76:22]
  reg  lru_48; // @[inst_cache.scala 76:22]
  reg  lru_49; // @[inst_cache.scala 76:22]
  reg  lru_50; // @[inst_cache.scala 76:22]
  reg  lru_51; // @[inst_cache.scala 76:22]
  reg  lru_52; // @[inst_cache.scala 76:22]
  reg  lru_53; // @[inst_cache.scala 76:22]
  reg  lru_54; // @[inst_cache.scala 76:22]
  reg  lru_55; // @[inst_cache.scala 76:22]
  reg  lru_56; // @[inst_cache.scala 76:22]
  reg  lru_57; // @[inst_cache.scala 76:22]
  reg  lru_58; // @[inst_cache.scala 76:22]
  reg  lru_59; // @[inst_cache.scala 76:22]
  reg  lru_60; // @[inst_cache.scala 76:22]
  reg  lru_61; // @[inst_cache.scala 76:22]
  reg  lru_62; // @[inst_cache.scala 76:22]
  reg  lru_63; // @[inst_cache.scala 76:22]
  reg  lru_64; // @[inst_cache.scala 76:22]
  reg  lru_65; // @[inst_cache.scala 76:22]
  reg  lru_66; // @[inst_cache.scala 76:22]
  reg  lru_67; // @[inst_cache.scala 76:22]
  reg  lru_68; // @[inst_cache.scala 76:22]
  reg  lru_69; // @[inst_cache.scala 76:22]
  reg  lru_70; // @[inst_cache.scala 76:22]
  reg  lru_71; // @[inst_cache.scala 76:22]
  reg  lru_72; // @[inst_cache.scala 76:22]
  reg  lru_73; // @[inst_cache.scala 76:22]
  reg  lru_74; // @[inst_cache.scala 76:22]
  reg  lru_75; // @[inst_cache.scala 76:22]
  reg  lru_76; // @[inst_cache.scala 76:22]
  reg  lru_77; // @[inst_cache.scala 76:22]
  reg  lru_78; // @[inst_cache.scala 76:22]
  reg  lru_79; // @[inst_cache.scala 76:22]
  reg  lru_80; // @[inst_cache.scala 76:22]
  reg  lru_81; // @[inst_cache.scala 76:22]
  reg  lru_82; // @[inst_cache.scala 76:22]
  reg  lru_83; // @[inst_cache.scala 76:22]
  reg  lru_84; // @[inst_cache.scala 76:22]
  reg  lru_85; // @[inst_cache.scala 76:22]
  reg  lru_86; // @[inst_cache.scala 76:22]
  reg  lru_87; // @[inst_cache.scala 76:22]
  reg  lru_88; // @[inst_cache.scala 76:22]
  reg  lru_89; // @[inst_cache.scala 76:22]
  reg  lru_90; // @[inst_cache.scala 76:22]
  reg  lru_91; // @[inst_cache.scala 76:22]
  reg  lru_92; // @[inst_cache.scala 76:22]
  reg  lru_93; // @[inst_cache.scala 76:22]
  reg  lru_94; // @[inst_cache.scala 76:22]
  reg  lru_95; // @[inst_cache.scala 76:22]
  reg  lru_96; // @[inst_cache.scala 76:22]
  reg  lru_97; // @[inst_cache.scala 76:22]
  reg  lru_98; // @[inst_cache.scala 76:22]
  reg  lru_99; // @[inst_cache.scala 76:22]
  reg  lru_100; // @[inst_cache.scala 76:22]
  reg  lru_101; // @[inst_cache.scala 76:22]
  reg  lru_102; // @[inst_cache.scala 76:22]
  reg  lru_103; // @[inst_cache.scala 76:22]
  reg  lru_104; // @[inst_cache.scala 76:22]
  reg  lru_105; // @[inst_cache.scala 76:22]
  reg  lru_106; // @[inst_cache.scala 76:22]
  reg  lru_107; // @[inst_cache.scala 76:22]
  reg  lru_108; // @[inst_cache.scala 76:22]
  reg  lru_109; // @[inst_cache.scala 76:22]
  reg  lru_110; // @[inst_cache.scala 76:22]
  reg  lru_111; // @[inst_cache.scala 76:22]
  reg  lru_112; // @[inst_cache.scala 76:22]
  reg  lru_113; // @[inst_cache.scala 76:22]
  reg  lru_114; // @[inst_cache.scala 76:22]
  reg  lru_115; // @[inst_cache.scala 76:22]
  reg  lru_116; // @[inst_cache.scala 76:22]
  reg  lru_117; // @[inst_cache.scala 76:22]
  reg  lru_118; // @[inst_cache.scala 76:22]
  reg  lru_119; // @[inst_cache.scala 76:22]
  reg  lru_120; // @[inst_cache.scala 76:22]
  reg  lru_121; // @[inst_cache.scala 76:22]
  reg  lru_122; // @[inst_cache.scala 76:22]
  reg  lru_123; // @[inst_cache.scala 76:22]
  reg  lru_124; // @[inst_cache.scala 76:22]
  reg  lru_125; // @[inst_cache.scala 76:22]
  reg  lru_126; // @[inst_cache.scala 76:22]
  reg  lru_127; // @[inst_cache.scala 76:22]
  reg [3:0] work_state; // @[inst_cache.scala 108:29]
  reg [2:0] write_counter; // @[inst_cache.scala 110:33]
  reg [39:0] wait_data_L; // @[inst_cache.scala 111:31]
  wire  stage1_flush = ~io_sram_req & io_stage1_valid_flush; // @[inst_cache.scala 115:35]
  reg  stage1_stall_reg; // @[inst_cache.scala 122:35]
  reg [63:0] stage1_addr_line_mapping; // @[Reg.scala 28:20]
  reg [63:0] stage1_sram_phy_addr_reg; // @[inst_cache.scala 126:43]
  reg  stage1_sram_cache_reg; // @[Reg.scala 28:20]
  wire  _stage1_sram_req_reg_T_1 = io_sram_req | stage1_flush; // @[inst_cache.scala 128:106]
  reg  stage1_sram_req_reg; // @[Reg.scala 28:20]
  reg  stage1_finished; // @[inst_cache.scala 131:34]
  wire  _stage1_finished_T_1 = work_state == 4'h7; // @[inst_cache.scala 147:67]
  wire  _stage1_finished_T_2 = work_state == 4'h3; // @[inst_cache.scala 147:103]
  wire  _access_work_state_T = work_state == 4'h2; // @[inst_cache.scala 251:41]
  wire  _access_work_state_T_6 = io_port_rlast & io_port_rvalid; // @[inst_cache.scala 252:71]
  wire [2:0] _access_work_state_T_7 = io_port_rlast & io_port_rvalid ? 3'h4 : 3'h3; // @[inst_cache.scala 252:49]
  wire  _access_work_state_T_8 = work_state == 4'h4; // @[inst_cache.scala 253:23]
  wire  _hit_T = icache_tag_io_hit; // @[inst_cache.scala 178:33]
  wire  _hit_T_2 = icache_tag_io_hit & icache_tag_io_valid; // @[inst_cache.scala 178:40]
  wire  _hit_T_3 = icache_tag_1_io_hit; // @[inst_cache.scala 179:27]
  wire  _hit_T_5 = icache_tag_1_io_hit & icache_tag_1_io_valid; // @[inst_cache.scala 179:34]
  wire  hit = icache_tag_io_hit & icache_tag_io_valid | _hit_T_5; // @[inst_cache.scala 178:70]
  wire [2:0] _access_work_state_T_13 = stage1_finished ? 3'h4 : 3'h2; // @[inst_cache.scala 253:145]
  wire [2:0] _access_work_state_T_14 = stage1_sram_cache_reg ? 3'h1 : _access_work_state_T_13; // @[inst_cache.scala 253:99]
  wire [2:0] _access_work_state_T_15 = stage1_sram_req_reg ? _access_work_state_T_14 : 3'h1; // @[inst_cache.scala 253:68]
  wire [2:0] _access_work_state_T_18 = stage1_finished ? 3'h4 : 3'h5; // @[inst_cache.scala 254:79]
  wire [2:0] _access_work_state_T_20 = stage1_sram_cache_reg ? _access_work_state_T_18 : _access_work_state_T_13; // @[inst_cache.scala 254:46]
  wire [2:0] _access_work_state_T_21 = stage1_sram_req_reg ? _access_work_state_T_20 : 3'h1; // @[inst_cache.scala 254:15]
  wire [2:0] _access_work_state_T_22 = hit ? _access_work_state_T_15 : _access_work_state_T_21; // @[inst_cache.scala 253:46]
  wire  _access_work_state_T_23 = work_state == 4'h1; // @[inst_cache.scala 256:23]
  wire [1:0] _access_work_state_T_28 = stage1_sram_cache_reg ? 2'h1 : 2'h2; // @[inst_cache.scala 256:95]
  wire [1:0] _access_work_state_T_29 = stage1_sram_req_reg ? _access_work_state_T_28 : 2'h1; // @[inst_cache.scala 256:64]
  wire [2:0] _access_work_state_T_32 = stage1_sram_cache_reg ? 3'h5 : 3'h2; // @[inst_cache.scala 257:46]
  wire [2:0] _access_work_state_T_33 = stage1_sram_req_reg ? _access_work_state_T_32 : 3'h1; // @[inst_cache.scala 257:15]
  wire [2:0] _access_work_state_T_34 = hit ? {{1'd0}, _access_work_state_T_29} : _access_work_state_T_33; // @[inst_cache.scala 256:42]
  wire  _access_work_state_T_35 = work_state == 4'h5; // @[inst_cache.scala 258:23]
  wire  _access_work_state_T_38 = work_state == 4'h6; // @[inst_cache.scala 259:23]
  wire [3:0] _access_work_state_T_42 = _access_work_state_T_6 ? 4'h7 : work_state; // @[inst_cache.scala 259:54]
  wire [3:0] _access_work_state_T_44 = _stage1_finished_T_1 ? 4'h4 : work_state; // @[inst_cache.scala 260:12]
  wire [3:0] _access_work_state_T_45 = work_state == 4'h6 ? _access_work_state_T_42 : _access_work_state_T_44; // @[inst_cache.scala 259:12]
  wire [3:0] _access_work_state_T_46 = work_state == 4'h5 & io_port_arready ? 4'h6 : _access_work_state_T_45; // @[inst_cache.scala 258:12]
  wire [3:0] _access_work_state_T_47 = work_state == 4'h1 ? {{1'd0}, _access_work_state_T_34} : _access_work_state_T_46; // @[inst_cache.scala 256:12]
  wire [3:0] _access_work_state_T_48 = work_state == 4'h4 ? {{1'd0}, _access_work_state_T_22} : _access_work_state_T_47; // @[inst_cache.scala 253:12]
  wire [3:0] _access_work_state_T_49 = _stage1_finished_T_2 ? {{1'd0}, _access_work_state_T_7} : _access_work_state_T_48
    ; // @[inst_cache.scala 252:12]
  wire [3:0] access_work_state = work_state == 4'h2 & io_port_arready ? 4'h3 : _access_work_state_T_49; // @[inst_cache.scala 251:30]
  wire  _stage2_stall_T = access_work_state == 4'h1; // @[inst_cache.scala 152:40]
  wire  _stage2_stall_T_5 = ~io_inst_buffer_full; // @[inst_cache.scala 153:11]
  wire  stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4) & _stage2_stall_T_5; // @[inst_cache.scala 152:129]
  wire [6:0] decoder_inst_data_0_opD = io_port_rdata[6:0]; // @[macros.scala 532:24]
  wire [2:0] decoder_inst_data_0_Funct3D = io_port_rdata[14:12]; // @[macros.scala 533:28]
  wire [1:0] _decoder_inst_data_0_T_4 = 3'h1 == decoder_inst_data_0_Funct3D ? 2'h2 : {{1'd0}, 3'h0 ==
    decoder_inst_data_0_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _decoder_inst_data_0_T_6 = 3'h4 == decoder_inst_data_0_Funct3D ? 3'h4 : {{1'd0}, _decoder_inst_data_0_T_4}; // @[Mux.scala 81:58]
  wire [3:0] _decoder_inst_data_0_T_8 = 3'h5 == decoder_inst_data_0_Funct3D ? 4'h8 : {{1'd0}, _decoder_inst_data_0_T_6}; // @[Mux.scala 81:58]
  wire [4:0] _decoder_inst_data_0_T_10 = 3'h6 == decoder_inst_data_0_Funct3D ? 5'h10 : {{1'd0}, _decoder_inst_data_0_T_8
    }; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_0_T_12 = 3'h7 == decoder_inst_data_0_Funct3D ? 6'h20 : {{1'd0},
    _decoder_inst_data_0_T_10}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_0_T_14 = 7'h63 == decoder_inst_data_0_opD ? _decoder_inst_data_0_T_12 : 6'h0; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_0_T_18 = decoder_inst_data_0_opD == 7'h67 & decoder_inst_data_0_Funct3D == 3'h0; // @[macros.scala 505:30]
  wire  _decoder_inst_data_0_T_20 = _decoder_inst_data_0_T_18 | decoder_inst_data_0_opD == 7'h6f; // @[macros.scala 510:27]
  wire  _decoder_inst_data_0_T_22 = decoder_inst_data_0_opD == 7'h63; // @[macros.scala 528:13]
  wire [39:0] decoder_inst_data_0 = {_decoder_inst_data_0_T_14,_decoder_inst_data_0_T_20,_decoder_inst_data_0_T_22,
    io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [6:0] decoder_inst_data_1_opD = io_port_rdata[38:32]; // @[macros.scala 532:24]
  wire [2:0] decoder_inst_data_1_Funct3D = io_port_rdata[46:44]; // @[macros.scala 533:28]
  wire [1:0] _decoder_inst_data_1_T_4 = 3'h1 == decoder_inst_data_1_Funct3D ? 2'h2 : {{1'd0}, 3'h0 ==
    decoder_inst_data_1_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _decoder_inst_data_1_T_6 = 3'h4 == decoder_inst_data_1_Funct3D ? 3'h4 : {{1'd0}, _decoder_inst_data_1_T_4}; // @[Mux.scala 81:58]
  wire [3:0] _decoder_inst_data_1_T_8 = 3'h5 == decoder_inst_data_1_Funct3D ? 4'h8 : {{1'd0}, _decoder_inst_data_1_T_6}; // @[Mux.scala 81:58]
  wire [4:0] _decoder_inst_data_1_T_10 = 3'h6 == decoder_inst_data_1_Funct3D ? 5'h10 : {{1'd0}, _decoder_inst_data_1_T_8
    }; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_1_T_12 = 3'h7 == decoder_inst_data_1_Funct3D ? 6'h20 : {{1'd0},
    _decoder_inst_data_1_T_10}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_1_T_14 = 7'h63 == decoder_inst_data_1_opD ? _decoder_inst_data_1_T_12 : 6'h0; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_1_T_18 = decoder_inst_data_1_opD == 7'h67 & decoder_inst_data_1_Funct3D == 3'h0; // @[macros.scala 505:30]
  wire  _decoder_inst_data_1_T_20 = _decoder_inst_data_1_T_18 | decoder_inst_data_1_opD == 7'h6f; // @[macros.scala 510:27]
  wire  _decoder_inst_data_1_T_22 = decoder_inst_data_1_opD == 7'h63; // @[macros.scala 528:13]
  wire [39:0] decoder_inst_data_1 = {_decoder_inst_data_1_T_14,_decoder_inst_data_1_T_20,_decoder_inst_data_1_T_22,
    io_port_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [39:0] decoder_inst_data = stage1_addr_line_mapping[2] ? decoder_inst_data_1 : decoder_inst_data_0; // @[inst_cache.scala 163:33]
  wire  _GEN_4 = 7'h1 == stage1_addr_line_mapping[10:4] ? lru_1 : lru_0; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_5 = 7'h2 == stage1_addr_line_mapping[10:4] ? lru_2 : _GEN_4; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_6 = 7'h3 == stage1_addr_line_mapping[10:4] ? lru_3 : _GEN_5; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_7 = 7'h4 == stage1_addr_line_mapping[10:4] ? lru_4 : _GEN_6; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_8 = 7'h5 == stage1_addr_line_mapping[10:4] ? lru_5 : _GEN_7; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_9 = 7'h6 == stage1_addr_line_mapping[10:4] ? lru_6 : _GEN_8; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_10 = 7'h7 == stage1_addr_line_mapping[10:4] ? lru_7 : _GEN_9; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_11 = 7'h8 == stage1_addr_line_mapping[10:4] ? lru_8 : _GEN_10; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_12 = 7'h9 == stage1_addr_line_mapping[10:4] ? lru_9 : _GEN_11; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_13 = 7'ha == stage1_addr_line_mapping[10:4] ? lru_10 : _GEN_12; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_14 = 7'hb == stage1_addr_line_mapping[10:4] ? lru_11 : _GEN_13; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_15 = 7'hc == stage1_addr_line_mapping[10:4] ? lru_12 : _GEN_14; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_16 = 7'hd == stage1_addr_line_mapping[10:4] ? lru_13 : _GEN_15; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_17 = 7'he == stage1_addr_line_mapping[10:4] ? lru_14 : _GEN_16; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_18 = 7'hf == stage1_addr_line_mapping[10:4] ? lru_15 : _GEN_17; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_19 = 7'h10 == stage1_addr_line_mapping[10:4] ? lru_16 : _GEN_18; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_20 = 7'h11 == stage1_addr_line_mapping[10:4] ? lru_17 : _GEN_19; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_21 = 7'h12 == stage1_addr_line_mapping[10:4] ? lru_18 : _GEN_20; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_22 = 7'h13 == stage1_addr_line_mapping[10:4] ? lru_19 : _GEN_21; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_23 = 7'h14 == stage1_addr_line_mapping[10:4] ? lru_20 : _GEN_22; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_24 = 7'h15 == stage1_addr_line_mapping[10:4] ? lru_21 : _GEN_23; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_25 = 7'h16 == stage1_addr_line_mapping[10:4] ? lru_22 : _GEN_24; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_26 = 7'h17 == stage1_addr_line_mapping[10:4] ? lru_23 : _GEN_25; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_27 = 7'h18 == stage1_addr_line_mapping[10:4] ? lru_24 : _GEN_26; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_28 = 7'h19 == stage1_addr_line_mapping[10:4] ? lru_25 : _GEN_27; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_29 = 7'h1a == stage1_addr_line_mapping[10:4] ? lru_26 : _GEN_28; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_30 = 7'h1b == stage1_addr_line_mapping[10:4] ? lru_27 : _GEN_29; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_31 = 7'h1c == stage1_addr_line_mapping[10:4] ? lru_28 : _GEN_30; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_32 = 7'h1d == stage1_addr_line_mapping[10:4] ? lru_29 : _GEN_31; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_33 = 7'h1e == stage1_addr_line_mapping[10:4] ? lru_30 : _GEN_32; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_34 = 7'h1f == stage1_addr_line_mapping[10:4] ? lru_31 : _GEN_33; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_35 = 7'h20 == stage1_addr_line_mapping[10:4] ? lru_32 : _GEN_34; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_36 = 7'h21 == stage1_addr_line_mapping[10:4] ? lru_33 : _GEN_35; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_37 = 7'h22 == stage1_addr_line_mapping[10:4] ? lru_34 : _GEN_36; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_38 = 7'h23 == stage1_addr_line_mapping[10:4] ? lru_35 : _GEN_37; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_39 = 7'h24 == stage1_addr_line_mapping[10:4] ? lru_36 : _GEN_38; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_40 = 7'h25 == stage1_addr_line_mapping[10:4] ? lru_37 : _GEN_39; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_41 = 7'h26 == stage1_addr_line_mapping[10:4] ? lru_38 : _GEN_40; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_42 = 7'h27 == stage1_addr_line_mapping[10:4] ? lru_39 : _GEN_41; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_43 = 7'h28 == stage1_addr_line_mapping[10:4] ? lru_40 : _GEN_42; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_44 = 7'h29 == stage1_addr_line_mapping[10:4] ? lru_41 : _GEN_43; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_45 = 7'h2a == stage1_addr_line_mapping[10:4] ? lru_42 : _GEN_44; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_46 = 7'h2b == stage1_addr_line_mapping[10:4] ? lru_43 : _GEN_45; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_47 = 7'h2c == stage1_addr_line_mapping[10:4] ? lru_44 : _GEN_46; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_48 = 7'h2d == stage1_addr_line_mapping[10:4] ? lru_45 : _GEN_47; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_49 = 7'h2e == stage1_addr_line_mapping[10:4] ? lru_46 : _GEN_48; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_50 = 7'h2f == stage1_addr_line_mapping[10:4] ? lru_47 : _GEN_49; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_51 = 7'h30 == stage1_addr_line_mapping[10:4] ? lru_48 : _GEN_50; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_52 = 7'h31 == stage1_addr_line_mapping[10:4] ? lru_49 : _GEN_51; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_53 = 7'h32 == stage1_addr_line_mapping[10:4] ? lru_50 : _GEN_52; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_54 = 7'h33 == stage1_addr_line_mapping[10:4] ? lru_51 : _GEN_53; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_55 = 7'h34 == stage1_addr_line_mapping[10:4] ? lru_52 : _GEN_54; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_56 = 7'h35 == stage1_addr_line_mapping[10:4] ? lru_53 : _GEN_55; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_57 = 7'h36 == stage1_addr_line_mapping[10:4] ? lru_54 : _GEN_56; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_58 = 7'h37 == stage1_addr_line_mapping[10:4] ? lru_55 : _GEN_57; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_59 = 7'h38 == stage1_addr_line_mapping[10:4] ? lru_56 : _GEN_58; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_60 = 7'h39 == stage1_addr_line_mapping[10:4] ? lru_57 : _GEN_59; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_61 = 7'h3a == stage1_addr_line_mapping[10:4] ? lru_58 : _GEN_60; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_62 = 7'h3b == stage1_addr_line_mapping[10:4] ? lru_59 : _GEN_61; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_63 = 7'h3c == stage1_addr_line_mapping[10:4] ? lru_60 : _GEN_62; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_64 = 7'h3d == stage1_addr_line_mapping[10:4] ? lru_61 : _GEN_63; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_65 = 7'h3e == stage1_addr_line_mapping[10:4] ? lru_62 : _GEN_64; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_66 = 7'h3f == stage1_addr_line_mapping[10:4] ? lru_63 : _GEN_65; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_67 = 7'h40 == stage1_addr_line_mapping[10:4] ? lru_64 : _GEN_66; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_68 = 7'h41 == stage1_addr_line_mapping[10:4] ? lru_65 : _GEN_67; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_69 = 7'h42 == stage1_addr_line_mapping[10:4] ? lru_66 : _GEN_68; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_70 = 7'h43 == stage1_addr_line_mapping[10:4] ? lru_67 : _GEN_69; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_71 = 7'h44 == stage1_addr_line_mapping[10:4] ? lru_68 : _GEN_70; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_72 = 7'h45 == stage1_addr_line_mapping[10:4] ? lru_69 : _GEN_71; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_73 = 7'h46 == stage1_addr_line_mapping[10:4] ? lru_70 : _GEN_72; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_74 = 7'h47 == stage1_addr_line_mapping[10:4] ? lru_71 : _GEN_73; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_75 = 7'h48 == stage1_addr_line_mapping[10:4] ? lru_72 : _GEN_74; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_76 = 7'h49 == stage1_addr_line_mapping[10:4] ? lru_73 : _GEN_75; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_77 = 7'h4a == stage1_addr_line_mapping[10:4] ? lru_74 : _GEN_76; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_78 = 7'h4b == stage1_addr_line_mapping[10:4] ? lru_75 : _GEN_77; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_79 = 7'h4c == stage1_addr_line_mapping[10:4] ? lru_76 : _GEN_78; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_80 = 7'h4d == stage1_addr_line_mapping[10:4] ? lru_77 : _GEN_79; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_81 = 7'h4e == stage1_addr_line_mapping[10:4] ? lru_78 : _GEN_80; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_82 = 7'h4f == stage1_addr_line_mapping[10:4] ? lru_79 : _GEN_81; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_83 = 7'h50 == stage1_addr_line_mapping[10:4] ? lru_80 : _GEN_82; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_84 = 7'h51 == stage1_addr_line_mapping[10:4] ? lru_81 : _GEN_83; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_85 = 7'h52 == stage1_addr_line_mapping[10:4] ? lru_82 : _GEN_84; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_86 = 7'h53 == stage1_addr_line_mapping[10:4] ? lru_83 : _GEN_85; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_87 = 7'h54 == stage1_addr_line_mapping[10:4] ? lru_84 : _GEN_86; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_88 = 7'h55 == stage1_addr_line_mapping[10:4] ? lru_85 : _GEN_87; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_89 = 7'h56 == stage1_addr_line_mapping[10:4] ? lru_86 : _GEN_88; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_90 = 7'h57 == stage1_addr_line_mapping[10:4] ? lru_87 : _GEN_89; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_91 = 7'h58 == stage1_addr_line_mapping[10:4] ? lru_88 : _GEN_90; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_92 = 7'h59 == stage1_addr_line_mapping[10:4] ? lru_89 : _GEN_91; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_93 = 7'h5a == stage1_addr_line_mapping[10:4] ? lru_90 : _GEN_92; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_94 = 7'h5b == stage1_addr_line_mapping[10:4] ? lru_91 : _GEN_93; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_95 = 7'h5c == stage1_addr_line_mapping[10:4] ? lru_92 : _GEN_94; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_96 = 7'h5d == stage1_addr_line_mapping[10:4] ? lru_93 : _GEN_95; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_97 = 7'h5e == stage1_addr_line_mapping[10:4] ? lru_94 : _GEN_96; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_98 = 7'h5f == stage1_addr_line_mapping[10:4] ? lru_95 : _GEN_97; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_99 = 7'h60 == stage1_addr_line_mapping[10:4] ? lru_96 : _GEN_98; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_100 = 7'h61 == stage1_addr_line_mapping[10:4] ? lru_97 : _GEN_99; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_101 = 7'h62 == stage1_addr_line_mapping[10:4] ? lru_98 : _GEN_100; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_102 = 7'h63 == stage1_addr_line_mapping[10:4] ? lru_99 : _GEN_101; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_103 = 7'h64 == stage1_addr_line_mapping[10:4] ? lru_100 : _GEN_102; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_104 = 7'h65 == stage1_addr_line_mapping[10:4] ? lru_101 : _GEN_103; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_105 = 7'h66 == stage1_addr_line_mapping[10:4] ? lru_102 : _GEN_104; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_106 = 7'h67 == stage1_addr_line_mapping[10:4] ? lru_103 : _GEN_105; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_107 = 7'h68 == stage1_addr_line_mapping[10:4] ? lru_104 : _GEN_106; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_108 = 7'h69 == stage1_addr_line_mapping[10:4] ? lru_105 : _GEN_107; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_109 = 7'h6a == stage1_addr_line_mapping[10:4] ? lru_106 : _GEN_108; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_110 = 7'h6b == stage1_addr_line_mapping[10:4] ? lru_107 : _GEN_109; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_111 = 7'h6c == stage1_addr_line_mapping[10:4] ? lru_108 : _GEN_110; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_112 = 7'h6d == stage1_addr_line_mapping[10:4] ? lru_109 : _GEN_111; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_113 = 7'h6e == stage1_addr_line_mapping[10:4] ? lru_110 : _GEN_112; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_114 = 7'h6f == stage1_addr_line_mapping[10:4] ? lru_111 : _GEN_113; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_115 = 7'h70 == stage1_addr_line_mapping[10:4] ? lru_112 : _GEN_114; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_116 = 7'h71 == stage1_addr_line_mapping[10:4] ? lru_113 : _GEN_115; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_117 = 7'h72 == stage1_addr_line_mapping[10:4] ? lru_114 : _GEN_116; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_118 = 7'h73 == stage1_addr_line_mapping[10:4] ? lru_115 : _GEN_117; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_119 = 7'h74 == stage1_addr_line_mapping[10:4] ? lru_116 : _GEN_118; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_120 = 7'h75 == stage1_addr_line_mapping[10:4] ? lru_117 : _GEN_119; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_121 = 7'h76 == stage1_addr_line_mapping[10:4] ? lru_118 : _GEN_120; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_122 = 7'h77 == stage1_addr_line_mapping[10:4] ? lru_119 : _GEN_121; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_123 = 7'h78 == stage1_addr_line_mapping[10:4] ? lru_120 : _GEN_122; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_124 = 7'h79 == stage1_addr_line_mapping[10:4] ? lru_121 : _GEN_123; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_125 = 7'h7a == stage1_addr_line_mapping[10:4] ? lru_122 : _GEN_124; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_126 = 7'h7b == stage1_addr_line_mapping[10:4] ? lru_123 : _GEN_125; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_127 = 7'h7c == stage1_addr_line_mapping[10:4] ? lru_124 : _GEN_126; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_128 = 7'h7d == stage1_addr_line_mapping[10:4] ? lru_125 : _GEN_127; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_129 = 7'h7e == stage1_addr_line_mapping[10:4] ? lru_126 : _GEN_128; // @[inst_cache.scala 183:{12,12}]
  wire  _GEN_130 = 7'h7f == stage1_addr_line_mapping[10:4] ? lru_127 : _GEN_129; // @[inst_cache.scala 183:{12,12}]
  wire  _lru_T_4 = _hit_T_3 ? 1'h0 : _GEN_130; // @[inst_cache.scala 183:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[inst_cache.scala 182:12]
  wire  _lru_T_8 = ~_GEN_130; // @[inst_cache.scala 184:46]
  reg [2:0] stage2_sram_addr_reg; // @[inst_cache.scala 189:39]
  wire [2:0] _stage2_sram_addr_reg_T_2 = {stage1_addr_line_mapping[3],stage1_addr_line_mapping[1:0]}; // @[Cat.scala 31:58]
  reg  stage2_sram_req_reg; // @[inst_cache.scala 196:38]
  reg  stage2_hit0_reg; // @[inst_cache.scala 200:34]
  reg [1:0] stage2_write_en_reg; // @[inst_cache.scala 217:38]
  wire [39:0] icache_data_way0_0_rdata = icache_data_io_rdata; // @[inst_cache.scala 91:{36,36}]
  wire [39:0] icache_data_way0_1_rdata = icache_data_1_io_rdata; // @[inst_cache.scala 91:{36,36}]
  wire [39:0] _GEN_516 = stage2_sram_addr_reg[2] ? icache_data_way0_1_rdata : icache_data_way0_0_rdata; // @[inst_cache.scala 228:{25,25}]
  wire [39:0] icache_data_way1_0_rdata = icache_data_2_io_rdata; // @[inst_cache.scala 92:{36,36}]
  wire [39:0] icache_data_way1_1_rdata = icache_data_3_io_rdata; // @[inst_cache.scala 92:{36,36}]
  wire [39:0] _GEN_518 = stage2_sram_addr_reg[2] ? icache_data_way1_1_rdata : icache_data_way1_0_rdata; // @[inst_cache.scala 228:{25,25}]
  wire [39:0] hit_word_L = stage2_hit0_reg ? _GEN_516 : _GEN_518; // @[inst_cache.scala 228:25]
  reg  has_stage2_stall; // @[inst_cache.scala 230:35]
  reg [39:0] sram_rdata_L_Reg; // @[inst_cache.scala 233:35]
  wire [39:0] _access_sram_rdata_L_T_2 = _access_work_state_T_23 ? hit_word_L : 40'h0; // @[inst_cache.scala 236:84]
  wire [39:0] access_sram_rdata_L = _access_work_state_T_8 ? wait_data_L : _access_sram_rdata_L_T_2; // @[inst_cache.scala 236:35]
  wire  _icache_data_way0_0_wen_T_2 = _access_work_state_T_38 & io_port_rvalid; // @[inst_cache.scala 243:119]
  wire  _icache_data_way0_0_wen_T_6 = write_counter == 3'h0; // @[inst_cache.scala 244:69]
  wire  _icache_data_way0_0_wen_T_7 = _icache_data_way0_0_wen_T_2 & _lru_T_8 & write_counter == 3'h0; // @[inst_cache.scala 244:52]
  wire  _icache_data_way0_1_wen_T_6 = write_counter == 3'h1; // @[inst_cache.scala 244:69]
  wire  _icache_data_way0_1_wen_T_7 = _icache_data_way0_0_wen_T_2 & _lru_T_8 & write_counter == 3'h1; // @[inst_cache.scala 244:52]
  wire  _icache_data_way1_0_wen_T_7 = _icache_data_way0_0_wen_T_2 & _GEN_130 & _icache_data_way0_0_wen_T_6; // @[inst_cache.scala 246:52]
  wire  _icache_data_way1_1_wen_T_7 = _icache_data_way0_0_wen_T_2 & _GEN_130 & _icache_data_way0_1_wen_T_6; // @[inst_cache.scala 246:52]
  wire [2:0] _GEN_1287 = {{2'd0}, stage1_addr_line_mapping[3]}; // @[inst_cache.scala 266:95]
  wire [2:0] _write_counter_T_8 = write_counter + 3'h1; // @[inst_cache.scala 271:196]
  wire [21:0] _T_13 = {1'h1,stage1_addr_line_mapping[31:11]}; // @[Cat.scala 31:58]
  wire [63:0] _io_port_araddr_T_3 = {stage1_sram_phy_addr_reg[63:4],4'h0}; // @[Cat.scala 31:58]
  wire [63:0] _io_port_araddr_T_4 = _access_work_state_T_35 ? _io_port_araddr_T_3 : 64'h0; // @[inst_cache.scala 285:12]
  wire [63:0] _io_port_araddr_T_5 = _access_work_state_T ? stage1_sram_phy_addr_reg : _io_port_araddr_T_4; // @[inst_cache.scala 284:26]
  wire [1:0] _io_port_arsize_T_1 = stage1_sram_cache_reg ? 2'h3 : 2'h2; // @[inst_cache.scala 288:26]
  wire  _io_sram_write_en_T_3 = ~stage2_sram_req_reg & stage2_sram_addr_reg[1:0] != 2'h0; // @[inst_cache.scala 324:31]
  wire [1:0] _io_sram_write_en_T_5 = stage2_sram_req_reg | _io_sram_write_en_T_3 ? stage2_write_en_reg : 2'h0; // @[inst_cache.scala 323:57]
  ysyx_22040886_icache_tag icache_tag ( // @[inst_cache.scala 83:34]
    .clock(icache_tag_clock),
    .reset(icache_tag_reset),
    .io_wen(icache_tag_io_wen),
    .io_wdata(icache_tag_io_wdata),
    .io_addr(icache_tag_io_addr),
    .io_hit(icache_tag_io_hit),
    .io_valid(icache_tag_io_valid),
    .io_tag_all_flush(icache_tag_io_tag_all_flush)
  );
  ysyx_22040886_icache_tag icache_tag_1 ( // @[inst_cache.scala 85:34]
    .clock(icache_tag_1_clock),
    .reset(icache_tag_1_reset),
    .io_wen(icache_tag_1_io_wen),
    .io_wdata(icache_tag_1_io_wdata),
    .io_addr(icache_tag_1_io_addr),
    .io_hit(icache_tag_1_io_hit),
    .io_valid(icache_tag_1_io_valid),
    .io_tag_all_flush(icache_tag_1_io_tag_all_flush)
  );
  ysyx_22040886_icache_data icache_data ( // @[inst_cache.scala 91:55]
    .clock(icache_data_clock),
    .io_wen(icache_data_io_wen),
    .io_addr(icache_data_io_addr),
    .io_wdata(icache_data_io_wdata),
    .io_rdata(icache_data_io_rdata),
    .io_sram_addr(icache_data_io_sram_addr),
    .io_sram_wen(icache_data_io_sram_wen),
    .io_sram_wmask(icache_data_io_sram_wmask),
    .io_sram_wdata(icache_data_io_sram_wdata),
    .io_sram_rdata(icache_data_io_sram_rdata)
  );
  ysyx_22040886_icache_data icache_data_1 ( // @[inst_cache.scala 91:55]
    .clock(icache_data_1_clock),
    .io_wen(icache_data_1_io_wen),
    .io_addr(icache_data_1_io_addr),
    .io_wdata(icache_data_1_io_wdata),
    .io_rdata(icache_data_1_io_rdata),
    .io_sram_addr(icache_data_1_io_sram_addr),
    .io_sram_wen(icache_data_1_io_sram_wen),
    .io_sram_wmask(icache_data_1_io_sram_wmask),
    .io_sram_wdata(icache_data_1_io_sram_wdata),
    .io_sram_rdata(icache_data_1_io_sram_rdata)
  );
  ysyx_22040886_icache_data icache_data_2 ( // @[inst_cache.scala 92:55]
    .clock(icache_data_2_clock),
    .io_wen(icache_data_2_io_wen),
    .io_addr(icache_data_2_io_addr),
    .io_wdata(icache_data_2_io_wdata),
    .io_rdata(icache_data_2_io_rdata),
    .io_sram_addr(icache_data_2_io_sram_addr),
    .io_sram_wen(icache_data_2_io_sram_wen),
    .io_sram_wmask(icache_data_2_io_sram_wmask),
    .io_sram_wdata(icache_data_2_io_sram_wdata),
    .io_sram_rdata(icache_data_2_io_sram_rdata)
  );
  ysyx_22040886_icache_data icache_data_3 ( // @[inst_cache.scala 92:55]
    .clock(icache_data_3_clock),
    .io_wen(icache_data_3_io_wen),
    .io_addr(icache_data_3_io_addr),
    .io_wdata(icache_data_3_io_wdata),
    .io_rdata(icache_data_3_io_rdata),
    .io_sram_addr(icache_data_3_io_sram_addr),
    .io_sram_wen(icache_data_3_io_sram_wen),
    .io_sram_wmask(icache_data_3_io_sram_wmask),
    .io_sram_wdata(icache_data_3_io_sram_wdata),
    .io_sram_rdata(icache_data_3_io_sram_rdata)
  );
  assign io_port_araddr = _io_port_araddr_T_5[31:0]; // @[inst_cache.scala 284:20]
  assign io_port_arlen = {{7'd0}, stage1_sram_cache_reg}; // @[inst_cache.scala 287:20]
  assign io_port_arsize = {{1'd0}, _io_port_arsize_T_1}; // @[inst_cache.scala 288:20]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[inst_cache.scala 289:21]
  assign io_port_arvalid = _access_work_state_T | _access_work_state_T_35; // @[inst_cache.scala 294:59]
  assign io_stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4) & _stage2_stall_T_5; // @[inst_cache.scala 152:129]
  assign io_v_addr_for_tlb = stage1_addr_line_mapping; // @[inst_cache.scala 141:23]
  assign io_sram_write_en = io_inst_buffer_full ? 2'h0 : _io_sram_write_en_T_5; // @[inst_cache.scala 323:28]
  assign io_sram_rdata_L = _stage2_stall_T_5 & has_stage2_stall ? access_sram_rdata_L : sram_rdata_L_Reg; // @[inst_cache.scala 248:27]
  assign io_sram_0_addr = icache_data_io_sram_addr; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_0_wen = icache_data_io_sram_wen; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_0_wmask = icache_data_io_sram_wmask; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_0_wdata = icache_data_io_sram_wdata; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_1_addr = icache_data_1_io_sram_addr; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_1_wen = icache_data_1_io_sram_wen; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_1_wmask = icache_data_1_io_sram_wmask; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_1_wdata = icache_data_1_io_sram_wdata; // @[inst_cache.scala 91:{36,36}]
  assign io_sram_2_addr = icache_data_2_io_sram_addr; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_2_wen = icache_data_2_io_sram_wen; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_2_wmask = icache_data_2_io_sram_wmask; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_2_wdata = icache_data_2_io_sram_wdata; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_3_addr = icache_data_3_io_sram_addr; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_3_wen = icache_data_3_io_sram_wen; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_3_wmask = icache_data_3_io_sram_wmask; // @[inst_cache.scala 92:{36,36}]
  assign io_sram_3_wdata = icache_data_3_io_sram_wdata; // @[inst_cache.scala 92:{36,36}]
  assign icache_tag_clock = clock;
  assign icache_tag_reset = reset;
  assign icache_tag_io_wen = _stage1_finished_T_1 & _lru_T_8; // @[inst_cache.scala 272:63]
  assign icache_tag_io_wdata = _stage1_finished_T_1 ? _T_13 : 22'h0; // @[inst_cache.scala 274:30]
  assign icache_tag_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 158:25]
  assign icache_tag_io_tag_all_flush = io_tag_valid_flush; // @[inst_cache.scala 89:32]
  assign icache_tag_1_clock = clock;
  assign icache_tag_1_reset = reset;
  assign icache_tag_1_io_wen = _stage1_finished_T_1 & _GEN_130; // @[inst_cache.scala 273:63]
  assign icache_tag_1_io_wdata = _stage1_finished_T_1 ? _T_13 : 22'h0; // @[inst_cache.scala 275:30]
  assign icache_tag_1_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 159:25]
  assign icache_tag_1_io_tag_all_flush = io_tag_valid_flush; // @[inst_cache.scala 90:32]
  assign icache_data_clock = clock;
  assign icache_data_io_wen = _icache_data_way0_0_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 243:79]
  assign icache_data_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 168:34 91:36]
  assign icache_data_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_io_sram_rdata = io_sram_0_rdata; // @[inst_cache.scala 91:36 94:30]
  assign icache_data_1_clock = clock;
  assign icache_data_1_io_wen = _icache_data_way0_1_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 243:79]
  assign icache_data_1_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 168:34 91:36]
  assign icache_data_1_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_1_io_sram_rdata = io_sram_1_rdata; // @[inst_cache.scala 91:36 95:30]
  assign icache_data_2_clock = clock;
  assign icache_data_2_io_wen = _icache_data_way1_0_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 245:79]
  assign icache_data_2_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 173:34 92:36]
  assign icache_data_2_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_2_io_sram_rdata = io_sram_2_rdata; // @[inst_cache.scala 92:36 96:30]
  assign icache_data_3_clock = clock;
  assign icache_data_3_io_wen = _icache_data_way1_1_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 245:79]
  assign icache_data_3_io_addr = stage1_addr_line_mapping[31:0]; // @[inst_cache.scala 173:34 92:36]
  assign icache_data_3_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_3_io_sram_rdata = io_sram_3_rdata; // @[inst_cache.scala 92:36 97:30]
  always @(posedge clock) begin
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_0 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_0 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_0 <= ~_GEN_130;
      end else begin
        lru_0 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_1 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_1 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_1 <= ~_GEN_130;
      end else begin
        lru_1 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_2 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_2 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_2 <= ~_GEN_130;
      end else begin
        lru_2 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_3 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_3 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_3 <= ~_GEN_130;
      end else begin
        lru_3 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_4 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_4 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_4 <= ~_GEN_130;
      end else begin
        lru_4 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_5 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_5 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_5 <= ~_GEN_130;
      end else begin
        lru_5 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_6 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_6 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_6 <= ~_GEN_130;
      end else begin
        lru_6 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_7 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_7 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_7 <= ~_GEN_130;
      end else begin
        lru_7 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_8 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_8 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_8 <= ~_GEN_130;
      end else begin
        lru_8 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_9 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_9 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_9 <= ~_GEN_130;
      end else begin
        lru_9 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_10 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_10 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_10 <= ~_GEN_130;
      end else begin
        lru_10 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_11 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_11 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_11 <= ~_GEN_130;
      end else begin
        lru_11 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_12 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_12 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_12 <= ~_GEN_130;
      end else begin
        lru_12 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_13 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_13 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_13 <= ~_GEN_130;
      end else begin
        lru_13 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_14 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_14 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_14 <= ~_GEN_130;
      end else begin
        lru_14 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_15 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_15 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_15 <= ~_GEN_130;
      end else begin
        lru_15 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_16 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_16 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_16 <= ~_GEN_130;
      end else begin
        lru_16 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_17 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_17 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_17 <= ~_GEN_130;
      end else begin
        lru_17 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_18 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_18 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_18 <= ~_GEN_130;
      end else begin
        lru_18 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_19 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_19 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_19 <= ~_GEN_130;
      end else begin
        lru_19 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_20 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_20 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_20 <= ~_GEN_130;
      end else begin
        lru_20 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_21 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_21 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_21 <= ~_GEN_130;
      end else begin
        lru_21 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_22 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_22 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_22 <= ~_GEN_130;
      end else begin
        lru_22 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_23 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_23 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_23 <= ~_GEN_130;
      end else begin
        lru_23 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_24 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_24 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_24 <= ~_GEN_130;
      end else begin
        lru_24 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_25 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_25 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_25 <= ~_GEN_130;
      end else begin
        lru_25 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_26 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_26 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_26 <= ~_GEN_130;
      end else begin
        lru_26 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_27 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_27 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_27 <= ~_GEN_130;
      end else begin
        lru_27 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_28 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_28 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_28 <= ~_GEN_130;
      end else begin
        lru_28 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_29 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_29 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_29 <= ~_GEN_130;
      end else begin
        lru_29 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_30 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_30 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_30 <= ~_GEN_130;
      end else begin
        lru_30 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_31 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_31 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_31 <= ~_GEN_130;
      end else begin
        lru_31 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_32 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_32 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_32 <= ~_GEN_130;
      end else begin
        lru_32 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_33 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_33 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_33 <= ~_GEN_130;
      end else begin
        lru_33 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_34 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_34 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_34 <= ~_GEN_130;
      end else begin
        lru_34 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_35 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_35 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_35 <= ~_GEN_130;
      end else begin
        lru_35 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_36 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_36 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_36 <= ~_GEN_130;
      end else begin
        lru_36 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_37 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_37 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_37 <= ~_GEN_130;
      end else begin
        lru_37 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_38 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_38 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_38 <= ~_GEN_130;
      end else begin
        lru_38 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_39 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_39 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_39 <= ~_GEN_130;
      end else begin
        lru_39 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_40 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_40 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_40 <= ~_GEN_130;
      end else begin
        lru_40 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_41 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_41 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_41 <= ~_GEN_130;
      end else begin
        lru_41 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_42 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_42 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_42 <= ~_GEN_130;
      end else begin
        lru_42 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_43 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_43 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_43 <= ~_GEN_130;
      end else begin
        lru_43 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_44 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_44 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_44 <= ~_GEN_130;
      end else begin
        lru_44 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_45 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_45 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_45 <= ~_GEN_130;
      end else begin
        lru_45 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_46 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_46 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_46 <= ~_GEN_130;
      end else begin
        lru_46 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_47 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_47 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_47 <= ~_GEN_130;
      end else begin
        lru_47 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_48 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_48 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_48 <= ~_GEN_130;
      end else begin
        lru_48 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_49 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_49 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_49 <= ~_GEN_130;
      end else begin
        lru_49 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_50 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_50 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_50 <= ~_GEN_130;
      end else begin
        lru_50 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_51 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_51 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_51 <= ~_GEN_130;
      end else begin
        lru_51 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_52 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_52 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_52 <= ~_GEN_130;
      end else begin
        lru_52 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_53 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_53 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_53 <= ~_GEN_130;
      end else begin
        lru_53 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_54 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_54 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_54 <= ~_GEN_130;
      end else begin
        lru_54 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_55 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_55 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_55 <= ~_GEN_130;
      end else begin
        lru_55 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_56 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_56 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_56 <= ~_GEN_130;
      end else begin
        lru_56 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_57 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_57 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_57 <= ~_GEN_130;
      end else begin
        lru_57 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_58 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_58 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_58 <= ~_GEN_130;
      end else begin
        lru_58 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_59 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_59 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_59 <= ~_GEN_130;
      end else begin
        lru_59 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_60 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_60 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_60 <= ~_GEN_130;
      end else begin
        lru_60 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_61 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_61 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_61 <= ~_GEN_130;
      end else begin
        lru_61 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_62 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_62 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_62 <= ~_GEN_130;
      end else begin
        lru_62 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_63 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_63 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_63 <= ~_GEN_130;
      end else begin
        lru_63 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_64 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_64 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_64 <= ~_GEN_130;
      end else begin
        lru_64 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_65 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_65 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_65 <= ~_GEN_130;
      end else begin
        lru_65 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_66 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_66 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_66 <= ~_GEN_130;
      end else begin
        lru_66 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_67 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_67 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_67 <= ~_GEN_130;
      end else begin
        lru_67 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_68 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_68 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_68 <= ~_GEN_130;
      end else begin
        lru_68 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_69 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_69 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_69 <= ~_GEN_130;
      end else begin
        lru_69 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_70 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_70 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_70 <= ~_GEN_130;
      end else begin
        lru_70 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_71 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_71 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_71 <= ~_GEN_130;
      end else begin
        lru_71 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_72 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_72 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_72 <= ~_GEN_130;
      end else begin
        lru_72 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_73 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_73 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_73 <= ~_GEN_130;
      end else begin
        lru_73 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_74 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_74 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_74 <= ~_GEN_130;
      end else begin
        lru_74 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_75 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_75 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_75 <= ~_GEN_130;
      end else begin
        lru_75 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_76 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_76 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_76 <= ~_GEN_130;
      end else begin
        lru_76 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_77 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_77 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_77 <= ~_GEN_130;
      end else begin
        lru_77 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_78 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_78 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_78 <= ~_GEN_130;
      end else begin
        lru_78 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_79 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_79 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_79 <= ~_GEN_130;
      end else begin
        lru_79 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_80 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_80 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_80 <= ~_GEN_130;
      end else begin
        lru_80 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_81 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_81 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_81 <= ~_GEN_130;
      end else begin
        lru_81 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_82 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_82 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_82 <= ~_GEN_130;
      end else begin
        lru_82 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_83 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_83 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_83 <= ~_GEN_130;
      end else begin
        lru_83 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_84 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_84 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_84 <= ~_GEN_130;
      end else begin
        lru_84 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_85 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_85 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_85 <= ~_GEN_130;
      end else begin
        lru_85 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_86 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_86 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_86 <= ~_GEN_130;
      end else begin
        lru_86 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_87 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_87 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_87 <= ~_GEN_130;
      end else begin
        lru_87 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_88 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_88 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_88 <= ~_GEN_130;
      end else begin
        lru_88 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_89 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_89 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_89 <= ~_GEN_130;
      end else begin
        lru_89 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_90 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_90 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_90 <= ~_GEN_130;
      end else begin
        lru_90 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_91 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_91 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_91 <= ~_GEN_130;
      end else begin
        lru_91 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_92 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_92 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_92 <= ~_GEN_130;
      end else begin
        lru_92 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_93 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_93 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_93 <= ~_GEN_130;
      end else begin
        lru_93 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_94 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_94 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_94 <= ~_GEN_130;
      end else begin
        lru_94 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_95 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_95 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_95 <= ~_GEN_130;
      end else begin
        lru_95 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_96 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_96 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_96 <= ~_GEN_130;
      end else begin
        lru_96 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_97 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_97 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_97 <= ~_GEN_130;
      end else begin
        lru_97 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_98 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_98 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_98 <= ~_GEN_130;
      end else begin
        lru_98 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_99 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_99 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_99 <= ~_GEN_130;
      end else begin
        lru_99 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_100 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_100 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_100 <= ~_GEN_130;
      end else begin
        lru_100 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_101 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_101 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_101 <= ~_GEN_130;
      end else begin
        lru_101 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_102 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_102 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_102 <= ~_GEN_130;
      end else begin
        lru_102 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_103 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_103 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_103 <= ~_GEN_130;
      end else begin
        lru_103 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_104 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_104 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_104 <= ~_GEN_130;
      end else begin
        lru_104 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_105 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_105 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_105 <= ~_GEN_130;
      end else begin
        lru_105 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_106 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_106 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_106 <= ~_GEN_130;
      end else begin
        lru_106 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_107 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_107 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_107 <= ~_GEN_130;
      end else begin
        lru_107 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_108 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_108 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_108 <= ~_GEN_130;
      end else begin
        lru_108 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_109 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_109 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_109 <= ~_GEN_130;
      end else begin
        lru_109 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_110 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_110 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_110 <= ~_GEN_130;
      end else begin
        lru_110 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_111 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_111 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_111 <= ~_GEN_130;
      end else begin
        lru_111 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_112 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_112 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_112 <= ~_GEN_130;
      end else begin
        lru_112 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_113 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_113 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_113 <= ~_GEN_130;
      end else begin
        lru_113 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_114 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_114 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_114 <= ~_GEN_130;
      end else begin
        lru_114 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_115 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_115 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_115 <= ~_GEN_130;
      end else begin
        lru_115 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_116 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_116 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_116 <= ~_GEN_130;
      end else begin
        lru_116 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_117 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_117 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_117 <= ~_GEN_130;
      end else begin
        lru_117 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_118 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_118 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_118 <= ~_GEN_130;
      end else begin
        lru_118 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_119 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_119 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_119 <= ~_GEN_130;
      end else begin
        lru_119 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_120 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_120 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_120 <= ~_GEN_130;
      end else begin
        lru_120 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_121 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_121 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_121 <= ~_GEN_130;
      end else begin
        lru_121 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_122 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_122 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_122 <= ~_GEN_130;
      end else begin
        lru_122 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_123 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_123 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_123 <= ~_GEN_130;
      end else begin
        lru_123 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_124 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_124 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_124 <= ~_GEN_130;
      end else begin
        lru_124 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_125 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_125 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_125 <= ~_GEN_130;
      end else begin
        lru_125 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_126 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_126 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_126 <= ~_GEN_130;
      end else begin
        lru_126 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 76:22]
      lru_127 <= 1'h0; // @[inst_cache.scala 76:22]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 181:37]
      if (_stage2_stall_T) begin // @[inst_cache.scala 181:43]
        lru_127 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin // @[inst_cache.scala 184:12]
        lru_127 <= ~_GEN_130;
      end else begin
        lru_127 <= _GEN_130;
      end
    end
    if (reset) begin // @[inst_cache.scala 108:29]
      work_state <= 4'h1; // @[inst_cache.scala 108:29]
    end else if (work_state == 4'h2 & io_port_arready) begin // @[inst_cache.scala 251:30]
      work_state <= 4'h3;
    end else if (_stage1_finished_T_2) begin // @[inst_cache.scala 252:12]
      work_state <= {{1'd0}, _access_work_state_T_7};
    end else if (work_state == 4'h4) begin // @[inst_cache.scala 253:12]
      work_state <= {{1'd0}, _access_work_state_T_22};
    end else begin
      work_state <= _access_work_state_T_47;
    end
    if (reset) begin // @[inst_cache.scala 110:33]
      write_counter <= 3'h0; // @[inst_cache.scala 110:33]
    end else if (_access_work_state_T_38 | _stage1_finished_T_2) begin // @[inst_cache.scala 271:26]
      if (io_port_rvalid & io_port_rlast) begin // @[inst_cache.scala 271:106]
        write_counter <= 3'h0;
      end else if (io_port_rvalid) begin // @[inst_cache.scala 271:160]
        write_counter <= _write_counter_T_8;
      end
    end
    if (reset) begin // @[inst_cache.scala 111:31]
      wait_data_L <= 40'h0; // @[inst_cache.scala 111:31]
    end else if (_stage1_finished_T_2 & io_port_rvalid & _icache_data_way0_0_wen_T_6) begin // @[inst_cache.scala 265:23]
      wait_data_L <= decoder_inst_data;
    end else if (_icache_data_way0_0_wen_T_2 & write_counter == _GEN_1287) begin // @[inst_cache.scala 266:13]
      wait_data_L <= decoder_inst_data;
    end
    if (reset) begin // @[inst_cache.scala 122:35]
      stage1_stall_reg <= 1'h0; // @[inst_cache.scala 122:35]
    end else begin
      stage1_stall_reg <= io_sram_req; // @[inst_cache.scala 123:22]
    end
    if (reset) begin // @[Reg.scala 28:20]
      stage1_addr_line_mapping <= 64'h0; // @[Reg.scala 28:20]
    end else if (io_sram_req) begin // @[Reg.scala 29:18]
      if (stage1_flush) begin // @[inst_cache.scala 125:45]
        stage1_addr_line_mapping <= 64'h0;
      end else begin
        stage1_addr_line_mapping <= io_sram_addr;
      end
    end
    if (reset) begin // @[inst_cache.scala 126:43]
      stage1_sram_phy_addr_reg <= 64'h0; // @[inst_cache.scala 126:43]
    end else if (stage1_stall_reg) begin // @[inst_cache.scala 144:38]
      stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
    end
    if (reset) begin // @[Reg.scala 28:20]
      stage1_sram_cache_reg <= 1'h0; // @[Reg.scala 28:20]
    end else if (io_sram_req) begin // @[Reg.scala 29:18]
      if (stage1_flush) begin // @[inst_cache.scala 127:46]
        stage1_sram_cache_reg <= 1'h0;
      end else begin
        stage1_sram_cache_reg <= io_sram_cache;
      end
    end
    if (reset) begin // @[Reg.scala 28:20]
      stage1_sram_req_reg <= 1'h0; // @[Reg.scala 28:20]
    end else if (_stage1_sram_req_reg_T_1) begin // @[Reg.scala 29:18]
      if (stage1_flush) begin // @[inst_cache.scala 128:44]
        stage1_sram_req_reg <= 1'h0;
      end else begin
        stage1_sram_req_reg <= io_inst_ready_to_use;
      end
    end
    if (reset) begin // @[inst_cache.scala 131:34]
      stage1_finished <= 1'h0; // @[inst_cache.scala 131:34]
    end else if (io_sram_req) begin // @[inst_cache.scala 147:27]
      stage1_finished <= 1'h0;
    end else begin
      stage1_finished <= work_state == 4'h7 | work_state == 4'h3;
    end
    if (reset) begin // @[inst_cache.scala 189:39]
      stage2_sram_addr_reg <= 3'h0; // @[inst_cache.scala 189:39]
    end else if (io_stage2_flush) begin // @[inst_cache.scala 191:33]
      stage2_sram_addr_reg <= 3'h0;
    end else if (stage2_stall) begin // @[inst_cache.scala 191:54]
      stage2_sram_addr_reg <= _stage2_sram_addr_reg_T_2;
    end
    if (reset) begin // @[inst_cache.scala 196:38]
      stage2_sram_req_reg <= 1'h0; // @[inst_cache.scala 196:38]
    end else if (io_stage2_flush) begin // @[inst_cache.scala 197:31]
      stage2_sram_req_reg <= 1'h0;
    end else if (stage2_stall) begin // @[inst_cache.scala 197:52]
      stage2_sram_req_reg <= stage1_sram_req_reg;
    end else begin
      stage2_sram_req_reg <= io_sram_write_en == 2'h0 & stage2_sram_req_reg;
    end
    if (reset) begin // @[inst_cache.scala 200:34]
      stage2_hit0_reg <= 1'h0; // @[inst_cache.scala 200:34]
    end else if (io_stage2_flush) begin // @[inst_cache.scala 201:27]
      stage2_hit0_reg <= 1'h0;
    end else if (stage2_stall) begin // @[inst_cache.scala 201:48]
      stage2_hit0_reg <= _hit_T_2;
    end
    if (reset) begin // @[inst_cache.scala 217:38]
      stage2_write_en_reg <= 2'h0; // @[inst_cache.scala 217:38]
    end else if (io_stage1_valid_flush) begin // @[inst_cache.scala 219:31]
      stage2_write_en_reg <= 2'h0;
    end else if (stage2_stall) begin // @[inst_cache.scala 219:61]
      stage2_write_en_reg <= 2'h1;
    end
    if (reset) begin // @[inst_cache.scala 230:35]
      has_stage2_stall <= 1'h0; // @[inst_cache.scala 230:35]
    end else begin
      has_stage2_stall <= stage2_stall; // @[inst_cache.scala 231:22]
    end
    if (reset) begin // @[inst_cache.scala 233:35]
      sram_rdata_L_Reg <= 40'h0; // @[inst_cache.scala 233:35]
    end else if (has_stage2_stall) begin // @[inst_cache.scala 239:28]
      if (_access_work_state_T_8) begin // @[inst_cache.scala 236:35]
        sram_rdata_L_Reg <= wait_data_L;
      end else if (_access_work_state_T_23) begin // @[inst_cache.scala 236:84]
        sram_rdata_L_Reg <= hit_word_L;
      end else begin
        sram_rdata_L_Reg <= 40'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lru_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lru_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  work_state = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  write_counter = _RAND_129[2:0];
  _RAND_130 = {2{`RANDOM}};
  wait_data_L = _RAND_130[39:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_131[0:0];
  _RAND_132 = {2{`RANDOM}};
  stage1_addr_line_mapping = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_133[63:0];
  _RAND_134 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  stage1_finished = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  stage2_sram_addr_reg = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  stage2_sram_req_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  stage2_write_en_reg = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  has_stage2_stall = _RAND_141[0:0];
  _RAND_142 = {2{`RANDOM}};
  sram_rdata_L_Reg = _RAND_142[39:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_dcache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [21:0] io_wdata,
  input  [31:0] io_raddr,
  input  [31:0] io_waddr,
  output        io_hit,
  output        io_valid,
  output [20:0] io_tag,
  output        io_w_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] tag_regs0_0; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_1; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_2; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_3; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_4; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_5; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_6; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_7; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_8; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_9; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_10; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_11; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_12; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_13; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_14; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_15; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_16; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_17; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_18; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_19; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_20; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_21; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_22; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_23; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_24; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_25; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_26; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_27; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_28; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_29; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_30; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_31; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_32; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_33; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_34; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_35; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_36; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_37; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_38; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_39; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_40; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_41; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_42; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_43; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_44; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_45; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_46; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_47; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_48; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_49; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_50; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_51; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_52; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_53; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_54; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_55; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_56; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_57; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_58; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_59; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_60; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_61; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_62; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs0_63; // @[dcache_tag.scala 23:28]
  reg [21:0] tag_regs1_0; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_1; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_2; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_3; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_4; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_5; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_6; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_7; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_8; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_9; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_10; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_11; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_12; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_13; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_14; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_15; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_16; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_17; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_18; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_19; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_20; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_21; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_22; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_23; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_24; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_25; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_26; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_27; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_28; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_29; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_30; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_31; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_32; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_33; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_34; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_35; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_36; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_37; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_38; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_39; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_40; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_41; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_42; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_43; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_44; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_45; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_46; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_47; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_48; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_49; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_50; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_51; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_52; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_53; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_54; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_55; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_56; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_57; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_58; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_59; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_60; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_61; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_62; // @[dcache_tag.scala 24:28]
  reg [21:0] tag_regs1_63; // @[dcache_tag.scala 24:28]
  wire [21:0] _GEN_1 = 6'h1 == io_waddr[10:5] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_2 = 6'h2 == io_waddr[10:5] ? tag_regs0_2 : _GEN_1; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_3 = 6'h3 == io_waddr[10:5] ? tag_regs0_3 : _GEN_2; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_4 = 6'h4 == io_waddr[10:5] ? tag_regs0_4 : _GEN_3; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_5 = 6'h5 == io_waddr[10:5] ? tag_regs0_5 : _GEN_4; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_6 = 6'h6 == io_waddr[10:5] ? tag_regs0_6 : _GEN_5; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_7 = 6'h7 == io_waddr[10:5] ? tag_regs0_7 : _GEN_6; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_8 = 6'h8 == io_waddr[10:5] ? tag_regs0_8 : _GEN_7; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_9 = 6'h9 == io_waddr[10:5] ? tag_regs0_9 : _GEN_8; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_10 = 6'ha == io_waddr[10:5] ? tag_regs0_10 : _GEN_9; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_11 = 6'hb == io_waddr[10:5] ? tag_regs0_11 : _GEN_10; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_12 = 6'hc == io_waddr[10:5] ? tag_regs0_12 : _GEN_11; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_13 = 6'hd == io_waddr[10:5] ? tag_regs0_13 : _GEN_12; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_14 = 6'he == io_waddr[10:5] ? tag_regs0_14 : _GEN_13; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_15 = 6'hf == io_waddr[10:5] ? tag_regs0_15 : _GEN_14; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_16 = 6'h10 == io_waddr[10:5] ? tag_regs0_16 : _GEN_15; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_17 = 6'h11 == io_waddr[10:5] ? tag_regs0_17 : _GEN_16; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_18 = 6'h12 == io_waddr[10:5] ? tag_regs0_18 : _GEN_17; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_19 = 6'h13 == io_waddr[10:5] ? tag_regs0_19 : _GEN_18; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_20 = 6'h14 == io_waddr[10:5] ? tag_regs0_20 : _GEN_19; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_21 = 6'h15 == io_waddr[10:5] ? tag_regs0_21 : _GEN_20; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_22 = 6'h16 == io_waddr[10:5] ? tag_regs0_22 : _GEN_21; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_23 = 6'h17 == io_waddr[10:5] ? tag_regs0_23 : _GEN_22; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_24 = 6'h18 == io_waddr[10:5] ? tag_regs0_24 : _GEN_23; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_25 = 6'h19 == io_waddr[10:5] ? tag_regs0_25 : _GEN_24; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_26 = 6'h1a == io_waddr[10:5] ? tag_regs0_26 : _GEN_25; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_27 = 6'h1b == io_waddr[10:5] ? tag_regs0_27 : _GEN_26; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_28 = 6'h1c == io_waddr[10:5] ? tag_regs0_28 : _GEN_27; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_29 = 6'h1d == io_waddr[10:5] ? tag_regs0_29 : _GEN_28; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_30 = 6'h1e == io_waddr[10:5] ? tag_regs0_30 : _GEN_29; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_31 = 6'h1f == io_waddr[10:5] ? tag_regs0_31 : _GEN_30; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_32 = 6'h20 == io_waddr[10:5] ? tag_regs0_32 : _GEN_31; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_33 = 6'h21 == io_waddr[10:5] ? tag_regs0_33 : _GEN_32; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_34 = 6'h22 == io_waddr[10:5] ? tag_regs0_34 : _GEN_33; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_35 = 6'h23 == io_waddr[10:5] ? tag_regs0_35 : _GEN_34; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_36 = 6'h24 == io_waddr[10:5] ? tag_regs0_36 : _GEN_35; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_37 = 6'h25 == io_waddr[10:5] ? tag_regs0_37 : _GEN_36; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_38 = 6'h26 == io_waddr[10:5] ? tag_regs0_38 : _GEN_37; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_39 = 6'h27 == io_waddr[10:5] ? tag_regs0_39 : _GEN_38; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_40 = 6'h28 == io_waddr[10:5] ? tag_regs0_40 : _GEN_39; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_41 = 6'h29 == io_waddr[10:5] ? tag_regs0_41 : _GEN_40; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_42 = 6'h2a == io_waddr[10:5] ? tag_regs0_42 : _GEN_41; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_43 = 6'h2b == io_waddr[10:5] ? tag_regs0_43 : _GEN_42; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_44 = 6'h2c == io_waddr[10:5] ? tag_regs0_44 : _GEN_43; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_45 = 6'h2d == io_waddr[10:5] ? tag_regs0_45 : _GEN_44; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_46 = 6'h2e == io_waddr[10:5] ? tag_regs0_46 : _GEN_45; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_47 = 6'h2f == io_waddr[10:5] ? tag_regs0_47 : _GEN_46; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_48 = 6'h30 == io_waddr[10:5] ? tag_regs0_48 : _GEN_47; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_49 = 6'h31 == io_waddr[10:5] ? tag_regs0_49 : _GEN_48; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_50 = 6'h32 == io_waddr[10:5] ? tag_regs0_50 : _GEN_49; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_51 = 6'h33 == io_waddr[10:5] ? tag_regs0_51 : _GEN_50; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_52 = 6'h34 == io_waddr[10:5] ? tag_regs0_52 : _GEN_51; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_53 = 6'h35 == io_waddr[10:5] ? tag_regs0_53 : _GEN_52; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_54 = 6'h36 == io_waddr[10:5] ? tag_regs0_54 : _GEN_53; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_55 = 6'h37 == io_waddr[10:5] ? tag_regs0_55 : _GEN_54; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_56 = 6'h38 == io_waddr[10:5] ? tag_regs0_56 : _GEN_55; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_57 = 6'h39 == io_waddr[10:5] ? tag_regs0_57 : _GEN_56; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_58 = 6'h3a == io_waddr[10:5] ? tag_regs0_58 : _GEN_57; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_59 = 6'h3b == io_waddr[10:5] ? tag_regs0_59 : _GEN_58; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_60 = 6'h3c == io_waddr[10:5] ? tag_regs0_60 : _GEN_59; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_61 = 6'h3d == io_waddr[10:5] ? tag_regs0_61 : _GEN_60; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_62 = 6'h3e == io_waddr[10:5] ? tag_regs0_62 : _GEN_61; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_63 = 6'h3f == io_waddr[10:5] ? tag_regs0_63 : _GEN_62; // @[dcache_tag.scala 27:{37,37}]
  wire [21:0] _GEN_129 = 6'h1 == io_waddr[10:5] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_130 = 6'h2 == io_waddr[10:5] ? tag_regs1_2 : _GEN_129; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_131 = 6'h3 == io_waddr[10:5] ? tag_regs1_3 : _GEN_130; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_132 = 6'h4 == io_waddr[10:5] ? tag_regs1_4 : _GEN_131; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_133 = 6'h5 == io_waddr[10:5] ? tag_regs1_5 : _GEN_132; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_134 = 6'h6 == io_waddr[10:5] ? tag_regs1_6 : _GEN_133; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_135 = 6'h7 == io_waddr[10:5] ? tag_regs1_7 : _GEN_134; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_136 = 6'h8 == io_waddr[10:5] ? tag_regs1_8 : _GEN_135; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_137 = 6'h9 == io_waddr[10:5] ? tag_regs1_9 : _GEN_136; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_138 = 6'ha == io_waddr[10:5] ? tag_regs1_10 : _GEN_137; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_139 = 6'hb == io_waddr[10:5] ? tag_regs1_11 : _GEN_138; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_140 = 6'hc == io_waddr[10:5] ? tag_regs1_12 : _GEN_139; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_141 = 6'hd == io_waddr[10:5] ? tag_regs1_13 : _GEN_140; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_142 = 6'he == io_waddr[10:5] ? tag_regs1_14 : _GEN_141; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_143 = 6'hf == io_waddr[10:5] ? tag_regs1_15 : _GEN_142; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_144 = 6'h10 == io_waddr[10:5] ? tag_regs1_16 : _GEN_143; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_145 = 6'h11 == io_waddr[10:5] ? tag_regs1_17 : _GEN_144; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_146 = 6'h12 == io_waddr[10:5] ? tag_regs1_18 : _GEN_145; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_147 = 6'h13 == io_waddr[10:5] ? tag_regs1_19 : _GEN_146; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_148 = 6'h14 == io_waddr[10:5] ? tag_regs1_20 : _GEN_147; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_149 = 6'h15 == io_waddr[10:5] ? tag_regs1_21 : _GEN_148; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_150 = 6'h16 == io_waddr[10:5] ? tag_regs1_22 : _GEN_149; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_151 = 6'h17 == io_waddr[10:5] ? tag_regs1_23 : _GEN_150; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_152 = 6'h18 == io_waddr[10:5] ? tag_regs1_24 : _GEN_151; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_153 = 6'h19 == io_waddr[10:5] ? tag_regs1_25 : _GEN_152; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_154 = 6'h1a == io_waddr[10:5] ? tag_regs1_26 : _GEN_153; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_155 = 6'h1b == io_waddr[10:5] ? tag_regs1_27 : _GEN_154; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_156 = 6'h1c == io_waddr[10:5] ? tag_regs1_28 : _GEN_155; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_157 = 6'h1d == io_waddr[10:5] ? tag_regs1_29 : _GEN_156; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_158 = 6'h1e == io_waddr[10:5] ? tag_regs1_30 : _GEN_157; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_159 = 6'h1f == io_waddr[10:5] ? tag_regs1_31 : _GEN_158; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_160 = 6'h20 == io_waddr[10:5] ? tag_regs1_32 : _GEN_159; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_161 = 6'h21 == io_waddr[10:5] ? tag_regs1_33 : _GEN_160; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_162 = 6'h22 == io_waddr[10:5] ? tag_regs1_34 : _GEN_161; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_163 = 6'h23 == io_waddr[10:5] ? tag_regs1_35 : _GEN_162; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_164 = 6'h24 == io_waddr[10:5] ? tag_regs1_36 : _GEN_163; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_165 = 6'h25 == io_waddr[10:5] ? tag_regs1_37 : _GEN_164; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_166 = 6'h26 == io_waddr[10:5] ? tag_regs1_38 : _GEN_165; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_167 = 6'h27 == io_waddr[10:5] ? tag_regs1_39 : _GEN_166; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_168 = 6'h28 == io_waddr[10:5] ? tag_regs1_40 : _GEN_167; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_169 = 6'h29 == io_waddr[10:5] ? tag_regs1_41 : _GEN_168; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_170 = 6'h2a == io_waddr[10:5] ? tag_regs1_42 : _GEN_169; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_171 = 6'h2b == io_waddr[10:5] ? tag_regs1_43 : _GEN_170; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_172 = 6'h2c == io_waddr[10:5] ? tag_regs1_44 : _GEN_171; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_173 = 6'h2d == io_waddr[10:5] ? tag_regs1_45 : _GEN_172; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_174 = 6'h2e == io_waddr[10:5] ? tag_regs1_46 : _GEN_173; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_175 = 6'h2f == io_waddr[10:5] ? tag_regs1_47 : _GEN_174; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_176 = 6'h30 == io_waddr[10:5] ? tag_regs1_48 : _GEN_175; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_177 = 6'h31 == io_waddr[10:5] ? tag_regs1_49 : _GEN_176; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_178 = 6'h32 == io_waddr[10:5] ? tag_regs1_50 : _GEN_177; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_179 = 6'h33 == io_waddr[10:5] ? tag_regs1_51 : _GEN_178; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_180 = 6'h34 == io_waddr[10:5] ? tag_regs1_52 : _GEN_179; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_181 = 6'h35 == io_waddr[10:5] ? tag_regs1_53 : _GEN_180; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_182 = 6'h36 == io_waddr[10:5] ? tag_regs1_54 : _GEN_181; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_183 = 6'h37 == io_waddr[10:5] ? tag_regs1_55 : _GEN_182; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_184 = 6'h38 == io_waddr[10:5] ? tag_regs1_56 : _GEN_183; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_185 = 6'h39 == io_waddr[10:5] ? tag_regs1_57 : _GEN_184; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_186 = 6'h3a == io_waddr[10:5] ? tag_regs1_58 : _GEN_185; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_187 = 6'h3b == io_waddr[10:5] ? tag_regs1_59 : _GEN_186; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_188 = 6'h3c == io_waddr[10:5] ? tag_regs1_60 : _GEN_187; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_189 = 6'h3d == io_waddr[10:5] ? tag_regs1_61 : _GEN_188; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_190 = 6'h3e == io_waddr[10:5] ? tag_regs1_62 : _GEN_189; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_191 = 6'h3f == io_waddr[10:5] ? tag_regs1_63 : _GEN_190; // @[dcache_tag.scala 28:{37,37}]
  wire [21:0] _GEN_385 = 6'h1 == io_raddr[10:5] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_386 = 6'h2 == io_raddr[10:5] ? tag_regs1_2 : _GEN_385; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_387 = 6'h3 == io_raddr[10:5] ? tag_regs1_3 : _GEN_386; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_388 = 6'h4 == io_raddr[10:5] ? tag_regs1_4 : _GEN_387; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_389 = 6'h5 == io_raddr[10:5] ? tag_regs1_5 : _GEN_388; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_390 = 6'h6 == io_raddr[10:5] ? tag_regs1_6 : _GEN_389; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_391 = 6'h7 == io_raddr[10:5] ? tag_regs1_7 : _GEN_390; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_392 = 6'h8 == io_raddr[10:5] ? tag_regs1_8 : _GEN_391; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_393 = 6'h9 == io_raddr[10:5] ? tag_regs1_9 : _GEN_392; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_394 = 6'ha == io_raddr[10:5] ? tag_regs1_10 : _GEN_393; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_395 = 6'hb == io_raddr[10:5] ? tag_regs1_11 : _GEN_394; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_396 = 6'hc == io_raddr[10:5] ? tag_regs1_12 : _GEN_395; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_397 = 6'hd == io_raddr[10:5] ? tag_regs1_13 : _GEN_396; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_398 = 6'he == io_raddr[10:5] ? tag_regs1_14 : _GEN_397; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_399 = 6'hf == io_raddr[10:5] ? tag_regs1_15 : _GEN_398; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_400 = 6'h10 == io_raddr[10:5] ? tag_regs1_16 : _GEN_399; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_401 = 6'h11 == io_raddr[10:5] ? tag_regs1_17 : _GEN_400; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_402 = 6'h12 == io_raddr[10:5] ? tag_regs1_18 : _GEN_401; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_403 = 6'h13 == io_raddr[10:5] ? tag_regs1_19 : _GEN_402; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_404 = 6'h14 == io_raddr[10:5] ? tag_regs1_20 : _GEN_403; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_405 = 6'h15 == io_raddr[10:5] ? tag_regs1_21 : _GEN_404; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_406 = 6'h16 == io_raddr[10:5] ? tag_regs1_22 : _GEN_405; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_407 = 6'h17 == io_raddr[10:5] ? tag_regs1_23 : _GEN_406; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_408 = 6'h18 == io_raddr[10:5] ? tag_regs1_24 : _GEN_407; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_409 = 6'h19 == io_raddr[10:5] ? tag_regs1_25 : _GEN_408; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_410 = 6'h1a == io_raddr[10:5] ? tag_regs1_26 : _GEN_409; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_411 = 6'h1b == io_raddr[10:5] ? tag_regs1_27 : _GEN_410; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_412 = 6'h1c == io_raddr[10:5] ? tag_regs1_28 : _GEN_411; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_413 = 6'h1d == io_raddr[10:5] ? tag_regs1_29 : _GEN_412; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_414 = 6'h1e == io_raddr[10:5] ? tag_regs1_30 : _GEN_413; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_415 = 6'h1f == io_raddr[10:5] ? tag_regs1_31 : _GEN_414; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_416 = 6'h20 == io_raddr[10:5] ? tag_regs1_32 : _GEN_415; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_417 = 6'h21 == io_raddr[10:5] ? tag_regs1_33 : _GEN_416; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_418 = 6'h22 == io_raddr[10:5] ? tag_regs1_34 : _GEN_417; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_419 = 6'h23 == io_raddr[10:5] ? tag_regs1_35 : _GEN_418; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_420 = 6'h24 == io_raddr[10:5] ? tag_regs1_36 : _GEN_419; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_421 = 6'h25 == io_raddr[10:5] ? tag_regs1_37 : _GEN_420; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_422 = 6'h26 == io_raddr[10:5] ? tag_regs1_38 : _GEN_421; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_423 = 6'h27 == io_raddr[10:5] ? tag_regs1_39 : _GEN_422; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_424 = 6'h28 == io_raddr[10:5] ? tag_regs1_40 : _GEN_423; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_425 = 6'h29 == io_raddr[10:5] ? tag_regs1_41 : _GEN_424; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_426 = 6'h2a == io_raddr[10:5] ? tag_regs1_42 : _GEN_425; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_427 = 6'h2b == io_raddr[10:5] ? tag_regs1_43 : _GEN_426; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_428 = 6'h2c == io_raddr[10:5] ? tag_regs1_44 : _GEN_427; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_429 = 6'h2d == io_raddr[10:5] ? tag_regs1_45 : _GEN_428; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_430 = 6'h2e == io_raddr[10:5] ? tag_regs1_46 : _GEN_429; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_431 = 6'h2f == io_raddr[10:5] ? tag_regs1_47 : _GEN_430; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_432 = 6'h30 == io_raddr[10:5] ? tag_regs1_48 : _GEN_431; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_433 = 6'h31 == io_raddr[10:5] ? tag_regs1_49 : _GEN_432; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_434 = 6'h32 == io_raddr[10:5] ? tag_regs1_50 : _GEN_433; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_435 = 6'h33 == io_raddr[10:5] ? tag_regs1_51 : _GEN_434; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_436 = 6'h34 == io_raddr[10:5] ? tag_regs1_52 : _GEN_435; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_437 = 6'h35 == io_raddr[10:5] ? tag_regs1_53 : _GEN_436; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_438 = 6'h36 == io_raddr[10:5] ? tag_regs1_54 : _GEN_437; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_439 = 6'h37 == io_raddr[10:5] ? tag_regs1_55 : _GEN_438; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_440 = 6'h38 == io_raddr[10:5] ? tag_regs1_56 : _GEN_439; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_441 = 6'h39 == io_raddr[10:5] ? tag_regs1_57 : _GEN_440; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_442 = 6'h3a == io_raddr[10:5] ? tag_regs1_58 : _GEN_441; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_443 = 6'h3b == io_raddr[10:5] ? tag_regs1_59 : _GEN_442; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_444 = 6'h3c == io_raddr[10:5] ? tag_regs1_60 : _GEN_443; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_445 = 6'h3d == io_raddr[10:5] ? tag_regs1_61 : _GEN_444; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_446 = 6'h3e == io_raddr[10:5] ? tag_regs1_62 : _GEN_445; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_447 = 6'h3f == io_raddr[10:5] ? tag_regs1_63 : _GEN_446; // @[dcache_tag.scala 38:{44,44}]
  wire [21:0] _GEN_449 = 6'h1 == io_raddr[10:5] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_450 = 6'h2 == io_raddr[10:5] ? tag_regs0_2 : _GEN_449; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_451 = 6'h3 == io_raddr[10:5] ? tag_regs0_3 : _GEN_450; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_452 = 6'h4 == io_raddr[10:5] ? tag_regs0_4 : _GEN_451; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_453 = 6'h5 == io_raddr[10:5] ? tag_regs0_5 : _GEN_452; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_454 = 6'h6 == io_raddr[10:5] ? tag_regs0_6 : _GEN_453; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_455 = 6'h7 == io_raddr[10:5] ? tag_regs0_7 : _GEN_454; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_456 = 6'h8 == io_raddr[10:5] ? tag_regs0_8 : _GEN_455; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_457 = 6'h9 == io_raddr[10:5] ? tag_regs0_9 : _GEN_456; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_458 = 6'ha == io_raddr[10:5] ? tag_regs0_10 : _GEN_457; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_459 = 6'hb == io_raddr[10:5] ? tag_regs0_11 : _GEN_458; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_460 = 6'hc == io_raddr[10:5] ? tag_regs0_12 : _GEN_459; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_461 = 6'hd == io_raddr[10:5] ? tag_regs0_13 : _GEN_460; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_462 = 6'he == io_raddr[10:5] ? tag_regs0_14 : _GEN_461; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_463 = 6'hf == io_raddr[10:5] ? tag_regs0_15 : _GEN_462; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_464 = 6'h10 == io_raddr[10:5] ? tag_regs0_16 : _GEN_463; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_465 = 6'h11 == io_raddr[10:5] ? tag_regs0_17 : _GEN_464; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_466 = 6'h12 == io_raddr[10:5] ? tag_regs0_18 : _GEN_465; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_467 = 6'h13 == io_raddr[10:5] ? tag_regs0_19 : _GEN_466; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_468 = 6'h14 == io_raddr[10:5] ? tag_regs0_20 : _GEN_467; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_469 = 6'h15 == io_raddr[10:5] ? tag_regs0_21 : _GEN_468; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_470 = 6'h16 == io_raddr[10:5] ? tag_regs0_22 : _GEN_469; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_471 = 6'h17 == io_raddr[10:5] ? tag_regs0_23 : _GEN_470; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_472 = 6'h18 == io_raddr[10:5] ? tag_regs0_24 : _GEN_471; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_473 = 6'h19 == io_raddr[10:5] ? tag_regs0_25 : _GEN_472; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_474 = 6'h1a == io_raddr[10:5] ? tag_regs0_26 : _GEN_473; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_475 = 6'h1b == io_raddr[10:5] ? tag_regs0_27 : _GEN_474; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_476 = 6'h1c == io_raddr[10:5] ? tag_regs0_28 : _GEN_475; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_477 = 6'h1d == io_raddr[10:5] ? tag_regs0_29 : _GEN_476; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_478 = 6'h1e == io_raddr[10:5] ? tag_regs0_30 : _GEN_477; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_479 = 6'h1f == io_raddr[10:5] ? tag_regs0_31 : _GEN_478; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_480 = 6'h20 == io_raddr[10:5] ? tag_regs0_32 : _GEN_479; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_481 = 6'h21 == io_raddr[10:5] ? tag_regs0_33 : _GEN_480; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_482 = 6'h22 == io_raddr[10:5] ? tag_regs0_34 : _GEN_481; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_483 = 6'h23 == io_raddr[10:5] ? tag_regs0_35 : _GEN_482; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_484 = 6'h24 == io_raddr[10:5] ? tag_regs0_36 : _GEN_483; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_485 = 6'h25 == io_raddr[10:5] ? tag_regs0_37 : _GEN_484; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_486 = 6'h26 == io_raddr[10:5] ? tag_regs0_38 : _GEN_485; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_487 = 6'h27 == io_raddr[10:5] ? tag_regs0_39 : _GEN_486; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_488 = 6'h28 == io_raddr[10:5] ? tag_regs0_40 : _GEN_487; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_489 = 6'h29 == io_raddr[10:5] ? tag_regs0_41 : _GEN_488; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_490 = 6'h2a == io_raddr[10:5] ? tag_regs0_42 : _GEN_489; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_491 = 6'h2b == io_raddr[10:5] ? tag_regs0_43 : _GEN_490; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_492 = 6'h2c == io_raddr[10:5] ? tag_regs0_44 : _GEN_491; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_493 = 6'h2d == io_raddr[10:5] ? tag_regs0_45 : _GEN_492; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_494 = 6'h2e == io_raddr[10:5] ? tag_regs0_46 : _GEN_493; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_495 = 6'h2f == io_raddr[10:5] ? tag_regs0_47 : _GEN_494; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_496 = 6'h30 == io_raddr[10:5] ? tag_regs0_48 : _GEN_495; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_497 = 6'h31 == io_raddr[10:5] ? tag_regs0_49 : _GEN_496; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_498 = 6'h32 == io_raddr[10:5] ? tag_regs0_50 : _GEN_497; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_499 = 6'h33 == io_raddr[10:5] ? tag_regs0_51 : _GEN_498; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_500 = 6'h34 == io_raddr[10:5] ? tag_regs0_52 : _GEN_499; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_501 = 6'h35 == io_raddr[10:5] ? tag_regs0_53 : _GEN_500; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_502 = 6'h36 == io_raddr[10:5] ? tag_regs0_54 : _GEN_501; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_503 = 6'h37 == io_raddr[10:5] ? tag_regs0_55 : _GEN_502; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_504 = 6'h38 == io_raddr[10:5] ? tag_regs0_56 : _GEN_503; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_505 = 6'h39 == io_raddr[10:5] ? tag_regs0_57 : _GEN_504; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_506 = 6'h3a == io_raddr[10:5] ? tag_regs0_58 : _GEN_505; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_507 = 6'h3b == io_raddr[10:5] ? tag_regs0_59 : _GEN_506; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_508 = 6'h3c == io_raddr[10:5] ? tag_regs0_60 : _GEN_507; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_509 = 6'h3d == io_raddr[10:5] ? tag_regs0_61 : _GEN_508; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_510 = 6'h3e == io_raddr[10:5] ? tag_regs0_62 : _GEN_509; // @[dcache_tag.scala 38:{63,63}]
  wire [21:0] _GEN_511 = 6'h3f == io_raddr[10:5] ? tag_regs0_63 : _GEN_510; // @[dcache_tag.scala 38:{63,63}]
  wire  _io_hit_T_6 = ~io_raddr[4]; // @[dcache_tag.scala 39:91]
  wire  _io_hit_T_10 = _io_hit_T_6 & _GEN_511[20:0] == io_raddr[31:11]; // @[dcache_tag.scala 40:9]
  assign io_hit = io_raddr[4] & _GEN_447[20:0] == io_raddr[31:11] | _io_hit_T_10; // @[dcache_tag.scala 39:87]
  assign io_valid = io_raddr[4] ? _GEN_447[21] : _GEN_511[21]; // @[dcache_tag.scala 38:20]
  assign io_tag = io_waddr[4] ? _GEN_191[20:0] : _GEN_63[20:0]; // @[dcache_tag.scala 35:18]
  assign io_w_valid = io_waddr[4] ? _GEN_191[21] : _GEN_63[21]; // @[dcache_tag.scala 36:22]
  always @(posedge clock) begin
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_0 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h0 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_0 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_0 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_0 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_1 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_1 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_1 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_1 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_2 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_2 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_2 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_2 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_3 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_3 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_3 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_3 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_4 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h4 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_4 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_4 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_4 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_5 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h5 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_5 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_5 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_5 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_6 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h6 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_6 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_6 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_6 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_7 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h7 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_7 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_7 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_7 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_8 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h8 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_8 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_8 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_8 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_9 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h9 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_9 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_9 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_9 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_10 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'ha == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_10 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_10 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_10 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_11 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'hb == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_11 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_11 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_11 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_12 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'hc == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_12 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_12 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_12 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_13 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'hd == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_13 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_13 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_13 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_14 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'he == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_14 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_14 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_14 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_15 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'hf == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_15 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_15 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_15 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_16 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h10 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_16 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_16 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_16 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_17 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h11 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_17 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_17 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_17 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_18 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h12 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_18 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_18 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_18 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_19 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h13 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_19 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_19 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_19 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_20 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h14 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_20 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_20 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_20 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_21 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h15 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_21 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_21 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_21 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_22 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h16 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_22 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_22 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_22 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_23 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h17 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_23 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_23 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_23 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_24 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h18 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_24 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_24 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_24 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_25 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h19 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_25 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_25 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_25 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_26 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1a == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_26 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_26 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_26 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_27 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1b == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_27 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_27 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_27 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_28 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1c == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_28 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_28 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_28 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_29 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1d == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_29 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_29 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_29 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_30 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1e == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_30 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_30 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_30 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_31 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h1f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_31 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_31 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_31 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_32 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h20 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_32 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_32 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_32 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_33 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h21 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_33 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_33 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_33 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_34 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h22 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_34 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_34 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_34 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_35 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h23 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_35 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_35 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_35 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_36 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h24 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_36 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_36 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_36 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_37 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h25 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_37 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_37 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_37 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_38 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h26 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_38 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_38 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_38 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_39 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h27 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_39 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_39 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_39 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_40 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h28 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_40 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_40 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_40 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_41 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h29 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_41 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_41 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_41 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_42 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2a == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_42 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_42 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_42 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_43 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2b == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_43 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_43 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_43 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_44 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2c == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_44 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_44 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_44 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_45 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2d == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_45 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_45 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_45 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_46 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2e == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_46 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_46 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_46 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_47 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h2f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_47 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_47 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_47 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_48 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h30 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_48 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_48 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_48 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_49 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h31 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_49 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_49 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_49 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_50 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h32 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_50 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_50 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_50 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_51 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h33 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_51 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_51 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_51 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_52 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h34 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_52 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_52 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_52 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_53 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h35 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_53 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_53 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_53 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_54 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h36 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_54 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_54 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_54 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_55 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h37 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_55 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_55 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_55 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_56 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h38 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_56 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_56 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_56 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_57 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h39 == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_57 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_57 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_57 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_58 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3a == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_58 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_58 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_58 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_59 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3b == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_59 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_59 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_59 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_60 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3c == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_60 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_60 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_60 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_61 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3d == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_61 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_61 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_61 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_62 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3e == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_62 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_62 <= tag_regs0_63; // @[dcache_tag.scala 27:37]
      end else begin
        tag_regs0_62 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 23:28]
      tag_regs0_63 <= 22'h0; // @[dcache_tag.scala 23:28]
    end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 27:31]
      if (io_wen & ~io_waddr[4]) begin // @[dcache_tag.scala 27:37]
        tag_regs0_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[10:5])) begin // @[dcache_tag.scala 27:37]
        tag_regs0_63 <= _GEN_62;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_0 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h0 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_0 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_0 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_0 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_1 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_1 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_1 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_1 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_2 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_2 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_2 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_2 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_3 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_3 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_3 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_3 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_4 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h4 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_4 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_4 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_4 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_5 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h5 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_5 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_5 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_5 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_6 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h6 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_6 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_6 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_6 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_7 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h7 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_7 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_7 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_7 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_8 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h8 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_8 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_8 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_8 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_9 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h9 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_9 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_9 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_9 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_10 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'ha == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_10 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_10 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_10 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_11 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'hb == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_11 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_11 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_11 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_12 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'hc == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_12 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_12 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_12 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_13 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'hd == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_13 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_13 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_13 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_14 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'he == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_14 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_14 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_14 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_15 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'hf == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_15 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_15 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_15 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_16 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h10 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_16 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_16 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_16 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_17 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h11 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_17 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_17 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_17 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_18 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h12 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_18 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_18 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_18 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_19 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h13 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_19 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_19 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_19 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_20 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h14 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_20 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_20 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_20 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_21 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h15 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_21 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_21 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_21 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_22 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h16 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_22 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_22 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_22 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_23 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h17 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_23 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_23 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_23 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_24 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h18 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_24 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_24 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_24 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_25 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h19 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_25 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_25 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_25 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_26 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1a == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_26 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_26 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_26 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_27 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1b == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_27 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_27 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_27 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_28 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1c == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_28 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_28 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_28 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_29 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1d == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_29 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_29 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_29 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_30 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1e == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_30 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_30 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_30 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_31 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h1f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_31 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_31 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_31 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_32 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h20 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_32 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_32 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_32 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_33 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h21 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_33 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_33 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_33 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_34 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h22 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_34 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_34 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_34 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_35 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h23 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_35 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_35 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_35 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_36 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h24 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_36 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_36 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_36 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_37 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h25 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_37 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_37 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_37 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_38 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h26 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_38 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_38 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_38 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_39 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h27 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_39 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_39 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_39 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_40 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h28 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_40 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_40 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_40 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_41 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h29 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_41 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_41 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_41 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_42 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2a == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_42 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_42 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_42 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_43 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2b == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_43 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_43 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_43 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_44 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2c == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_44 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_44 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_44 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_45 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2d == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_45 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_45 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_45 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_46 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2e == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_46 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_46 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_46 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_47 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h2f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_47 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_47 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_47 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_48 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h30 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_48 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_48 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_48 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_49 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h31 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_49 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_49 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_49 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_50 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h32 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_50 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_50 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_50 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_51 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h33 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_51 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_51 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_51 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_52 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h34 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_52 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_52 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_52 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_53 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h35 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_53 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_53 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_53 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_54 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h36 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_54 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_54 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_54 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_55 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h37 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_55 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_55 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_55 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_56 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h38 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_56 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_56 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_56 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_57 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h39 == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_57 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_57 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_57 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_58 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3a == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_58 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_58 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_58 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_59 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3b == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_59 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_59 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_59 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_60 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3c == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_60 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_60 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_60 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_61 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3d == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_61 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_61 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_61 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_62 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3e == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_62 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_62 <= tag_regs1_63; // @[dcache_tag.scala 28:37]
      end else begin
        tag_regs1_62 <= _GEN_190;
      end
    end
    if (reset) begin // @[dcache_tag.scala 24:28]
      tag_regs1_63 <= 22'h0; // @[dcache_tag.scala 24:28]
    end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 28:31]
      if (io_wen & io_waddr[4]) begin // @[dcache_tag.scala 28:37]
        tag_regs1_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[10:5])) begin // @[dcache_tag.scala 28:37]
        tag_regs1_63 <= _GEN_190;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_regs0_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_regs0_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_regs0_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_regs0_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_regs0_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_regs0_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_regs0_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_regs0_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_regs0_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_regs0_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_regs0_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_regs0_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_regs0_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_regs0_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_regs0_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_regs0_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_regs0_16 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_regs0_17 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_regs0_18 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_regs0_19 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_regs0_20 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_regs0_21 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_regs0_22 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_regs0_23 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_regs0_24 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_regs0_25 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_regs0_26 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_regs0_27 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_regs0_28 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_regs0_29 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_regs0_30 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_regs0_31 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_regs0_32 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_regs0_33 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_regs0_34 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_regs0_35 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_regs0_36 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_regs0_37 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_regs0_38 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_regs0_39 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_regs0_40 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_regs0_41 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_regs0_42 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_regs0_43 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_regs0_44 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_regs0_45 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_regs0_46 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_regs0_47 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_regs0_48 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_regs0_49 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_regs0_50 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_regs0_51 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_regs0_52 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_regs0_53 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_regs0_54 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_regs0_55 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_regs0_56 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_regs0_57 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_regs0_58 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_regs0_59 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_regs0_60 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_regs0_61 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_regs0_62 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_regs0_63 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  tag_regs1_0 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  tag_regs1_1 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tag_regs1_2 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tag_regs1_3 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tag_regs1_4 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tag_regs1_5 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tag_regs1_6 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tag_regs1_7 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tag_regs1_8 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tag_regs1_9 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tag_regs1_10 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tag_regs1_11 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tag_regs1_12 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tag_regs1_13 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tag_regs1_14 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tag_regs1_15 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tag_regs1_16 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tag_regs1_17 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tag_regs1_18 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tag_regs1_19 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tag_regs1_20 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tag_regs1_21 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tag_regs1_22 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tag_regs1_23 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tag_regs1_24 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tag_regs1_25 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tag_regs1_26 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tag_regs1_27 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tag_regs1_28 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tag_regs1_29 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tag_regs1_30 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tag_regs1_31 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tag_regs1_32 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tag_regs1_33 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tag_regs1_34 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tag_regs1_35 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tag_regs1_36 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tag_regs1_37 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tag_regs1_38 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tag_regs1_39 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tag_regs1_40 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tag_regs1_41 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tag_regs1_42 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tag_regs1_43 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tag_regs1_44 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tag_regs1_45 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tag_regs1_46 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tag_regs1_47 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tag_regs1_48 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tag_regs1_49 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tag_regs1_50 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tag_regs1_51 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tag_regs1_52 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tag_regs1_53 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tag_regs1_54 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tag_regs1_55 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tag_regs1_56 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tag_regs1_57 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tag_regs1_58 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tag_regs1_59 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tag_regs1_60 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tag_regs1_61 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tag_regs1_62 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tag_regs1_63 = _RAND_127[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_dcache_data(
  input          clock,
  input  [7:0]   io_wen,
  input  [31:0]  io_addr,
  input  [63:0]  io_wdata,
  output [63:0]  io_rdata,
  output [5:0]   io_sram_addr,
  output         io_sram_wen,
  output [127:0] io_sram_wmask,
  output [127:0] io_sram_wdata,
  input  [127:0] io_sram_rdata
);
  wire  dcache_data_ram_0_clock; // @[dcache_data.scala 34:35]
  wire [7:0] dcache_data_ram_0_io_wea; // @[dcache_data.scala 34:35]
  wire [6:0] dcache_data_ram_0_io_addra; // @[dcache_data.scala 34:35]
  wire [63:0] dcache_data_ram_0_io_dina; // @[dcache_data.scala 34:35]
  wire [63:0] dcache_data_ram_0_io_douta; // @[dcache_data.scala 34:35]
  wire [5:0] dcache_data_ram_0_io_sram_port_addr; // @[dcache_data.scala 34:35]
  wire  dcache_data_ram_0_io_sram_port_wen; // @[dcache_data.scala 34:35]
  wire [127:0] dcache_data_ram_0_io_sram_port_wmask; // @[dcache_data.scala 34:35]
  wire [127:0] dcache_data_ram_0_io_sram_port_wdata; // @[dcache_data.scala 34:35]
  wire [127:0] dcache_data_ram_0_io_sram_port_rdata; // @[dcache_data.scala 34:35]
  ysyx_22040886_ysyx_sram_with_mask dcache_data_ram_0 ( // @[dcache_data.scala 34:35]
    .clock(dcache_data_ram_0_clock),
    .io_wea(dcache_data_ram_0_io_wea),
    .io_addra(dcache_data_ram_0_io_addra),
    .io_dina(dcache_data_ram_0_io_dina),
    .io_douta(dcache_data_ram_0_io_douta),
    .io_sram_port_addr(dcache_data_ram_0_io_sram_port_addr),
    .io_sram_port_wen(dcache_data_ram_0_io_sram_port_wen),
    .io_sram_port_wmask(dcache_data_ram_0_io_sram_port_wmask),
    .io_sram_port_wdata(dcache_data_ram_0_io_sram_port_wdata),
    .io_sram_port_rdata(dcache_data_ram_0_io_sram_port_rdata)
  );
  assign io_rdata = dcache_data_ram_0_io_douta; // @[dcache_data.scala 41:16]
  assign io_sram_addr = dcache_data_ram_0_io_sram_port_addr; // @[dcache_data.scala 39:13]
  assign io_sram_wen = dcache_data_ram_0_io_sram_port_wen; // @[dcache_data.scala 39:13]
  assign io_sram_wmask = dcache_data_ram_0_io_sram_port_wmask; // @[dcache_data.scala 39:13]
  assign io_sram_wdata = dcache_data_ram_0_io_sram_port_wdata; // @[dcache_data.scala 39:13]
  assign dcache_data_ram_0_clock = clock;
  assign dcache_data_ram_0_io_wea = io_wen; // @[dcache_data.scala 36:31]
  assign dcache_data_ram_0_io_addra = io_addr[10:4]; // @[dcache_data.scala 37:42]
  assign dcache_data_ram_0_io_dina = io_wdata; // @[dcache_data.scala 38:31]
  assign dcache_data_ram_0_io_sram_port_rdata = io_sram_rdata; // @[dcache_data.scala 39:13]
endmodule
module ysyx_22040886_data_cache(
  input          clock,
  input          reset,
  output [31:0]  io_port_araddr,
  output [7:0]   io_port_arlen,
  output [2:0]   io_port_arsize,
  output [1:0]   io_port_arburst,
  output         io_port_arvalid,
  input          io_port_arready,
  input  [63:0]  io_port_rdata,
  input          io_port_rlast,
  input          io_port_rvalid,
  output [31:0]  io_port_awaddr,
  output [7:0]   io_port_awlen,
  output [2:0]   io_port_awsize,
  output [1:0]   io_port_awburst,
  output         io_port_awvalid,
  input          io_port_awready,
  output [63:0]  io_port_wdata,
  output [7:0]   io_port_wstrb,
  output         io_port_wlast,
  output         io_port_wvalid,
  input          io_port_wready,
  input          io_port_bvalid,
  output         io_stage2_stall,
  output [31:0]  io_v_addr_for_tlb,
  input  [31:0]  io_p_addr_for_tlb,
  input  [7:0]   io_data_wstrb,
  input          io_sram_req,
  input          io_sram_wr,
  input  [2:0]   io_sram_size,
  input  [31:0]  io_sram_addr,
  input  [63:0]  io_sram_wdata,
  output [63:0]  io_sram_rdata,
  input          io_sram_cache,
  input          io_fence_i_control,
  output [5:0]   io_sram_0_addr,
  output         io_sram_0_wen,
  output [127:0] io_sram_0_wmask,
  output [127:0] io_sram_0_wdata,
  input  [127:0] io_sram_0_rdata,
  output [5:0]   io_sram_1_addr,
  output         io_sram_1_wen,
  output [127:0] io_sram_1_wmask,
  output [127:0] io_sram_1_wdata,
  input  [127:0] io_sram_1_rdata,
  output [5:0]   io_sram_2_addr,
  output         io_sram_2_wen,
  output [127:0] io_sram_2_wmask,
  output [127:0] io_sram_2_wdata,
  input  [127:0] io_sram_2_rdata,
  output [5:0]   io_sram_3_addr,
  output         io_sram_3_wen,
  output [127:0] io_sram_3_wmask,
  output [127:0] io_sram_3_wdata,
  input  [127:0] io_sram_3_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [63:0] _RAND_406;
  reg [31:0] _RAND_407;
`endif // RANDOMIZE_REG_INIT
  wire  dcache_tag_clock; // @[data_cache.scala 62:30]
  wire  dcache_tag_reset; // @[data_cache.scala 62:30]
  wire  dcache_tag_io_wen; // @[data_cache.scala 62:30]
  wire [21:0] dcache_tag_io_wdata; // @[data_cache.scala 62:30]
  wire [31:0] dcache_tag_io_raddr; // @[data_cache.scala 62:30]
  wire [31:0] dcache_tag_io_waddr; // @[data_cache.scala 62:30]
  wire  dcache_tag_io_hit; // @[data_cache.scala 62:30]
  wire  dcache_tag_io_valid; // @[data_cache.scala 62:30]
  wire [20:0] dcache_tag_io_tag; // @[data_cache.scala 62:30]
  wire  dcache_tag_io_w_valid; // @[data_cache.scala 62:30]
  wire  dcache_tag_1_clock; // @[data_cache.scala 63:30]
  wire  dcache_tag_1_reset; // @[data_cache.scala 63:30]
  wire  dcache_tag_1_io_wen; // @[data_cache.scala 63:30]
  wire [21:0] dcache_tag_1_io_wdata; // @[data_cache.scala 63:30]
  wire [31:0] dcache_tag_1_io_raddr; // @[data_cache.scala 63:30]
  wire [31:0] dcache_tag_1_io_waddr; // @[data_cache.scala 63:30]
  wire  dcache_tag_1_io_hit; // @[data_cache.scala 63:30]
  wire  dcache_tag_1_io_valid; // @[data_cache.scala 63:30]
  wire [20:0] dcache_tag_1_io_tag; // @[data_cache.scala 63:30]
  wire  dcache_tag_1_io_w_valid; // @[data_cache.scala 63:30]
  wire  dcache_data_clock; // @[data_cache.scala 95:62]
  wire [7:0] dcache_data_io_wen; // @[data_cache.scala 95:62]
  wire [31:0] dcache_data_io_addr; // @[data_cache.scala 95:62]
  wire [63:0] dcache_data_io_wdata; // @[data_cache.scala 95:62]
  wire [63:0] dcache_data_io_rdata; // @[data_cache.scala 95:62]
  wire [5:0] dcache_data_io_sram_addr; // @[data_cache.scala 95:62]
  wire  dcache_data_io_sram_wen; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_io_sram_wmask; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_io_sram_wdata; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_io_sram_rdata; // @[data_cache.scala 95:62]
  wire  dcache_data_1_clock; // @[data_cache.scala 95:62]
  wire [7:0] dcache_data_1_io_wen; // @[data_cache.scala 95:62]
  wire [31:0] dcache_data_1_io_addr; // @[data_cache.scala 95:62]
  wire [63:0] dcache_data_1_io_wdata; // @[data_cache.scala 95:62]
  wire [63:0] dcache_data_1_io_rdata; // @[data_cache.scala 95:62]
  wire [5:0] dcache_data_1_io_sram_addr; // @[data_cache.scala 95:62]
  wire  dcache_data_1_io_sram_wen; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_1_io_sram_wmask; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_1_io_sram_wdata; // @[data_cache.scala 95:62]
  wire [127:0] dcache_data_1_io_sram_rdata; // @[data_cache.scala 95:62]
  wire  dcache_data_2_clock; // @[data_cache.scala 96:62]
  wire [7:0] dcache_data_2_io_wen; // @[data_cache.scala 96:62]
  wire [31:0] dcache_data_2_io_addr; // @[data_cache.scala 96:62]
  wire [63:0] dcache_data_2_io_wdata; // @[data_cache.scala 96:62]
  wire [63:0] dcache_data_2_io_rdata; // @[data_cache.scala 96:62]
  wire [5:0] dcache_data_2_io_sram_addr; // @[data_cache.scala 96:62]
  wire  dcache_data_2_io_sram_wen; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_2_io_sram_wmask; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_2_io_sram_wdata; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_2_io_sram_rdata; // @[data_cache.scala 96:62]
  wire  dcache_data_3_clock; // @[data_cache.scala 96:62]
  wire [7:0] dcache_data_3_io_wen; // @[data_cache.scala 96:62]
  wire [31:0] dcache_data_3_io_addr; // @[data_cache.scala 96:62]
  wire [63:0] dcache_data_3_io_wdata; // @[data_cache.scala 96:62]
  wire [63:0] dcache_data_3_io_rdata; // @[data_cache.scala 96:62]
  wire [5:0] dcache_data_3_io_sram_addr; // @[data_cache.scala 96:62]
  wire  dcache_data_3_io_sram_wen; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_3_io_sram_wmask; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_3_io_sram_wdata; // @[data_cache.scala 96:62]
  wire [127:0] dcache_data_3_io_sram_rdata; // @[data_cache.scala 96:62]
  reg [4:0] work_state; // @[data_cache.scala 55:29]
  reg [2:0] write_counter; // @[data_cache.scala 57:33]
  reg [2:0] read_counter; // @[data_cache.scala 58:32]
  reg [63:0] wait_data; // @[data_cache.scala 59:29]
  reg  lru_0; // @[data_cache.scala 65:22]
  reg  lru_1; // @[data_cache.scala 65:22]
  reg  lru_2; // @[data_cache.scala 65:22]
  reg  lru_3; // @[data_cache.scala 65:22]
  reg  lru_4; // @[data_cache.scala 65:22]
  reg  lru_5; // @[data_cache.scala 65:22]
  reg  lru_6; // @[data_cache.scala 65:22]
  reg  lru_7; // @[data_cache.scala 65:22]
  reg  lru_8; // @[data_cache.scala 65:22]
  reg  lru_9; // @[data_cache.scala 65:22]
  reg  lru_10; // @[data_cache.scala 65:22]
  reg  lru_11; // @[data_cache.scala 65:22]
  reg  lru_12; // @[data_cache.scala 65:22]
  reg  lru_13; // @[data_cache.scala 65:22]
  reg  lru_14; // @[data_cache.scala 65:22]
  reg  lru_15; // @[data_cache.scala 65:22]
  reg  lru_16; // @[data_cache.scala 65:22]
  reg  lru_17; // @[data_cache.scala 65:22]
  reg  lru_18; // @[data_cache.scala 65:22]
  reg  lru_19; // @[data_cache.scala 65:22]
  reg  lru_20; // @[data_cache.scala 65:22]
  reg  lru_21; // @[data_cache.scala 65:22]
  reg  lru_22; // @[data_cache.scala 65:22]
  reg  lru_23; // @[data_cache.scala 65:22]
  reg  lru_24; // @[data_cache.scala 65:22]
  reg  lru_25; // @[data_cache.scala 65:22]
  reg  lru_26; // @[data_cache.scala 65:22]
  reg  lru_27; // @[data_cache.scala 65:22]
  reg  lru_28; // @[data_cache.scala 65:22]
  reg  lru_29; // @[data_cache.scala 65:22]
  reg  lru_30; // @[data_cache.scala 65:22]
  reg  lru_31; // @[data_cache.scala 65:22]
  reg  lru_32; // @[data_cache.scala 65:22]
  reg  lru_33; // @[data_cache.scala 65:22]
  reg  lru_34; // @[data_cache.scala 65:22]
  reg  lru_35; // @[data_cache.scala 65:22]
  reg  lru_36; // @[data_cache.scala 65:22]
  reg  lru_37; // @[data_cache.scala 65:22]
  reg  lru_38; // @[data_cache.scala 65:22]
  reg  lru_39; // @[data_cache.scala 65:22]
  reg  lru_40; // @[data_cache.scala 65:22]
  reg  lru_41; // @[data_cache.scala 65:22]
  reg  lru_42; // @[data_cache.scala 65:22]
  reg  lru_43; // @[data_cache.scala 65:22]
  reg  lru_44; // @[data_cache.scala 65:22]
  reg  lru_45; // @[data_cache.scala 65:22]
  reg  lru_46; // @[data_cache.scala 65:22]
  reg  lru_47; // @[data_cache.scala 65:22]
  reg  lru_48; // @[data_cache.scala 65:22]
  reg  lru_49; // @[data_cache.scala 65:22]
  reg  lru_50; // @[data_cache.scala 65:22]
  reg  lru_51; // @[data_cache.scala 65:22]
  reg  lru_52; // @[data_cache.scala 65:22]
  reg  lru_53; // @[data_cache.scala 65:22]
  reg  lru_54; // @[data_cache.scala 65:22]
  reg  lru_55; // @[data_cache.scala 65:22]
  reg  lru_56; // @[data_cache.scala 65:22]
  reg  lru_57; // @[data_cache.scala 65:22]
  reg  lru_58; // @[data_cache.scala 65:22]
  reg  lru_59; // @[data_cache.scala 65:22]
  reg  lru_60; // @[data_cache.scala 65:22]
  reg  lru_61; // @[data_cache.scala 65:22]
  reg  lru_62; // @[data_cache.scala 65:22]
  reg  lru_63; // @[data_cache.scala 65:22]
  reg  lru_64; // @[data_cache.scala 65:22]
  reg  lru_65; // @[data_cache.scala 65:22]
  reg  lru_66; // @[data_cache.scala 65:22]
  reg  lru_67; // @[data_cache.scala 65:22]
  reg  lru_68; // @[data_cache.scala 65:22]
  reg  lru_69; // @[data_cache.scala 65:22]
  reg  lru_70; // @[data_cache.scala 65:22]
  reg  lru_71; // @[data_cache.scala 65:22]
  reg  lru_72; // @[data_cache.scala 65:22]
  reg  lru_73; // @[data_cache.scala 65:22]
  reg  lru_74; // @[data_cache.scala 65:22]
  reg  lru_75; // @[data_cache.scala 65:22]
  reg  lru_76; // @[data_cache.scala 65:22]
  reg  lru_77; // @[data_cache.scala 65:22]
  reg  lru_78; // @[data_cache.scala 65:22]
  reg  lru_79; // @[data_cache.scala 65:22]
  reg  lru_80; // @[data_cache.scala 65:22]
  reg  lru_81; // @[data_cache.scala 65:22]
  reg  lru_82; // @[data_cache.scala 65:22]
  reg  lru_83; // @[data_cache.scala 65:22]
  reg  lru_84; // @[data_cache.scala 65:22]
  reg  lru_85; // @[data_cache.scala 65:22]
  reg  lru_86; // @[data_cache.scala 65:22]
  reg  lru_87; // @[data_cache.scala 65:22]
  reg  lru_88; // @[data_cache.scala 65:22]
  reg  lru_89; // @[data_cache.scala 65:22]
  reg  lru_90; // @[data_cache.scala 65:22]
  reg  lru_91; // @[data_cache.scala 65:22]
  reg  lru_92; // @[data_cache.scala 65:22]
  reg  lru_93; // @[data_cache.scala 65:22]
  reg  lru_94; // @[data_cache.scala 65:22]
  reg  lru_95; // @[data_cache.scala 65:22]
  reg  lru_96; // @[data_cache.scala 65:22]
  reg  lru_97; // @[data_cache.scala 65:22]
  reg  lru_98; // @[data_cache.scala 65:22]
  reg  lru_99; // @[data_cache.scala 65:22]
  reg  lru_100; // @[data_cache.scala 65:22]
  reg  lru_101; // @[data_cache.scala 65:22]
  reg  lru_102; // @[data_cache.scala 65:22]
  reg  lru_103; // @[data_cache.scala 65:22]
  reg  lru_104; // @[data_cache.scala 65:22]
  reg  lru_105; // @[data_cache.scala 65:22]
  reg  lru_106; // @[data_cache.scala 65:22]
  reg  lru_107; // @[data_cache.scala 65:22]
  reg  lru_108; // @[data_cache.scala 65:22]
  reg  lru_109; // @[data_cache.scala 65:22]
  reg  lru_110; // @[data_cache.scala 65:22]
  reg  lru_111; // @[data_cache.scala 65:22]
  reg  lru_112; // @[data_cache.scala 65:22]
  reg  lru_113; // @[data_cache.scala 65:22]
  reg  lru_114; // @[data_cache.scala 65:22]
  reg  lru_115; // @[data_cache.scala 65:22]
  reg  lru_116; // @[data_cache.scala 65:22]
  reg  lru_117; // @[data_cache.scala 65:22]
  reg  lru_118; // @[data_cache.scala 65:22]
  reg  lru_119; // @[data_cache.scala 65:22]
  reg  lru_120; // @[data_cache.scala 65:22]
  reg  lru_121; // @[data_cache.scala 65:22]
  reg  lru_122; // @[data_cache.scala 65:22]
  reg  lru_123; // @[data_cache.scala 65:22]
  reg  lru_124; // @[data_cache.scala 65:22]
  reg  lru_125; // @[data_cache.scala 65:22]
  reg  lru_126; // @[data_cache.scala 65:22]
  reg  lru_127; // @[data_cache.scala 65:22]
  reg  way0_dirty_0; // @[data_cache.scala 66:29]
  reg  way0_dirty_1; // @[data_cache.scala 66:29]
  reg  way0_dirty_2; // @[data_cache.scala 66:29]
  reg  way0_dirty_3; // @[data_cache.scala 66:29]
  reg  way0_dirty_4; // @[data_cache.scala 66:29]
  reg  way0_dirty_5; // @[data_cache.scala 66:29]
  reg  way0_dirty_6; // @[data_cache.scala 66:29]
  reg  way0_dirty_7; // @[data_cache.scala 66:29]
  reg  way0_dirty_8; // @[data_cache.scala 66:29]
  reg  way0_dirty_9; // @[data_cache.scala 66:29]
  reg  way0_dirty_10; // @[data_cache.scala 66:29]
  reg  way0_dirty_11; // @[data_cache.scala 66:29]
  reg  way0_dirty_12; // @[data_cache.scala 66:29]
  reg  way0_dirty_13; // @[data_cache.scala 66:29]
  reg  way0_dirty_14; // @[data_cache.scala 66:29]
  reg  way0_dirty_15; // @[data_cache.scala 66:29]
  reg  way0_dirty_16; // @[data_cache.scala 66:29]
  reg  way0_dirty_17; // @[data_cache.scala 66:29]
  reg  way0_dirty_18; // @[data_cache.scala 66:29]
  reg  way0_dirty_19; // @[data_cache.scala 66:29]
  reg  way0_dirty_20; // @[data_cache.scala 66:29]
  reg  way0_dirty_21; // @[data_cache.scala 66:29]
  reg  way0_dirty_22; // @[data_cache.scala 66:29]
  reg  way0_dirty_23; // @[data_cache.scala 66:29]
  reg  way0_dirty_24; // @[data_cache.scala 66:29]
  reg  way0_dirty_25; // @[data_cache.scala 66:29]
  reg  way0_dirty_26; // @[data_cache.scala 66:29]
  reg  way0_dirty_27; // @[data_cache.scala 66:29]
  reg  way0_dirty_28; // @[data_cache.scala 66:29]
  reg  way0_dirty_29; // @[data_cache.scala 66:29]
  reg  way0_dirty_30; // @[data_cache.scala 66:29]
  reg  way0_dirty_31; // @[data_cache.scala 66:29]
  reg  way0_dirty_32; // @[data_cache.scala 66:29]
  reg  way0_dirty_33; // @[data_cache.scala 66:29]
  reg  way0_dirty_34; // @[data_cache.scala 66:29]
  reg  way0_dirty_35; // @[data_cache.scala 66:29]
  reg  way0_dirty_36; // @[data_cache.scala 66:29]
  reg  way0_dirty_37; // @[data_cache.scala 66:29]
  reg  way0_dirty_38; // @[data_cache.scala 66:29]
  reg  way0_dirty_39; // @[data_cache.scala 66:29]
  reg  way0_dirty_40; // @[data_cache.scala 66:29]
  reg  way0_dirty_41; // @[data_cache.scala 66:29]
  reg  way0_dirty_42; // @[data_cache.scala 66:29]
  reg  way0_dirty_43; // @[data_cache.scala 66:29]
  reg  way0_dirty_44; // @[data_cache.scala 66:29]
  reg  way0_dirty_45; // @[data_cache.scala 66:29]
  reg  way0_dirty_46; // @[data_cache.scala 66:29]
  reg  way0_dirty_47; // @[data_cache.scala 66:29]
  reg  way0_dirty_48; // @[data_cache.scala 66:29]
  reg  way0_dirty_49; // @[data_cache.scala 66:29]
  reg  way0_dirty_50; // @[data_cache.scala 66:29]
  reg  way0_dirty_51; // @[data_cache.scala 66:29]
  reg  way0_dirty_52; // @[data_cache.scala 66:29]
  reg  way0_dirty_53; // @[data_cache.scala 66:29]
  reg  way0_dirty_54; // @[data_cache.scala 66:29]
  reg  way0_dirty_55; // @[data_cache.scala 66:29]
  reg  way0_dirty_56; // @[data_cache.scala 66:29]
  reg  way0_dirty_57; // @[data_cache.scala 66:29]
  reg  way0_dirty_58; // @[data_cache.scala 66:29]
  reg  way0_dirty_59; // @[data_cache.scala 66:29]
  reg  way0_dirty_60; // @[data_cache.scala 66:29]
  reg  way0_dirty_61; // @[data_cache.scala 66:29]
  reg  way0_dirty_62; // @[data_cache.scala 66:29]
  reg  way0_dirty_63; // @[data_cache.scala 66:29]
  reg  way0_dirty_64; // @[data_cache.scala 66:29]
  reg  way0_dirty_65; // @[data_cache.scala 66:29]
  reg  way0_dirty_66; // @[data_cache.scala 66:29]
  reg  way0_dirty_67; // @[data_cache.scala 66:29]
  reg  way0_dirty_68; // @[data_cache.scala 66:29]
  reg  way0_dirty_69; // @[data_cache.scala 66:29]
  reg  way0_dirty_70; // @[data_cache.scala 66:29]
  reg  way0_dirty_71; // @[data_cache.scala 66:29]
  reg  way0_dirty_72; // @[data_cache.scala 66:29]
  reg  way0_dirty_73; // @[data_cache.scala 66:29]
  reg  way0_dirty_74; // @[data_cache.scala 66:29]
  reg  way0_dirty_75; // @[data_cache.scala 66:29]
  reg  way0_dirty_76; // @[data_cache.scala 66:29]
  reg  way0_dirty_77; // @[data_cache.scala 66:29]
  reg  way0_dirty_78; // @[data_cache.scala 66:29]
  reg  way0_dirty_79; // @[data_cache.scala 66:29]
  reg  way0_dirty_80; // @[data_cache.scala 66:29]
  reg  way0_dirty_81; // @[data_cache.scala 66:29]
  reg  way0_dirty_82; // @[data_cache.scala 66:29]
  reg  way0_dirty_83; // @[data_cache.scala 66:29]
  reg  way0_dirty_84; // @[data_cache.scala 66:29]
  reg  way0_dirty_85; // @[data_cache.scala 66:29]
  reg  way0_dirty_86; // @[data_cache.scala 66:29]
  reg  way0_dirty_87; // @[data_cache.scala 66:29]
  reg  way0_dirty_88; // @[data_cache.scala 66:29]
  reg  way0_dirty_89; // @[data_cache.scala 66:29]
  reg  way0_dirty_90; // @[data_cache.scala 66:29]
  reg  way0_dirty_91; // @[data_cache.scala 66:29]
  reg  way0_dirty_92; // @[data_cache.scala 66:29]
  reg  way0_dirty_93; // @[data_cache.scala 66:29]
  reg  way0_dirty_94; // @[data_cache.scala 66:29]
  reg  way0_dirty_95; // @[data_cache.scala 66:29]
  reg  way0_dirty_96; // @[data_cache.scala 66:29]
  reg  way0_dirty_97; // @[data_cache.scala 66:29]
  reg  way0_dirty_98; // @[data_cache.scala 66:29]
  reg  way0_dirty_99; // @[data_cache.scala 66:29]
  reg  way0_dirty_100; // @[data_cache.scala 66:29]
  reg  way0_dirty_101; // @[data_cache.scala 66:29]
  reg  way0_dirty_102; // @[data_cache.scala 66:29]
  reg  way0_dirty_103; // @[data_cache.scala 66:29]
  reg  way0_dirty_104; // @[data_cache.scala 66:29]
  reg  way0_dirty_105; // @[data_cache.scala 66:29]
  reg  way0_dirty_106; // @[data_cache.scala 66:29]
  reg  way0_dirty_107; // @[data_cache.scala 66:29]
  reg  way0_dirty_108; // @[data_cache.scala 66:29]
  reg  way0_dirty_109; // @[data_cache.scala 66:29]
  reg  way0_dirty_110; // @[data_cache.scala 66:29]
  reg  way0_dirty_111; // @[data_cache.scala 66:29]
  reg  way0_dirty_112; // @[data_cache.scala 66:29]
  reg  way0_dirty_113; // @[data_cache.scala 66:29]
  reg  way0_dirty_114; // @[data_cache.scala 66:29]
  reg  way0_dirty_115; // @[data_cache.scala 66:29]
  reg  way0_dirty_116; // @[data_cache.scala 66:29]
  reg  way0_dirty_117; // @[data_cache.scala 66:29]
  reg  way0_dirty_118; // @[data_cache.scala 66:29]
  reg  way0_dirty_119; // @[data_cache.scala 66:29]
  reg  way0_dirty_120; // @[data_cache.scala 66:29]
  reg  way0_dirty_121; // @[data_cache.scala 66:29]
  reg  way0_dirty_122; // @[data_cache.scala 66:29]
  reg  way0_dirty_123; // @[data_cache.scala 66:29]
  reg  way0_dirty_124; // @[data_cache.scala 66:29]
  reg  way0_dirty_125; // @[data_cache.scala 66:29]
  reg  way0_dirty_126; // @[data_cache.scala 66:29]
  reg  way0_dirty_127; // @[data_cache.scala 66:29]
  reg  way1_dirty_0; // @[data_cache.scala 67:29]
  reg  way1_dirty_1; // @[data_cache.scala 67:29]
  reg  way1_dirty_2; // @[data_cache.scala 67:29]
  reg  way1_dirty_3; // @[data_cache.scala 67:29]
  reg  way1_dirty_4; // @[data_cache.scala 67:29]
  reg  way1_dirty_5; // @[data_cache.scala 67:29]
  reg  way1_dirty_6; // @[data_cache.scala 67:29]
  reg  way1_dirty_7; // @[data_cache.scala 67:29]
  reg  way1_dirty_8; // @[data_cache.scala 67:29]
  reg  way1_dirty_9; // @[data_cache.scala 67:29]
  reg  way1_dirty_10; // @[data_cache.scala 67:29]
  reg  way1_dirty_11; // @[data_cache.scala 67:29]
  reg  way1_dirty_12; // @[data_cache.scala 67:29]
  reg  way1_dirty_13; // @[data_cache.scala 67:29]
  reg  way1_dirty_14; // @[data_cache.scala 67:29]
  reg  way1_dirty_15; // @[data_cache.scala 67:29]
  reg  way1_dirty_16; // @[data_cache.scala 67:29]
  reg  way1_dirty_17; // @[data_cache.scala 67:29]
  reg  way1_dirty_18; // @[data_cache.scala 67:29]
  reg  way1_dirty_19; // @[data_cache.scala 67:29]
  reg  way1_dirty_20; // @[data_cache.scala 67:29]
  reg  way1_dirty_21; // @[data_cache.scala 67:29]
  reg  way1_dirty_22; // @[data_cache.scala 67:29]
  reg  way1_dirty_23; // @[data_cache.scala 67:29]
  reg  way1_dirty_24; // @[data_cache.scala 67:29]
  reg  way1_dirty_25; // @[data_cache.scala 67:29]
  reg  way1_dirty_26; // @[data_cache.scala 67:29]
  reg  way1_dirty_27; // @[data_cache.scala 67:29]
  reg  way1_dirty_28; // @[data_cache.scala 67:29]
  reg  way1_dirty_29; // @[data_cache.scala 67:29]
  reg  way1_dirty_30; // @[data_cache.scala 67:29]
  reg  way1_dirty_31; // @[data_cache.scala 67:29]
  reg  way1_dirty_32; // @[data_cache.scala 67:29]
  reg  way1_dirty_33; // @[data_cache.scala 67:29]
  reg  way1_dirty_34; // @[data_cache.scala 67:29]
  reg  way1_dirty_35; // @[data_cache.scala 67:29]
  reg  way1_dirty_36; // @[data_cache.scala 67:29]
  reg  way1_dirty_37; // @[data_cache.scala 67:29]
  reg  way1_dirty_38; // @[data_cache.scala 67:29]
  reg  way1_dirty_39; // @[data_cache.scala 67:29]
  reg  way1_dirty_40; // @[data_cache.scala 67:29]
  reg  way1_dirty_41; // @[data_cache.scala 67:29]
  reg  way1_dirty_42; // @[data_cache.scala 67:29]
  reg  way1_dirty_43; // @[data_cache.scala 67:29]
  reg  way1_dirty_44; // @[data_cache.scala 67:29]
  reg  way1_dirty_45; // @[data_cache.scala 67:29]
  reg  way1_dirty_46; // @[data_cache.scala 67:29]
  reg  way1_dirty_47; // @[data_cache.scala 67:29]
  reg  way1_dirty_48; // @[data_cache.scala 67:29]
  reg  way1_dirty_49; // @[data_cache.scala 67:29]
  reg  way1_dirty_50; // @[data_cache.scala 67:29]
  reg  way1_dirty_51; // @[data_cache.scala 67:29]
  reg  way1_dirty_52; // @[data_cache.scala 67:29]
  reg  way1_dirty_53; // @[data_cache.scala 67:29]
  reg  way1_dirty_54; // @[data_cache.scala 67:29]
  reg  way1_dirty_55; // @[data_cache.scala 67:29]
  reg  way1_dirty_56; // @[data_cache.scala 67:29]
  reg  way1_dirty_57; // @[data_cache.scala 67:29]
  reg  way1_dirty_58; // @[data_cache.scala 67:29]
  reg  way1_dirty_59; // @[data_cache.scala 67:29]
  reg  way1_dirty_60; // @[data_cache.scala 67:29]
  reg  way1_dirty_61; // @[data_cache.scala 67:29]
  reg  way1_dirty_62; // @[data_cache.scala 67:29]
  reg  way1_dirty_63; // @[data_cache.scala 67:29]
  reg  way1_dirty_64; // @[data_cache.scala 67:29]
  reg  way1_dirty_65; // @[data_cache.scala 67:29]
  reg  way1_dirty_66; // @[data_cache.scala 67:29]
  reg  way1_dirty_67; // @[data_cache.scala 67:29]
  reg  way1_dirty_68; // @[data_cache.scala 67:29]
  reg  way1_dirty_69; // @[data_cache.scala 67:29]
  reg  way1_dirty_70; // @[data_cache.scala 67:29]
  reg  way1_dirty_71; // @[data_cache.scala 67:29]
  reg  way1_dirty_72; // @[data_cache.scala 67:29]
  reg  way1_dirty_73; // @[data_cache.scala 67:29]
  reg  way1_dirty_74; // @[data_cache.scala 67:29]
  reg  way1_dirty_75; // @[data_cache.scala 67:29]
  reg  way1_dirty_76; // @[data_cache.scala 67:29]
  reg  way1_dirty_77; // @[data_cache.scala 67:29]
  reg  way1_dirty_78; // @[data_cache.scala 67:29]
  reg  way1_dirty_79; // @[data_cache.scala 67:29]
  reg  way1_dirty_80; // @[data_cache.scala 67:29]
  reg  way1_dirty_81; // @[data_cache.scala 67:29]
  reg  way1_dirty_82; // @[data_cache.scala 67:29]
  reg  way1_dirty_83; // @[data_cache.scala 67:29]
  reg  way1_dirty_84; // @[data_cache.scala 67:29]
  reg  way1_dirty_85; // @[data_cache.scala 67:29]
  reg  way1_dirty_86; // @[data_cache.scala 67:29]
  reg  way1_dirty_87; // @[data_cache.scala 67:29]
  reg  way1_dirty_88; // @[data_cache.scala 67:29]
  reg  way1_dirty_89; // @[data_cache.scala 67:29]
  reg  way1_dirty_90; // @[data_cache.scala 67:29]
  reg  way1_dirty_91; // @[data_cache.scala 67:29]
  reg  way1_dirty_92; // @[data_cache.scala 67:29]
  reg  way1_dirty_93; // @[data_cache.scala 67:29]
  reg  way1_dirty_94; // @[data_cache.scala 67:29]
  reg  way1_dirty_95; // @[data_cache.scala 67:29]
  reg  way1_dirty_96; // @[data_cache.scala 67:29]
  reg  way1_dirty_97; // @[data_cache.scala 67:29]
  reg  way1_dirty_98; // @[data_cache.scala 67:29]
  reg  way1_dirty_99; // @[data_cache.scala 67:29]
  reg  way1_dirty_100; // @[data_cache.scala 67:29]
  reg  way1_dirty_101; // @[data_cache.scala 67:29]
  reg  way1_dirty_102; // @[data_cache.scala 67:29]
  reg  way1_dirty_103; // @[data_cache.scala 67:29]
  reg  way1_dirty_104; // @[data_cache.scala 67:29]
  reg  way1_dirty_105; // @[data_cache.scala 67:29]
  reg  way1_dirty_106; // @[data_cache.scala 67:29]
  reg  way1_dirty_107; // @[data_cache.scala 67:29]
  reg  way1_dirty_108; // @[data_cache.scala 67:29]
  reg  way1_dirty_109; // @[data_cache.scala 67:29]
  reg  way1_dirty_110; // @[data_cache.scala 67:29]
  reg  way1_dirty_111; // @[data_cache.scala 67:29]
  reg  way1_dirty_112; // @[data_cache.scala 67:29]
  reg  way1_dirty_113; // @[data_cache.scala 67:29]
  reg  way1_dirty_114; // @[data_cache.scala 67:29]
  reg  way1_dirty_115; // @[data_cache.scala 67:29]
  reg  way1_dirty_116; // @[data_cache.scala 67:29]
  reg  way1_dirty_117; // @[data_cache.scala 67:29]
  reg  way1_dirty_118; // @[data_cache.scala 67:29]
  reg  way1_dirty_119; // @[data_cache.scala 67:29]
  reg  way1_dirty_120; // @[data_cache.scala 67:29]
  reg  way1_dirty_121; // @[data_cache.scala 67:29]
  reg  way1_dirty_122; // @[data_cache.scala 67:29]
  reg  way1_dirty_123; // @[data_cache.scala 67:29]
  reg  way1_dirty_124; // @[data_cache.scala 67:29]
  reg  way1_dirty_125; // @[data_cache.scala 67:29]
  reg  way1_dirty_126; // @[data_cache.scala 67:29]
  reg  way1_dirty_127; // @[data_cache.scala 67:29]
  reg [31:0] stage1_addr_line_mapping; // @[data_cache.scala 71:39]
  reg  stage1_sram_cache_reg; // @[data_cache.scala 72:40]
  reg [63:0] stage1_sram_wdata_reg; // @[data_cache.scala 73:40]
  reg [2:0] stage1_sram_size_reg; // @[data_cache.scala 74:39]
  reg  stage1_sram_wr_reg; // @[data_cache.scala 75:37]
  reg  stage1_sram_req_reg; // @[data_cache.scala 76:38]
  reg  stage1_sram_hit0_reg; // @[data_cache.scala 78:40]
  reg  stage1_sram_hit1_reg; // @[data_cache.scala 79:40]
  reg  stage1_sram_valid0_reg; // @[data_cache.scala 80:42]
  reg  stage1_sram_valid1_reg; // @[data_cache.scala 81:42]
  reg [7:0] stage1_wstrb_reg; // @[data_cache.scala 82:35]
  reg [31:0] stage1_sram_phy_addr_reg; // @[data_cache.scala 84:43]
  reg [7:0] data_write_back_counter; // @[data_cache.scala 146:42]
  wire  _data_cache_under_write_back_T = work_state == 5'h11; // @[data_cache.scala 148:51]
  wire  _data_cache_under_write_back_T_1 = work_state == 5'h15; // @[data_cache.scala 148:93]
  wire  _data_cache_under_write_back_T_3 = work_state == 5'h12; // @[data_cache.scala 148:135]
  wire  _data_cache_under_write_back_T_4 = work_state == 5'h11 | work_state == 5'h15 | work_state == 5'h12; // @[data_cache.scala 148:121]
  wire  _data_cache_under_write_back_T_5 = work_state == 5'h13; // @[data_cache.scala 149:23]
  wire  data_cache_under_write_back = _data_cache_under_write_back_T_4 | work_state == 5'h13 | work_state == 5'h14; // @[data_cache.scala 149:53]
  wire  _GEN_1 = 7'h1 == data_write_back_counter[6:0] ? way1_dirty_1 : way1_dirty_0; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_2 = 7'h2 == data_write_back_counter[6:0] ? way1_dirty_2 : _GEN_1; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_3 = 7'h3 == data_write_back_counter[6:0] ? way1_dirty_3 : _GEN_2; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_4 = 7'h4 == data_write_back_counter[6:0] ? way1_dirty_4 : _GEN_3; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_5 = 7'h5 == data_write_back_counter[6:0] ? way1_dirty_5 : _GEN_4; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_6 = 7'h6 == data_write_back_counter[6:0] ? way1_dirty_6 : _GEN_5; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_7 = 7'h7 == data_write_back_counter[6:0] ? way1_dirty_7 : _GEN_6; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_8 = 7'h8 == data_write_back_counter[6:0] ? way1_dirty_8 : _GEN_7; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_9 = 7'h9 == data_write_back_counter[6:0] ? way1_dirty_9 : _GEN_8; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_10 = 7'ha == data_write_back_counter[6:0] ? way1_dirty_10 : _GEN_9; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_11 = 7'hb == data_write_back_counter[6:0] ? way1_dirty_11 : _GEN_10; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_12 = 7'hc == data_write_back_counter[6:0] ? way1_dirty_12 : _GEN_11; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_13 = 7'hd == data_write_back_counter[6:0] ? way1_dirty_13 : _GEN_12; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_14 = 7'he == data_write_back_counter[6:0] ? way1_dirty_14 : _GEN_13; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_15 = 7'hf == data_write_back_counter[6:0] ? way1_dirty_15 : _GEN_14; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_16 = 7'h10 == data_write_back_counter[6:0] ? way1_dirty_16 : _GEN_15; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_17 = 7'h11 == data_write_back_counter[6:0] ? way1_dirty_17 : _GEN_16; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_18 = 7'h12 == data_write_back_counter[6:0] ? way1_dirty_18 : _GEN_17; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_19 = 7'h13 == data_write_back_counter[6:0] ? way1_dirty_19 : _GEN_18; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_20 = 7'h14 == data_write_back_counter[6:0] ? way1_dirty_20 : _GEN_19; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_21 = 7'h15 == data_write_back_counter[6:0] ? way1_dirty_21 : _GEN_20; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_22 = 7'h16 == data_write_back_counter[6:0] ? way1_dirty_22 : _GEN_21; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_23 = 7'h17 == data_write_back_counter[6:0] ? way1_dirty_23 : _GEN_22; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_24 = 7'h18 == data_write_back_counter[6:0] ? way1_dirty_24 : _GEN_23; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_25 = 7'h19 == data_write_back_counter[6:0] ? way1_dirty_25 : _GEN_24; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_26 = 7'h1a == data_write_back_counter[6:0] ? way1_dirty_26 : _GEN_25; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_27 = 7'h1b == data_write_back_counter[6:0] ? way1_dirty_27 : _GEN_26; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_28 = 7'h1c == data_write_back_counter[6:0] ? way1_dirty_28 : _GEN_27; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_29 = 7'h1d == data_write_back_counter[6:0] ? way1_dirty_29 : _GEN_28; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_30 = 7'h1e == data_write_back_counter[6:0] ? way1_dirty_30 : _GEN_29; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_31 = 7'h1f == data_write_back_counter[6:0] ? way1_dirty_31 : _GEN_30; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_32 = 7'h20 == data_write_back_counter[6:0] ? way1_dirty_32 : _GEN_31; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_33 = 7'h21 == data_write_back_counter[6:0] ? way1_dirty_33 : _GEN_32; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_34 = 7'h22 == data_write_back_counter[6:0] ? way1_dirty_34 : _GEN_33; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_35 = 7'h23 == data_write_back_counter[6:0] ? way1_dirty_35 : _GEN_34; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_36 = 7'h24 == data_write_back_counter[6:0] ? way1_dirty_36 : _GEN_35; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_37 = 7'h25 == data_write_back_counter[6:0] ? way1_dirty_37 : _GEN_36; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_38 = 7'h26 == data_write_back_counter[6:0] ? way1_dirty_38 : _GEN_37; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_39 = 7'h27 == data_write_back_counter[6:0] ? way1_dirty_39 : _GEN_38; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_40 = 7'h28 == data_write_back_counter[6:0] ? way1_dirty_40 : _GEN_39; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_41 = 7'h29 == data_write_back_counter[6:0] ? way1_dirty_41 : _GEN_40; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_42 = 7'h2a == data_write_back_counter[6:0] ? way1_dirty_42 : _GEN_41; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_43 = 7'h2b == data_write_back_counter[6:0] ? way1_dirty_43 : _GEN_42; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_44 = 7'h2c == data_write_back_counter[6:0] ? way1_dirty_44 : _GEN_43; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_45 = 7'h2d == data_write_back_counter[6:0] ? way1_dirty_45 : _GEN_44; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_46 = 7'h2e == data_write_back_counter[6:0] ? way1_dirty_46 : _GEN_45; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_47 = 7'h2f == data_write_back_counter[6:0] ? way1_dirty_47 : _GEN_46; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_48 = 7'h30 == data_write_back_counter[6:0] ? way1_dirty_48 : _GEN_47; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_49 = 7'h31 == data_write_back_counter[6:0] ? way1_dirty_49 : _GEN_48; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_50 = 7'h32 == data_write_back_counter[6:0] ? way1_dirty_50 : _GEN_49; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_51 = 7'h33 == data_write_back_counter[6:0] ? way1_dirty_51 : _GEN_50; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_52 = 7'h34 == data_write_back_counter[6:0] ? way1_dirty_52 : _GEN_51; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_53 = 7'h35 == data_write_back_counter[6:0] ? way1_dirty_53 : _GEN_52; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_54 = 7'h36 == data_write_back_counter[6:0] ? way1_dirty_54 : _GEN_53; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_55 = 7'h37 == data_write_back_counter[6:0] ? way1_dirty_55 : _GEN_54; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_56 = 7'h38 == data_write_back_counter[6:0] ? way1_dirty_56 : _GEN_55; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_57 = 7'h39 == data_write_back_counter[6:0] ? way1_dirty_57 : _GEN_56; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_58 = 7'h3a == data_write_back_counter[6:0] ? way1_dirty_58 : _GEN_57; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_59 = 7'h3b == data_write_back_counter[6:0] ? way1_dirty_59 : _GEN_58; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_60 = 7'h3c == data_write_back_counter[6:0] ? way1_dirty_60 : _GEN_59; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_61 = 7'h3d == data_write_back_counter[6:0] ? way1_dirty_61 : _GEN_60; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_62 = 7'h3e == data_write_back_counter[6:0] ? way1_dirty_62 : _GEN_61; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_63 = 7'h3f == data_write_back_counter[6:0] ? way1_dirty_63 : _GEN_62; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_64 = 7'h40 == data_write_back_counter[6:0] ? way1_dirty_64 : _GEN_63; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_65 = 7'h41 == data_write_back_counter[6:0] ? way1_dirty_65 : _GEN_64; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_66 = 7'h42 == data_write_back_counter[6:0] ? way1_dirty_66 : _GEN_65; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_67 = 7'h43 == data_write_back_counter[6:0] ? way1_dirty_67 : _GEN_66; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_68 = 7'h44 == data_write_back_counter[6:0] ? way1_dirty_68 : _GEN_67; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_69 = 7'h45 == data_write_back_counter[6:0] ? way1_dirty_69 : _GEN_68; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_70 = 7'h46 == data_write_back_counter[6:0] ? way1_dirty_70 : _GEN_69; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_71 = 7'h47 == data_write_back_counter[6:0] ? way1_dirty_71 : _GEN_70; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_72 = 7'h48 == data_write_back_counter[6:0] ? way1_dirty_72 : _GEN_71; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_73 = 7'h49 == data_write_back_counter[6:0] ? way1_dirty_73 : _GEN_72; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_74 = 7'h4a == data_write_back_counter[6:0] ? way1_dirty_74 : _GEN_73; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_75 = 7'h4b == data_write_back_counter[6:0] ? way1_dirty_75 : _GEN_74; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_76 = 7'h4c == data_write_back_counter[6:0] ? way1_dirty_76 : _GEN_75; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_77 = 7'h4d == data_write_back_counter[6:0] ? way1_dirty_77 : _GEN_76; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_78 = 7'h4e == data_write_back_counter[6:0] ? way1_dirty_78 : _GEN_77; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_79 = 7'h4f == data_write_back_counter[6:0] ? way1_dirty_79 : _GEN_78; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_80 = 7'h50 == data_write_back_counter[6:0] ? way1_dirty_80 : _GEN_79; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_81 = 7'h51 == data_write_back_counter[6:0] ? way1_dirty_81 : _GEN_80; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_82 = 7'h52 == data_write_back_counter[6:0] ? way1_dirty_82 : _GEN_81; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_83 = 7'h53 == data_write_back_counter[6:0] ? way1_dirty_83 : _GEN_82; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_84 = 7'h54 == data_write_back_counter[6:0] ? way1_dirty_84 : _GEN_83; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_85 = 7'h55 == data_write_back_counter[6:0] ? way1_dirty_85 : _GEN_84; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_86 = 7'h56 == data_write_back_counter[6:0] ? way1_dirty_86 : _GEN_85; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_87 = 7'h57 == data_write_back_counter[6:0] ? way1_dirty_87 : _GEN_86; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_88 = 7'h58 == data_write_back_counter[6:0] ? way1_dirty_88 : _GEN_87; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_89 = 7'h59 == data_write_back_counter[6:0] ? way1_dirty_89 : _GEN_88; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_90 = 7'h5a == data_write_back_counter[6:0] ? way1_dirty_90 : _GEN_89; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_91 = 7'h5b == data_write_back_counter[6:0] ? way1_dirty_91 : _GEN_90; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_92 = 7'h5c == data_write_back_counter[6:0] ? way1_dirty_92 : _GEN_91; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_93 = 7'h5d == data_write_back_counter[6:0] ? way1_dirty_93 : _GEN_92; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_94 = 7'h5e == data_write_back_counter[6:0] ? way1_dirty_94 : _GEN_93; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_95 = 7'h5f == data_write_back_counter[6:0] ? way1_dirty_95 : _GEN_94; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_96 = 7'h60 == data_write_back_counter[6:0] ? way1_dirty_96 : _GEN_95; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_97 = 7'h61 == data_write_back_counter[6:0] ? way1_dirty_97 : _GEN_96; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_98 = 7'h62 == data_write_back_counter[6:0] ? way1_dirty_98 : _GEN_97; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_99 = 7'h63 == data_write_back_counter[6:0] ? way1_dirty_99 : _GEN_98; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_100 = 7'h64 == data_write_back_counter[6:0] ? way1_dirty_100 : _GEN_99; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_101 = 7'h65 == data_write_back_counter[6:0] ? way1_dirty_101 : _GEN_100; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_102 = 7'h66 == data_write_back_counter[6:0] ? way1_dirty_102 : _GEN_101; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_103 = 7'h67 == data_write_back_counter[6:0] ? way1_dirty_103 : _GEN_102; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_104 = 7'h68 == data_write_back_counter[6:0] ? way1_dirty_104 : _GEN_103; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_105 = 7'h69 == data_write_back_counter[6:0] ? way1_dirty_105 : _GEN_104; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_106 = 7'h6a == data_write_back_counter[6:0] ? way1_dirty_106 : _GEN_105; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_107 = 7'h6b == data_write_back_counter[6:0] ? way1_dirty_107 : _GEN_106; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_108 = 7'h6c == data_write_back_counter[6:0] ? way1_dirty_108 : _GEN_107; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_109 = 7'h6d == data_write_back_counter[6:0] ? way1_dirty_109 : _GEN_108; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_110 = 7'h6e == data_write_back_counter[6:0] ? way1_dirty_110 : _GEN_109; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_111 = 7'h6f == data_write_back_counter[6:0] ? way1_dirty_111 : _GEN_110; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_112 = 7'h70 == data_write_back_counter[6:0] ? way1_dirty_112 : _GEN_111; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_113 = 7'h71 == data_write_back_counter[6:0] ? way1_dirty_113 : _GEN_112; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_114 = 7'h72 == data_write_back_counter[6:0] ? way1_dirty_114 : _GEN_113; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_115 = 7'h73 == data_write_back_counter[6:0] ? way1_dirty_115 : _GEN_114; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_116 = 7'h74 == data_write_back_counter[6:0] ? way1_dirty_116 : _GEN_115; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_117 = 7'h75 == data_write_back_counter[6:0] ? way1_dirty_117 : _GEN_116; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_118 = 7'h76 == data_write_back_counter[6:0] ? way1_dirty_118 : _GEN_117; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_119 = 7'h77 == data_write_back_counter[6:0] ? way1_dirty_119 : _GEN_118; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_120 = 7'h78 == data_write_back_counter[6:0] ? way1_dirty_120 : _GEN_119; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_121 = 7'h79 == data_write_back_counter[6:0] ? way1_dirty_121 : _GEN_120; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_122 = 7'h7a == data_write_back_counter[6:0] ? way1_dirty_122 : _GEN_121; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_123 = 7'h7b == data_write_back_counter[6:0] ? way1_dirty_123 : _GEN_122; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_124 = 7'h7c == data_write_back_counter[6:0] ? way1_dirty_124 : _GEN_123; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_125 = 7'h7d == data_write_back_counter[6:0] ? way1_dirty_125 : _GEN_124; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_126 = 7'h7e == data_write_back_counter[6:0] ? way1_dirty_126 : _GEN_125; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_127 = 7'h7f == data_write_back_counter[6:0] ? way1_dirty_127 : _GEN_126; // @[data_cache.scala 159:{149,149}]
  wire  _GEN_129 = 7'h1 == data_write_back_counter[6:0] ? way0_dirty_1 : way0_dirty_0; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_130 = 7'h2 == data_write_back_counter[6:0] ? way0_dirty_2 : _GEN_129; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_131 = 7'h3 == data_write_back_counter[6:0] ? way0_dirty_3 : _GEN_130; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_132 = 7'h4 == data_write_back_counter[6:0] ? way0_dirty_4 : _GEN_131; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_133 = 7'h5 == data_write_back_counter[6:0] ? way0_dirty_5 : _GEN_132; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_134 = 7'h6 == data_write_back_counter[6:0] ? way0_dirty_6 : _GEN_133; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_135 = 7'h7 == data_write_back_counter[6:0] ? way0_dirty_7 : _GEN_134; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_136 = 7'h8 == data_write_back_counter[6:0] ? way0_dirty_8 : _GEN_135; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_137 = 7'h9 == data_write_back_counter[6:0] ? way0_dirty_9 : _GEN_136; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_138 = 7'ha == data_write_back_counter[6:0] ? way0_dirty_10 : _GEN_137; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_139 = 7'hb == data_write_back_counter[6:0] ? way0_dirty_11 : _GEN_138; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_140 = 7'hc == data_write_back_counter[6:0] ? way0_dirty_12 : _GEN_139; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_141 = 7'hd == data_write_back_counter[6:0] ? way0_dirty_13 : _GEN_140; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_142 = 7'he == data_write_back_counter[6:0] ? way0_dirty_14 : _GEN_141; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_143 = 7'hf == data_write_back_counter[6:0] ? way0_dirty_15 : _GEN_142; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_144 = 7'h10 == data_write_back_counter[6:0] ? way0_dirty_16 : _GEN_143; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_145 = 7'h11 == data_write_back_counter[6:0] ? way0_dirty_17 : _GEN_144; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_146 = 7'h12 == data_write_back_counter[6:0] ? way0_dirty_18 : _GEN_145; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_147 = 7'h13 == data_write_back_counter[6:0] ? way0_dirty_19 : _GEN_146; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_148 = 7'h14 == data_write_back_counter[6:0] ? way0_dirty_20 : _GEN_147; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_149 = 7'h15 == data_write_back_counter[6:0] ? way0_dirty_21 : _GEN_148; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_150 = 7'h16 == data_write_back_counter[6:0] ? way0_dirty_22 : _GEN_149; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_151 = 7'h17 == data_write_back_counter[6:0] ? way0_dirty_23 : _GEN_150; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_152 = 7'h18 == data_write_back_counter[6:0] ? way0_dirty_24 : _GEN_151; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_153 = 7'h19 == data_write_back_counter[6:0] ? way0_dirty_25 : _GEN_152; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_154 = 7'h1a == data_write_back_counter[6:0] ? way0_dirty_26 : _GEN_153; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_155 = 7'h1b == data_write_back_counter[6:0] ? way0_dirty_27 : _GEN_154; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_156 = 7'h1c == data_write_back_counter[6:0] ? way0_dirty_28 : _GEN_155; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_157 = 7'h1d == data_write_back_counter[6:0] ? way0_dirty_29 : _GEN_156; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_158 = 7'h1e == data_write_back_counter[6:0] ? way0_dirty_30 : _GEN_157; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_159 = 7'h1f == data_write_back_counter[6:0] ? way0_dirty_31 : _GEN_158; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_160 = 7'h20 == data_write_back_counter[6:0] ? way0_dirty_32 : _GEN_159; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_161 = 7'h21 == data_write_back_counter[6:0] ? way0_dirty_33 : _GEN_160; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_162 = 7'h22 == data_write_back_counter[6:0] ? way0_dirty_34 : _GEN_161; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_163 = 7'h23 == data_write_back_counter[6:0] ? way0_dirty_35 : _GEN_162; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_164 = 7'h24 == data_write_back_counter[6:0] ? way0_dirty_36 : _GEN_163; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_165 = 7'h25 == data_write_back_counter[6:0] ? way0_dirty_37 : _GEN_164; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_166 = 7'h26 == data_write_back_counter[6:0] ? way0_dirty_38 : _GEN_165; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_167 = 7'h27 == data_write_back_counter[6:0] ? way0_dirty_39 : _GEN_166; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_168 = 7'h28 == data_write_back_counter[6:0] ? way0_dirty_40 : _GEN_167; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_169 = 7'h29 == data_write_back_counter[6:0] ? way0_dirty_41 : _GEN_168; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_170 = 7'h2a == data_write_back_counter[6:0] ? way0_dirty_42 : _GEN_169; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_171 = 7'h2b == data_write_back_counter[6:0] ? way0_dirty_43 : _GEN_170; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_172 = 7'h2c == data_write_back_counter[6:0] ? way0_dirty_44 : _GEN_171; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_173 = 7'h2d == data_write_back_counter[6:0] ? way0_dirty_45 : _GEN_172; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_174 = 7'h2e == data_write_back_counter[6:0] ? way0_dirty_46 : _GEN_173; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_175 = 7'h2f == data_write_back_counter[6:0] ? way0_dirty_47 : _GEN_174; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_176 = 7'h30 == data_write_back_counter[6:0] ? way0_dirty_48 : _GEN_175; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_177 = 7'h31 == data_write_back_counter[6:0] ? way0_dirty_49 : _GEN_176; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_178 = 7'h32 == data_write_back_counter[6:0] ? way0_dirty_50 : _GEN_177; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_179 = 7'h33 == data_write_back_counter[6:0] ? way0_dirty_51 : _GEN_178; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_180 = 7'h34 == data_write_back_counter[6:0] ? way0_dirty_52 : _GEN_179; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_181 = 7'h35 == data_write_back_counter[6:0] ? way0_dirty_53 : _GEN_180; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_182 = 7'h36 == data_write_back_counter[6:0] ? way0_dirty_54 : _GEN_181; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_183 = 7'h37 == data_write_back_counter[6:0] ? way0_dirty_55 : _GEN_182; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_184 = 7'h38 == data_write_back_counter[6:0] ? way0_dirty_56 : _GEN_183; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_185 = 7'h39 == data_write_back_counter[6:0] ? way0_dirty_57 : _GEN_184; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_186 = 7'h3a == data_write_back_counter[6:0] ? way0_dirty_58 : _GEN_185; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_187 = 7'h3b == data_write_back_counter[6:0] ? way0_dirty_59 : _GEN_186; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_188 = 7'h3c == data_write_back_counter[6:0] ? way0_dirty_60 : _GEN_187; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_189 = 7'h3d == data_write_back_counter[6:0] ? way0_dirty_61 : _GEN_188; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_190 = 7'h3e == data_write_back_counter[6:0] ? way0_dirty_62 : _GEN_189; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_191 = 7'h3f == data_write_back_counter[6:0] ? way0_dirty_63 : _GEN_190; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_192 = 7'h40 == data_write_back_counter[6:0] ? way0_dirty_64 : _GEN_191; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_193 = 7'h41 == data_write_back_counter[6:0] ? way0_dirty_65 : _GEN_192; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_194 = 7'h42 == data_write_back_counter[6:0] ? way0_dirty_66 : _GEN_193; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_195 = 7'h43 == data_write_back_counter[6:0] ? way0_dirty_67 : _GEN_194; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_196 = 7'h44 == data_write_back_counter[6:0] ? way0_dirty_68 : _GEN_195; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_197 = 7'h45 == data_write_back_counter[6:0] ? way0_dirty_69 : _GEN_196; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_198 = 7'h46 == data_write_back_counter[6:0] ? way0_dirty_70 : _GEN_197; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_199 = 7'h47 == data_write_back_counter[6:0] ? way0_dirty_71 : _GEN_198; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_200 = 7'h48 == data_write_back_counter[6:0] ? way0_dirty_72 : _GEN_199; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_201 = 7'h49 == data_write_back_counter[6:0] ? way0_dirty_73 : _GEN_200; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_202 = 7'h4a == data_write_back_counter[6:0] ? way0_dirty_74 : _GEN_201; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_203 = 7'h4b == data_write_back_counter[6:0] ? way0_dirty_75 : _GEN_202; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_204 = 7'h4c == data_write_back_counter[6:0] ? way0_dirty_76 : _GEN_203; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_205 = 7'h4d == data_write_back_counter[6:0] ? way0_dirty_77 : _GEN_204; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_206 = 7'h4e == data_write_back_counter[6:0] ? way0_dirty_78 : _GEN_205; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_207 = 7'h4f == data_write_back_counter[6:0] ? way0_dirty_79 : _GEN_206; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_208 = 7'h50 == data_write_back_counter[6:0] ? way0_dirty_80 : _GEN_207; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_209 = 7'h51 == data_write_back_counter[6:0] ? way0_dirty_81 : _GEN_208; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_210 = 7'h52 == data_write_back_counter[6:0] ? way0_dirty_82 : _GEN_209; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_211 = 7'h53 == data_write_back_counter[6:0] ? way0_dirty_83 : _GEN_210; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_212 = 7'h54 == data_write_back_counter[6:0] ? way0_dirty_84 : _GEN_211; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_213 = 7'h55 == data_write_back_counter[6:0] ? way0_dirty_85 : _GEN_212; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_214 = 7'h56 == data_write_back_counter[6:0] ? way0_dirty_86 : _GEN_213; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_215 = 7'h57 == data_write_back_counter[6:0] ? way0_dirty_87 : _GEN_214; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_216 = 7'h58 == data_write_back_counter[6:0] ? way0_dirty_88 : _GEN_215; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_217 = 7'h59 == data_write_back_counter[6:0] ? way0_dirty_89 : _GEN_216; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_218 = 7'h5a == data_write_back_counter[6:0] ? way0_dirty_90 : _GEN_217; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_219 = 7'h5b == data_write_back_counter[6:0] ? way0_dirty_91 : _GEN_218; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_220 = 7'h5c == data_write_back_counter[6:0] ? way0_dirty_92 : _GEN_219; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_221 = 7'h5d == data_write_back_counter[6:0] ? way0_dirty_93 : _GEN_220; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_222 = 7'h5e == data_write_back_counter[6:0] ? way0_dirty_94 : _GEN_221; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_223 = 7'h5f == data_write_back_counter[6:0] ? way0_dirty_95 : _GEN_222; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_224 = 7'h60 == data_write_back_counter[6:0] ? way0_dirty_96 : _GEN_223; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_225 = 7'h61 == data_write_back_counter[6:0] ? way0_dirty_97 : _GEN_224; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_226 = 7'h62 == data_write_back_counter[6:0] ? way0_dirty_98 : _GEN_225; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_227 = 7'h63 == data_write_back_counter[6:0] ? way0_dirty_99 : _GEN_226; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_228 = 7'h64 == data_write_back_counter[6:0] ? way0_dirty_100 : _GEN_227; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_229 = 7'h65 == data_write_back_counter[6:0] ? way0_dirty_101 : _GEN_228; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_230 = 7'h66 == data_write_back_counter[6:0] ? way0_dirty_102 : _GEN_229; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_231 = 7'h67 == data_write_back_counter[6:0] ? way0_dirty_103 : _GEN_230; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_232 = 7'h68 == data_write_back_counter[6:0] ? way0_dirty_104 : _GEN_231; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_233 = 7'h69 == data_write_back_counter[6:0] ? way0_dirty_105 : _GEN_232; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_234 = 7'h6a == data_write_back_counter[6:0] ? way0_dirty_106 : _GEN_233; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_235 = 7'h6b == data_write_back_counter[6:0] ? way0_dirty_107 : _GEN_234; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_236 = 7'h6c == data_write_back_counter[6:0] ? way0_dirty_108 : _GEN_235; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_237 = 7'h6d == data_write_back_counter[6:0] ? way0_dirty_109 : _GEN_236; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_238 = 7'h6e == data_write_back_counter[6:0] ? way0_dirty_110 : _GEN_237; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_239 = 7'h6f == data_write_back_counter[6:0] ? way0_dirty_111 : _GEN_238; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_240 = 7'h70 == data_write_back_counter[6:0] ? way0_dirty_112 : _GEN_239; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_241 = 7'h71 == data_write_back_counter[6:0] ? way0_dirty_113 : _GEN_240; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_242 = 7'h72 == data_write_back_counter[6:0] ? way0_dirty_114 : _GEN_241; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_243 = 7'h73 == data_write_back_counter[6:0] ? way0_dirty_115 : _GEN_242; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_244 = 7'h74 == data_write_back_counter[6:0] ? way0_dirty_116 : _GEN_243; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_245 = 7'h75 == data_write_back_counter[6:0] ? way0_dirty_117 : _GEN_244; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_246 = 7'h76 == data_write_back_counter[6:0] ? way0_dirty_118 : _GEN_245; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_247 = 7'h77 == data_write_back_counter[6:0] ? way0_dirty_119 : _GEN_246; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_248 = 7'h78 == data_write_back_counter[6:0] ? way0_dirty_120 : _GEN_247; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_249 = 7'h79 == data_write_back_counter[6:0] ? way0_dirty_121 : _GEN_248; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_250 = 7'h7a == data_write_back_counter[6:0] ? way0_dirty_122 : _GEN_249; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_251 = 7'h7b == data_write_back_counter[6:0] ? way0_dirty_123 : _GEN_250; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_252 = 7'h7c == data_write_back_counter[6:0] ? way0_dirty_124 : _GEN_251; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_253 = 7'h7d == data_write_back_counter[6:0] ? way0_dirty_125 : _GEN_252; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_254 = 7'h7e == data_write_back_counter[6:0] ? way0_dirty_126 : _GEN_253; // @[data_cache.scala 160:{87,87}]
  wire  _GEN_255 = 7'h7f == data_write_back_counter[6:0] ? way0_dirty_127 : _GEN_254; // @[data_cache.scala 160:{87,87}]
  wire  _data_should_write_back_T_6 = dcache_tag_io_w_valid & _GEN_255; // @[data_cache.scala 160:30]
  wire  data_should_write_back = data_write_back_counter[7] ? dcache_tag_1_io_w_valid & _GEN_127 :
    _data_should_write_back_T_6; // @[data_cache.scala 159:34]
  wire  _data_write_back_counter_T_2 = _data_cache_under_write_back_T & ~data_should_write_back; // @[data_cache.scala 153:49]
  wire [7:0] _data_write_back_counter_T_4 = data_write_back_counter + 8'h1; // @[data_cache.scala 153:106]
  wire  data_all_write_back = data_write_back_counter == 8'hff; // @[data_cache.scala 158:55]
  wire  _hit_T = stage1_sram_hit0_reg & stage1_sram_valid0_reg; // @[data_cache.scala 238:37]
  wire  _hit_T_1 = stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 239:31]
  wire  hit = stage1_sram_hit0_reg & stage1_sram_valid0_reg | _hit_T_1; // @[data_cache.scala 238:64]
  wire [4:0] _state_ready_lookup_should_be_T_2 = stage1_sram_cache_reg ? 5'h19 : 5'h0; // @[data_cache.scala 249:82]
  wire [4:0] _state_ready_lookup_should_be_T_3 = stage1_sram_req_reg ? _state_ready_lookup_should_be_T_2 : 5'h19; // @[data_cache.scala 249:51]
  wire [4:0] _state_ready_lookup_should_be_T_5 = stage1_sram_req_reg ? 5'h0 : 5'h19; // @[data_cache.scala 250:16]
  wire [4:0] state_ready_lookup_should_be = hit ? _state_ready_lookup_should_be_T_3 : _state_ready_lookup_should_be_T_5; // @[data_cache.scala 249:43]
  wire [1:0] _access_work_state_for_stall_T_6 = io_port_bvalid ? 2'h3 : 2'h0; // @[data_cache.scala 286:40]
  wire [1:0] _access_work_state_for_stall_T_3 = io_port_rvalid ? 2'h3 : work_state[4:3]; // @[data_cache.scala 284:39]
  wire [1:0] _access_work_state_for_stall_T_9 = 5'h2 == work_state ? _access_work_state_for_stall_T_3 : work_state[4:3]; // @[Mux.scala 81:58]
  wire [1:0] _access_work_state_for_stall_T_11 = 5'h18 == work_state ? state_ready_lookup_should_be[4:3] :
    _access_work_state_for_stall_T_9; // @[Mux.scala 81:58]
  wire [1:0] _access_work_state_for_stall_T_13 = 5'h5 == work_state ? _access_work_state_for_stall_T_6 :
    _access_work_state_for_stall_T_11; // @[Mux.scala 81:58]
  wire [1:0] _access_work_state_for_stall_T_15 = 5'h19 == work_state ? state_ready_lookup_should_be[4:3] :
    _access_work_state_for_stall_T_13; // @[Mux.scala 81:58]
  wire [1:0] _access_work_state_for_stall_T_17 = 5'he == work_state ? 2'h3 : _access_work_state_for_stall_T_15; // @[Mux.scala 81:58]
  wire [1:0] access_work_state_for_stall = 5'h10 == work_state ? 2'h3 : _access_work_state_for_stall_T_17; // @[Mux.scala 81:58]
  wire  stage2_stall = access_work_state_for_stall == 2'h3; // @[data_cache.scala 295:48]
  reg  stage2_sram_write_reg; // @[data_cache.scala 176:40]
  reg  stage1_stall_reg; // @[data_cache.scala 183:35]
  reg  write_access_complete_reg; // @[data_cache.scala 186:44]
  wire  _stage1_sram_req_reg_T_1 = stage2_stall ? 1'h0 : stage1_sram_req_reg; // @[data_cache.scala 195:60]
  wire [4:0] _state_lookup_for_less_delay_T_1 = 5'h18 == work_state ? state_ready_lookup_should_be : work_state; // @[Mux.scala 81:58]
  wire [4:0] state_lookup_for_less_delay = 5'h19 == work_state ? state_ready_lookup_should_be :
    _state_lookup_for_less_delay_T_1; // @[Mux.scala 81:58]
  wire  _way0_dirty_T = state_lookup_for_less_delay == 5'h19; // @[data_cache.scala 204:79]
  wire  _way0_dirty_T_2 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg; // @[data_cache.scala 204:96]
  wire  _way0_dirty_T_4 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
    stage1_sram_valid0_reg; // @[data_cache.scala 204:149]
  wire  _way0_dirty_T_5 = work_state == 5'he; // @[data_cache.scala 205:24]
  wire  _GEN_258 = 7'h1 == stage1_addr_line_mapping[10:4] ? lru_1 : lru_0; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_259 = 7'h2 == stage1_addr_line_mapping[10:4] ? lru_2 : _GEN_258; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_260 = 7'h3 == stage1_addr_line_mapping[10:4] ? lru_3 : _GEN_259; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_261 = 7'h4 == stage1_addr_line_mapping[10:4] ? lru_4 : _GEN_260; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_262 = 7'h5 == stage1_addr_line_mapping[10:4] ? lru_5 : _GEN_261; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_263 = 7'h6 == stage1_addr_line_mapping[10:4] ? lru_6 : _GEN_262; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_264 = 7'h7 == stage1_addr_line_mapping[10:4] ? lru_7 : _GEN_263; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_265 = 7'h8 == stage1_addr_line_mapping[10:4] ? lru_8 : _GEN_264; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_266 = 7'h9 == stage1_addr_line_mapping[10:4] ? lru_9 : _GEN_265; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_267 = 7'ha == stage1_addr_line_mapping[10:4] ? lru_10 : _GEN_266; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_268 = 7'hb == stage1_addr_line_mapping[10:4] ? lru_11 : _GEN_267; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_269 = 7'hc == stage1_addr_line_mapping[10:4] ? lru_12 : _GEN_268; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_270 = 7'hd == stage1_addr_line_mapping[10:4] ? lru_13 : _GEN_269; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_271 = 7'he == stage1_addr_line_mapping[10:4] ? lru_14 : _GEN_270; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_272 = 7'hf == stage1_addr_line_mapping[10:4] ? lru_15 : _GEN_271; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_273 = 7'h10 == stage1_addr_line_mapping[10:4] ? lru_16 : _GEN_272; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_274 = 7'h11 == stage1_addr_line_mapping[10:4] ? lru_17 : _GEN_273; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_275 = 7'h12 == stage1_addr_line_mapping[10:4] ? lru_18 : _GEN_274; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_276 = 7'h13 == stage1_addr_line_mapping[10:4] ? lru_19 : _GEN_275; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_277 = 7'h14 == stage1_addr_line_mapping[10:4] ? lru_20 : _GEN_276; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_278 = 7'h15 == stage1_addr_line_mapping[10:4] ? lru_21 : _GEN_277; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_279 = 7'h16 == stage1_addr_line_mapping[10:4] ? lru_22 : _GEN_278; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_280 = 7'h17 == stage1_addr_line_mapping[10:4] ? lru_23 : _GEN_279; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_281 = 7'h18 == stage1_addr_line_mapping[10:4] ? lru_24 : _GEN_280; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_282 = 7'h19 == stage1_addr_line_mapping[10:4] ? lru_25 : _GEN_281; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_283 = 7'h1a == stage1_addr_line_mapping[10:4] ? lru_26 : _GEN_282; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_284 = 7'h1b == stage1_addr_line_mapping[10:4] ? lru_27 : _GEN_283; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_285 = 7'h1c == stage1_addr_line_mapping[10:4] ? lru_28 : _GEN_284; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_286 = 7'h1d == stage1_addr_line_mapping[10:4] ? lru_29 : _GEN_285; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_287 = 7'h1e == stage1_addr_line_mapping[10:4] ? lru_30 : _GEN_286; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_288 = 7'h1f == stage1_addr_line_mapping[10:4] ? lru_31 : _GEN_287; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_289 = 7'h20 == stage1_addr_line_mapping[10:4] ? lru_32 : _GEN_288; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_290 = 7'h21 == stage1_addr_line_mapping[10:4] ? lru_33 : _GEN_289; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_291 = 7'h22 == stage1_addr_line_mapping[10:4] ? lru_34 : _GEN_290; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_292 = 7'h23 == stage1_addr_line_mapping[10:4] ? lru_35 : _GEN_291; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_293 = 7'h24 == stage1_addr_line_mapping[10:4] ? lru_36 : _GEN_292; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_294 = 7'h25 == stage1_addr_line_mapping[10:4] ? lru_37 : _GEN_293; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_295 = 7'h26 == stage1_addr_line_mapping[10:4] ? lru_38 : _GEN_294; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_296 = 7'h27 == stage1_addr_line_mapping[10:4] ? lru_39 : _GEN_295; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_297 = 7'h28 == stage1_addr_line_mapping[10:4] ? lru_40 : _GEN_296; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_298 = 7'h29 == stage1_addr_line_mapping[10:4] ? lru_41 : _GEN_297; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_299 = 7'h2a == stage1_addr_line_mapping[10:4] ? lru_42 : _GEN_298; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_300 = 7'h2b == stage1_addr_line_mapping[10:4] ? lru_43 : _GEN_299; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_301 = 7'h2c == stage1_addr_line_mapping[10:4] ? lru_44 : _GEN_300; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_302 = 7'h2d == stage1_addr_line_mapping[10:4] ? lru_45 : _GEN_301; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_303 = 7'h2e == stage1_addr_line_mapping[10:4] ? lru_46 : _GEN_302; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_304 = 7'h2f == stage1_addr_line_mapping[10:4] ? lru_47 : _GEN_303; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_305 = 7'h30 == stage1_addr_line_mapping[10:4] ? lru_48 : _GEN_304; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_306 = 7'h31 == stage1_addr_line_mapping[10:4] ? lru_49 : _GEN_305; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_307 = 7'h32 == stage1_addr_line_mapping[10:4] ? lru_50 : _GEN_306; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_308 = 7'h33 == stage1_addr_line_mapping[10:4] ? lru_51 : _GEN_307; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_309 = 7'h34 == stage1_addr_line_mapping[10:4] ? lru_52 : _GEN_308; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_310 = 7'h35 == stage1_addr_line_mapping[10:4] ? lru_53 : _GEN_309; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_311 = 7'h36 == stage1_addr_line_mapping[10:4] ? lru_54 : _GEN_310; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_312 = 7'h37 == stage1_addr_line_mapping[10:4] ? lru_55 : _GEN_311; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_313 = 7'h38 == stage1_addr_line_mapping[10:4] ? lru_56 : _GEN_312; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_314 = 7'h39 == stage1_addr_line_mapping[10:4] ? lru_57 : _GEN_313; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_315 = 7'h3a == stage1_addr_line_mapping[10:4] ? lru_58 : _GEN_314; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_316 = 7'h3b == stage1_addr_line_mapping[10:4] ? lru_59 : _GEN_315; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_317 = 7'h3c == stage1_addr_line_mapping[10:4] ? lru_60 : _GEN_316; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_318 = 7'h3d == stage1_addr_line_mapping[10:4] ? lru_61 : _GEN_317; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_319 = 7'h3e == stage1_addr_line_mapping[10:4] ? lru_62 : _GEN_318; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_320 = 7'h3f == stage1_addr_line_mapping[10:4] ? lru_63 : _GEN_319; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_321 = 7'h40 == stage1_addr_line_mapping[10:4] ? lru_64 : _GEN_320; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_322 = 7'h41 == stage1_addr_line_mapping[10:4] ? lru_65 : _GEN_321; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_323 = 7'h42 == stage1_addr_line_mapping[10:4] ? lru_66 : _GEN_322; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_324 = 7'h43 == stage1_addr_line_mapping[10:4] ? lru_67 : _GEN_323; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_325 = 7'h44 == stage1_addr_line_mapping[10:4] ? lru_68 : _GEN_324; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_326 = 7'h45 == stage1_addr_line_mapping[10:4] ? lru_69 : _GEN_325; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_327 = 7'h46 == stage1_addr_line_mapping[10:4] ? lru_70 : _GEN_326; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_328 = 7'h47 == stage1_addr_line_mapping[10:4] ? lru_71 : _GEN_327; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_329 = 7'h48 == stage1_addr_line_mapping[10:4] ? lru_72 : _GEN_328; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_330 = 7'h49 == stage1_addr_line_mapping[10:4] ? lru_73 : _GEN_329; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_331 = 7'h4a == stage1_addr_line_mapping[10:4] ? lru_74 : _GEN_330; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_332 = 7'h4b == stage1_addr_line_mapping[10:4] ? lru_75 : _GEN_331; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_333 = 7'h4c == stage1_addr_line_mapping[10:4] ? lru_76 : _GEN_332; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_334 = 7'h4d == stage1_addr_line_mapping[10:4] ? lru_77 : _GEN_333; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_335 = 7'h4e == stage1_addr_line_mapping[10:4] ? lru_78 : _GEN_334; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_336 = 7'h4f == stage1_addr_line_mapping[10:4] ? lru_79 : _GEN_335; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_337 = 7'h50 == stage1_addr_line_mapping[10:4] ? lru_80 : _GEN_336; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_338 = 7'h51 == stage1_addr_line_mapping[10:4] ? lru_81 : _GEN_337; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_339 = 7'h52 == stage1_addr_line_mapping[10:4] ? lru_82 : _GEN_338; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_340 = 7'h53 == stage1_addr_line_mapping[10:4] ? lru_83 : _GEN_339; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_341 = 7'h54 == stage1_addr_line_mapping[10:4] ? lru_84 : _GEN_340; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_342 = 7'h55 == stage1_addr_line_mapping[10:4] ? lru_85 : _GEN_341; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_343 = 7'h56 == stage1_addr_line_mapping[10:4] ? lru_86 : _GEN_342; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_344 = 7'h57 == stage1_addr_line_mapping[10:4] ? lru_87 : _GEN_343; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_345 = 7'h58 == stage1_addr_line_mapping[10:4] ? lru_88 : _GEN_344; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_346 = 7'h59 == stage1_addr_line_mapping[10:4] ? lru_89 : _GEN_345; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_347 = 7'h5a == stage1_addr_line_mapping[10:4] ? lru_90 : _GEN_346; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_348 = 7'h5b == stage1_addr_line_mapping[10:4] ? lru_91 : _GEN_347; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_349 = 7'h5c == stage1_addr_line_mapping[10:4] ? lru_92 : _GEN_348; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_350 = 7'h5d == stage1_addr_line_mapping[10:4] ? lru_93 : _GEN_349; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_351 = 7'h5e == stage1_addr_line_mapping[10:4] ? lru_94 : _GEN_350; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_352 = 7'h5f == stage1_addr_line_mapping[10:4] ? lru_95 : _GEN_351; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_353 = 7'h60 == stage1_addr_line_mapping[10:4] ? lru_96 : _GEN_352; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_354 = 7'h61 == stage1_addr_line_mapping[10:4] ? lru_97 : _GEN_353; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_355 = 7'h62 == stage1_addr_line_mapping[10:4] ? lru_98 : _GEN_354; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_356 = 7'h63 == stage1_addr_line_mapping[10:4] ? lru_99 : _GEN_355; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_357 = 7'h64 == stage1_addr_line_mapping[10:4] ? lru_100 : _GEN_356; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_358 = 7'h65 == stage1_addr_line_mapping[10:4] ? lru_101 : _GEN_357; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_359 = 7'h66 == stage1_addr_line_mapping[10:4] ? lru_102 : _GEN_358; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_360 = 7'h67 == stage1_addr_line_mapping[10:4] ? lru_103 : _GEN_359; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_361 = 7'h68 == stage1_addr_line_mapping[10:4] ? lru_104 : _GEN_360; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_362 = 7'h69 == stage1_addr_line_mapping[10:4] ? lru_105 : _GEN_361; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_363 = 7'h6a == stage1_addr_line_mapping[10:4] ? lru_106 : _GEN_362; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_364 = 7'h6b == stage1_addr_line_mapping[10:4] ? lru_107 : _GEN_363; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_365 = 7'h6c == stage1_addr_line_mapping[10:4] ? lru_108 : _GEN_364; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_366 = 7'h6d == stage1_addr_line_mapping[10:4] ? lru_109 : _GEN_365; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_367 = 7'h6e == stage1_addr_line_mapping[10:4] ? lru_110 : _GEN_366; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_368 = 7'h6f == stage1_addr_line_mapping[10:4] ? lru_111 : _GEN_367; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_369 = 7'h70 == stage1_addr_line_mapping[10:4] ? lru_112 : _GEN_368; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_370 = 7'h71 == stage1_addr_line_mapping[10:4] ? lru_113 : _GEN_369; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_371 = 7'h72 == stage1_addr_line_mapping[10:4] ? lru_114 : _GEN_370; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_372 = 7'h73 == stage1_addr_line_mapping[10:4] ? lru_115 : _GEN_371; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_373 = 7'h74 == stage1_addr_line_mapping[10:4] ? lru_116 : _GEN_372; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_374 = 7'h75 == stage1_addr_line_mapping[10:4] ? lru_117 : _GEN_373; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_375 = 7'h76 == stage1_addr_line_mapping[10:4] ? lru_118 : _GEN_374; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_376 = 7'h77 == stage1_addr_line_mapping[10:4] ? lru_119 : _GEN_375; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_377 = 7'h78 == stage1_addr_line_mapping[10:4] ? lru_120 : _GEN_376; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_378 = 7'h79 == stage1_addr_line_mapping[10:4] ? lru_121 : _GEN_377; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_379 = 7'h7a == stage1_addr_line_mapping[10:4] ? lru_122 : _GEN_378; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_380 = 7'h7b == stage1_addr_line_mapping[10:4] ? lru_123 : _GEN_379; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_381 = 7'h7c == stage1_addr_line_mapping[10:4] ? lru_124 : _GEN_380; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_382 = 7'h7d == stage1_addr_line_mapping[10:4] ? lru_125 : _GEN_381; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_383 = 7'h7e == stage1_addr_line_mapping[10:4] ? lru_126 : _GEN_382; // @[data_cache.scala 205:{86,86}]
  wire  _GEN_384 = 7'h7f == stage1_addr_line_mapping[10:4] ? lru_127 : _GEN_383; // @[data_cache.scala 205:{86,86}]
  wire  _way0_dirty_T_7 = ~_GEN_384; // @[data_cache.scala 205:86]
  wire  _way0_dirty_T_9 = work_state == 5'h10; // @[data_cache.scala 206:24]
  wire  _way0_dirty_T_12 = work_state == 5'h10 & _way0_dirty_T_7; // @[data_cache.scala 206:52]
  wire  _GEN_514 = 7'h1 == stage1_addr_line_mapping[10:4] ? way0_dirty_1 : way0_dirty_0; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_515 = 7'h2 == stage1_addr_line_mapping[10:4] ? way0_dirty_2 : _GEN_514; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_516 = 7'h3 == stage1_addr_line_mapping[10:4] ? way0_dirty_3 : _GEN_515; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_517 = 7'h4 == stage1_addr_line_mapping[10:4] ? way0_dirty_4 : _GEN_516; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_518 = 7'h5 == stage1_addr_line_mapping[10:4] ? way0_dirty_5 : _GEN_517; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_519 = 7'h6 == stage1_addr_line_mapping[10:4] ? way0_dirty_6 : _GEN_518; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_520 = 7'h7 == stage1_addr_line_mapping[10:4] ? way0_dirty_7 : _GEN_519; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_521 = 7'h8 == stage1_addr_line_mapping[10:4] ? way0_dirty_8 : _GEN_520; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_522 = 7'h9 == stage1_addr_line_mapping[10:4] ? way0_dirty_9 : _GEN_521; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_523 = 7'ha == stage1_addr_line_mapping[10:4] ? way0_dirty_10 : _GEN_522; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_524 = 7'hb == stage1_addr_line_mapping[10:4] ? way0_dirty_11 : _GEN_523; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_525 = 7'hc == stage1_addr_line_mapping[10:4] ? way0_dirty_12 : _GEN_524; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_526 = 7'hd == stage1_addr_line_mapping[10:4] ? way0_dirty_13 : _GEN_525; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_527 = 7'he == stage1_addr_line_mapping[10:4] ? way0_dirty_14 : _GEN_526; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_528 = 7'hf == stage1_addr_line_mapping[10:4] ? way0_dirty_15 : _GEN_527; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_529 = 7'h10 == stage1_addr_line_mapping[10:4] ? way0_dirty_16 : _GEN_528; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_530 = 7'h11 == stage1_addr_line_mapping[10:4] ? way0_dirty_17 : _GEN_529; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_531 = 7'h12 == stage1_addr_line_mapping[10:4] ? way0_dirty_18 : _GEN_530; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_532 = 7'h13 == stage1_addr_line_mapping[10:4] ? way0_dirty_19 : _GEN_531; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_533 = 7'h14 == stage1_addr_line_mapping[10:4] ? way0_dirty_20 : _GEN_532; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_534 = 7'h15 == stage1_addr_line_mapping[10:4] ? way0_dirty_21 : _GEN_533; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_535 = 7'h16 == stage1_addr_line_mapping[10:4] ? way0_dirty_22 : _GEN_534; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_536 = 7'h17 == stage1_addr_line_mapping[10:4] ? way0_dirty_23 : _GEN_535; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_537 = 7'h18 == stage1_addr_line_mapping[10:4] ? way0_dirty_24 : _GEN_536; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_538 = 7'h19 == stage1_addr_line_mapping[10:4] ? way0_dirty_25 : _GEN_537; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_539 = 7'h1a == stage1_addr_line_mapping[10:4] ? way0_dirty_26 : _GEN_538; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_540 = 7'h1b == stage1_addr_line_mapping[10:4] ? way0_dirty_27 : _GEN_539; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_541 = 7'h1c == stage1_addr_line_mapping[10:4] ? way0_dirty_28 : _GEN_540; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_542 = 7'h1d == stage1_addr_line_mapping[10:4] ? way0_dirty_29 : _GEN_541; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_543 = 7'h1e == stage1_addr_line_mapping[10:4] ? way0_dirty_30 : _GEN_542; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_544 = 7'h1f == stage1_addr_line_mapping[10:4] ? way0_dirty_31 : _GEN_543; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_545 = 7'h20 == stage1_addr_line_mapping[10:4] ? way0_dirty_32 : _GEN_544; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_546 = 7'h21 == stage1_addr_line_mapping[10:4] ? way0_dirty_33 : _GEN_545; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_547 = 7'h22 == stage1_addr_line_mapping[10:4] ? way0_dirty_34 : _GEN_546; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_548 = 7'h23 == stage1_addr_line_mapping[10:4] ? way0_dirty_35 : _GEN_547; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_549 = 7'h24 == stage1_addr_line_mapping[10:4] ? way0_dirty_36 : _GEN_548; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_550 = 7'h25 == stage1_addr_line_mapping[10:4] ? way0_dirty_37 : _GEN_549; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_551 = 7'h26 == stage1_addr_line_mapping[10:4] ? way0_dirty_38 : _GEN_550; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_552 = 7'h27 == stage1_addr_line_mapping[10:4] ? way0_dirty_39 : _GEN_551; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_553 = 7'h28 == stage1_addr_line_mapping[10:4] ? way0_dirty_40 : _GEN_552; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_554 = 7'h29 == stage1_addr_line_mapping[10:4] ? way0_dirty_41 : _GEN_553; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_555 = 7'h2a == stage1_addr_line_mapping[10:4] ? way0_dirty_42 : _GEN_554; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_556 = 7'h2b == stage1_addr_line_mapping[10:4] ? way0_dirty_43 : _GEN_555; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_557 = 7'h2c == stage1_addr_line_mapping[10:4] ? way0_dirty_44 : _GEN_556; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_558 = 7'h2d == stage1_addr_line_mapping[10:4] ? way0_dirty_45 : _GEN_557; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_559 = 7'h2e == stage1_addr_line_mapping[10:4] ? way0_dirty_46 : _GEN_558; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_560 = 7'h2f == stage1_addr_line_mapping[10:4] ? way0_dirty_47 : _GEN_559; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_561 = 7'h30 == stage1_addr_line_mapping[10:4] ? way0_dirty_48 : _GEN_560; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_562 = 7'h31 == stage1_addr_line_mapping[10:4] ? way0_dirty_49 : _GEN_561; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_563 = 7'h32 == stage1_addr_line_mapping[10:4] ? way0_dirty_50 : _GEN_562; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_564 = 7'h33 == stage1_addr_line_mapping[10:4] ? way0_dirty_51 : _GEN_563; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_565 = 7'h34 == stage1_addr_line_mapping[10:4] ? way0_dirty_52 : _GEN_564; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_566 = 7'h35 == stage1_addr_line_mapping[10:4] ? way0_dirty_53 : _GEN_565; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_567 = 7'h36 == stage1_addr_line_mapping[10:4] ? way0_dirty_54 : _GEN_566; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_568 = 7'h37 == stage1_addr_line_mapping[10:4] ? way0_dirty_55 : _GEN_567; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_569 = 7'h38 == stage1_addr_line_mapping[10:4] ? way0_dirty_56 : _GEN_568; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_570 = 7'h39 == stage1_addr_line_mapping[10:4] ? way0_dirty_57 : _GEN_569; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_571 = 7'h3a == stage1_addr_line_mapping[10:4] ? way0_dirty_58 : _GEN_570; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_572 = 7'h3b == stage1_addr_line_mapping[10:4] ? way0_dirty_59 : _GEN_571; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_573 = 7'h3c == stage1_addr_line_mapping[10:4] ? way0_dirty_60 : _GEN_572; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_574 = 7'h3d == stage1_addr_line_mapping[10:4] ? way0_dirty_61 : _GEN_573; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_575 = 7'h3e == stage1_addr_line_mapping[10:4] ? way0_dirty_62 : _GEN_574; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_576 = 7'h3f == stage1_addr_line_mapping[10:4] ? way0_dirty_63 : _GEN_575; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_577 = 7'h40 == stage1_addr_line_mapping[10:4] ? way0_dirty_64 : _GEN_576; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_578 = 7'h41 == stage1_addr_line_mapping[10:4] ? way0_dirty_65 : _GEN_577; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_579 = 7'h42 == stage1_addr_line_mapping[10:4] ? way0_dirty_66 : _GEN_578; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_580 = 7'h43 == stage1_addr_line_mapping[10:4] ? way0_dirty_67 : _GEN_579; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_581 = 7'h44 == stage1_addr_line_mapping[10:4] ? way0_dirty_68 : _GEN_580; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_582 = 7'h45 == stage1_addr_line_mapping[10:4] ? way0_dirty_69 : _GEN_581; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_583 = 7'h46 == stage1_addr_line_mapping[10:4] ? way0_dirty_70 : _GEN_582; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_584 = 7'h47 == stage1_addr_line_mapping[10:4] ? way0_dirty_71 : _GEN_583; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_585 = 7'h48 == stage1_addr_line_mapping[10:4] ? way0_dirty_72 : _GEN_584; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_586 = 7'h49 == stage1_addr_line_mapping[10:4] ? way0_dirty_73 : _GEN_585; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_587 = 7'h4a == stage1_addr_line_mapping[10:4] ? way0_dirty_74 : _GEN_586; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_588 = 7'h4b == stage1_addr_line_mapping[10:4] ? way0_dirty_75 : _GEN_587; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_589 = 7'h4c == stage1_addr_line_mapping[10:4] ? way0_dirty_76 : _GEN_588; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_590 = 7'h4d == stage1_addr_line_mapping[10:4] ? way0_dirty_77 : _GEN_589; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_591 = 7'h4e == stage1_addr_line_mapping[10:4] ? way0_dirty_78 : _GEN_590; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_592 = 7'h4f == stage1_addr_line_mapping[10:4] ? way0_dirty_79 : _GEN_591; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_593 = 7'h50 == stage1_addr_line_mapping[10:4] ? way0_dirty_80 : _GEN_592; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_594 = 7'h51 == stage1_addr_line_mapping[10:4] ? way0_dirty_81 : _GEN_593; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_595 = 7'h52 == stage1_addr_line_mapping[10:4] ? way0_dirty_82 : _GEN_594; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_596 = 7'h53 == stage1_addr_line_mapping[10:4] ? way0_dirty_83 : _GEN_595; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_597 = 7'h54 == stage1_addr_line_mapping[10:4] ? way0_dirty_84 : _GEN_596; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_598 = 7'h55 == stage1_addr_line_mapping[10:4] ? way0_dirty_85 : _GEN_597; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_599 = 7'h56 == stage1_addr_line_mapping[10:4] ? way0_dirty_86 : _GEN_598; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_600 = 7'h57 == stage1_addr_line_mapping[10:4] ? way0_dirty_87 : _GEN_599; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_601 = 7'h58 == stage1_addr_line_mapping[10:4] ? way0_dirty_88 : _GEN_600; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_602 = 7'h59 == stage1_addr_line_mapping[10:4] ? way0_dirty_89 : _GEN_601; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_603 = 7'h5a == stage1_addr_line_mapping[10:4] ? way0_dirty_90 : _GEN_602; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_604 = 7'h5b == stage1_addr_line_mapping[10:4] ? way0_dirty_91 : _GEN_603; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_605 = 7'h5c == stage1_addr_line_mapping[10:4] ? way0_dirty_92 : _GEN_604; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_606 = 7'h5d == stage1_addr_line_mapping[10:4] ? way0_dirty_93 : _GEN_605; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_607 = 7'h5e == stage1_addr_line_mapping[10:4] ? way0_dirty_94 : _GEN_606; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_608 = 7'h5f == stage1_addr_line_mapping[10:4] ? way0_dirty_95 : _GEN_607; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_609 = 7'h60 == stage1_addr_line_mapping[10:4] ? way0_dirty_96 : _GEN_608; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_610 = 7'h61 == stage1_addr_line_mapping[10:4] ? way0_dirty_97 : _GEN_609; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_611 = 7'h62 == stage1_addr_line_mapping[10:4] ? way0_dirty_98 : _GEN_610; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_612 = 7'h63 == stage1_addr_line_mapping[10:4] ? way0_dirty_99 : _GEN_611; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_613 = 7'h64 == stage1_addr_line_mapping[10:4] ? way0_dirty_100 : _GEN_612; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_614 = 7'h65 == stage1_addr_line_mapping[10:4] ? way0_dirty_101 : _GEN_613; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_615 = 7'h66 == stage1_addr_line_mapping[10:4] ? way0_dirty_102 : _GEN_614; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_616 = 7'h67 == stage1_addr_line_mapping[10:4] ? way0_dirty_103 : _GEN_615; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_617 = 7'h68 == stage1_addr_line_mapping[10:4] ? way0_dirty_104 : _GEN_616; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_618 = 7'h69 == stage1_addr_line_mapping[10:4] ? way0_dirty_105 : _GEN_617; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_619 = 7'h6a == stage1_addr_line_mapping[10:4] ? way0_dirty_106 : _GEN_618; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_620 = 7'h6b == stage1_addr_line_mapping[10:4] ? way0_dirty_107 : _GEN_619; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_621 = 7'h6c == stage1_addr_line_mapping[10:4] ? way0_dirty_108 : _GEN_620; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_622 = 7'h6d == stage1_addr_line_mapping[10:4] ? way0_dirty_109 : _GEN_621; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_623 = 7'h6e == stage1_addr_line_mapping[10:4] ? way0_dirty_110 : _GEN_622; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_624 = 7'h6f == stage1_addr_line_mapping[10:4] ? way0_dirty_111 : _GEN_623; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_625 = 7'h70 == stage1_addr_line_mapping[10:4] ? way0_dirty_112 : _GEN_624; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_626 = 7'h71 == stage1_addr_line_mapping[10:4] ? way0_dirty_113 : _GEN_625; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_627 = 7'h72 == stage1_addr_line_mapping[10:4] ? way0_dirty_114 : _GEN_626; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_628 = 7'h73 == stage1_addr_line_mapping[10:4] ? way0_dirty_115 : _GEN_627; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_629 = 7'h74 == stage1_addr_line_mapping[10:4] ? way0_dirty_116 : _GEN_628; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_630 = 7'h75 == stage1_addr_line_mapping[10:4] ? way0_dirty_117 : _GEN_629; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_631 = 7'h76 == stage1_addr_line_mapping[10:4] ? way0_dirty_118 : _GEN_630; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_632 = 7'h77 == stage1_addr_line_mapping[10:4] ? way0_dirty_119 : _GEN_631; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_633 = 7'h78 == stage1_addr_line_mapping[10:4] ? way0_dirty_120 : _GEN_632; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_634 = 7'h79 == stage1_addr_line_mapping[10:4] ? way0_dirty_121 : _GEN_633; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_635 = 7'h7a == stage1_addr_line_mapping[10:4] ? way0_dirty_122 : _GEN_634; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_636 = 7'h7b == stage1_addr_line_mapping[10:4] ? way0_dirty_123 : _GEN_635; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_637 = 7'h7c == stage1_addr_line_mapping[10:4] ? way0_dirty_124 : _GEN_636; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_638 = 7'h7d == stage1_addr_line_mapping[10:4] ? way0_dirty_125 : _GEN_637; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_639 = 7'h7e == stage1_addr_line_mapping[10:4] ? way0_dirty_126 : _GEN_638; // @[data_cache.scala 206:{12,12}]
  wire  _GEN_640 = 7'h7f == stage1_addr_line_mapping[10:4] ? way0_dirty_127 : _GEN_639; // @[data_cache.scala 206:{12,12}]
  wire  _way0_dirty_T_14 = work_state == 5'h10 & _way0_dirty_T_7 | _GEN_640; // @[data_cache.scala 206:12]
  wire  _way0_dirty_T_15 = work_state == 5'he & ~_GEN_384 ? 1'h0 : _way0_dirty_T_14; // @[data_cache.scala 205:12]
  wire  _way1_dirty_T_4 = _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 208:149]
  wire  _way1_dirty_T_12 = _way0_dirty_T_9 & _GEN_384; // @[data_cache.scala 210:52]
  wire  _GEN_1026 = 7'h1 == stage1_addr_line_mapping[10:4] ? way1_dirty_1 : way1_dirty_0; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1027 = 7'h2 == stage1_addr_line_mapping[10:4] ? way1_dirty_2 : _GEN_1026; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1028 = 7'h3 == stage1_addr_line_mapping[10:4] ? way1_dirty_3 : _GEN_1027; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1029 = 7'h4 == stage1_addr_line_mapping[10:4] ? way1_dirty_4 : _GEN_1028; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1030 = 7'h5 == stage1_addr_line_mapping[10:4] ? way1_dirty_5 : _GEN_1029; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1031 = 7'h6 == stage1_addr_line_mapping[10:4] ? way1_dirty_6 : _GEN_1030; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1032 = 7'h7 == stage1_addr_line_mapping[10:4] ? way1_dirty_7 : _GEN_1031; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1033 = 7'h8 == stage1_addr_line_mapping[10:4] ? way1_dirty_8 : _GEN_1032; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1034 = 7'h9 == stage1_addr_line_mapping[10:4] ? way1_dirty_9 : _GEN_1033; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1035 = 7'ha == stage1_addr_line_mapping[10:4] ? way1_dirty_10 : _GEN_1034; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1036 = 7'hb == stage1_addr_line_mapping[10:4] ? way1_dirty_11 : _GEN_1035; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1037 = 7'hc == stage1_addr_line_mapping[10:4] ? way1_dirty_12 : _GEN_1036; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1038 = 7'hd == stage1_addr_line_mapping[10:4] ? way1_dirty_13 : _GEN_1037; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1039 = 7'he == stage1_addr_line_mapping[10:4] ? way1_dirty_14 : _GEN_1038; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1040 = 7'hf == stage1_addr_line_mapping[10:4] ? way1_dirty_15 : _GEN_1039; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1041 = 7'h10 == stage1_addr_line_mapping[10:4] ? way1_dirty_16 : _GEN_1040; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1042 = 7'h11 == stage1_addr_line_mapping[10:4] ? way1_dirty_17 : _GEN_1041; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1043 = 7'h12 == stage1_addr_line_mapping[10:4] ? way1_dirty_18 : _GEN_1042; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1044 = 7'h13 == stage1_addr_line_mapping[10:4] ? way1_dirty_19 : _GEN_1043; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1045 = 7'h14 == stage1_addr_line_mapping[10:4] ? way1_dirty_20 : _GEN_1044; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1046 = 7'h15 == stage1_addr_line_mapping[10:4] ? way1_dirty_21 : _GEN_1045; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1047 = 7'h16 == stage1_addr_line_mapping[10:4] ? way1_dirty_22 : _GEN_1046; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1048 = 7'h17 == stage1_addr_line_mapping[10:4] ? way1_dirty_23 : _GEN_1047; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1049 = 7'h18 == stage1_addr_line_mapping[10:4] ? way1_dirty_24 : _GEN_1048; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1050 = 7'h19 == stage1_addr_line_mapping[10:4] ? way1_dirty_25 : _GEN_1049; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1051 = 7'h1a == stage1_addr_line_mapping[10:4] ? way1_dirty_26 : _GEN_1050; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1052 = 7'h1b == stage1_addr_line_mapping[10:4] ? way1_dirty_27 : _GEN_1051; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1053 = 7'h1c == stage1_addr_line_mapping[10:4] ? way1_dirty_28 : _GEN_1052; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1054 = 7'h1d == stage1_addr_line_mapping[10:4] ? way1_dirty_29 : _GEN_1053; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1055 = 7'h1e == stage1_addr_line_mapping[10:4] ? way1_dirty_30 : _GEN_1054; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1056 = 7'h1f == stage1_addr_line_mapping[10:4] ? way1_dirty_31 : _GEN_1055; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1057 = 7'h20 == stage1_addr_line_mapping[10:4] ? way1_dirty_32 : _GEN_1056; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1058 = 7'h21 == stage1_addr_line_mapping[10:4] ? way1_dirty_33 : _GEN_1057; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1059 = 7'h22 == stage1_addr_line_mapping[10:4] ? way1_dirty_34 : _GEN_1058; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1060 = 7'h23 == stage1_addr_line_mapping[10:4] ? way1_dirty_35 : _GEN_1059; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1061 = 7'h24 == stage1_addr_line_mapping[10:4] ? way1_dirty_36 : _GEN_1060; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1062 = 7'h25 == stage1_addr_line_mapping[10:4] ? way1_dirty_37 : _GEN_1061; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1063 = 7'h26 == stage1_addr_line_mapping[10:4] ? way1_dirty_38 : _GEN_1062; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1064 = 7'h27 == stage1_addr_line_mapping[10:4] ? way1_dirty_39 : _GEN_1063; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1065 = 7'h28 == stage1_addr_line_mapping[10:4] ? way1_dirty_40 : _GEN_1064; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1066 = 7'h29 == stage1_addr_line_mapping[10:4] ? way1_dirty_41 : _GEN_1065; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1067 = 7'h2a == stage1_addr_line_mapping[10:4] ? way1_dirty_42 : _GEN_1066; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1068 = 7'h2b == stage1_addr_line_mapping[10:4] ? way1_dirty_43 : _GEN_1067; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1069 = 7'h2c == stage1_addr_line_mapping[10:4] ? way1_dirty_44 : _GEN_1068; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1070 = 7'h2d == stage1_addr_line_mapping[10:4] ? way1_dirty_45 : _GEN_1069; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1071 = 7'h2e == stage1_addr_line_mapping[10:4] ? way1_dirty_46 : _GEN_1070; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1072 = 7'h2f == stage1_addr_line_mapping[10:4] ? way1_dirty_47 : _GEN_1071; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1073 = 7'h30 == stage1_addr_line_mapping[10:4] ? way1_dirty_48 : _GEN_1072; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1074 = 7'h31 == stage1_addr_line_mapping[10:4] ? way1_dirty_49 : _GEN_1073; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1075 = 7'h32 == stage1_addr_line_mapping[10:4] ? way1_dirty_50 : _GEN_1074; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1076 = 7'h33 == stage1_addr_line_mapping[10:4] ? way1_dirty_51 : _GEN_1075; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1077 = 7'h34 == stage1_addr_line_mapping[10:4] ? way1_dirty_52 : _GEN_1076; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1078 = 7'h35 == stage1_addr_line_mapping[10:4] ? way1_dirty_53 : _GEN_1077; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1079 = 7'h36 == stage1_addr_line_mapping[10:4] ? way1_dirty_54 : _GEN_1078; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1080 = 7'h37 == stage1_addr_line_mapping[10:4] ? way1_dirty_55 : _GEN_1079; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1081 = 7'h38 == stage1_addr_line_mapping[10:4] ? way1_dirty_56 : _GEN_1080; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1082 = 7'h39 == stage1_addr_line_mapping[10:4] ? way1_dirty_57 : _GEN_1081; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1083 = 7'h3a == stage1_addr_line_mapping[10:4] ? way1_dirty_58 : _GEN_1082; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1084 = 7'h3b == stage1_addr_line_mapping[10:4] ? way1_dirty_59 : _GEN_1083; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1085 = 7'h3c == stage1_addr_line_mapping[10:4] ? way1_dirty_60 : _GEN_1084; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1086 = 7'h3d == stage1_addr_line_mapping[10:4] ? way1_dirty_61 : _GEN_1085; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1087 = 7'h3e == stage1_addr_line_mapping[10:4] ? way1_dirty_62 : _GEN_1086; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1088 = 7'h3f == stage1_addr_line_mapping[10:4] ? way1_dirty_63 : _GEN_1087; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1089 = 7'h40 == stage1_addr_line_mapping[10:4] ? way1_dirty_64 : _GEN_1088; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1090 = 7'h41 == stage1_addr_line_mapping[10:4] ? way1_dirty_65 : _GEN_1089; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1091 = 7'h42 == stage1_addr_line_mapping[10:4] ? way1_dirty_66 : _GEN_1090; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1092 = 7'h43 == stage1_addr_line_mapping[10:4] ? way1_dirty_67 : _GEN_1091; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1093 = 7'h44 == stage1_addr_line_mapping[10:4] ? way1_dirty_68 : _GEN_1092; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1094 = 7'h45 == stage1_addr_line_mapping[10:4] ? way1_dirty_69 : _GEN_1093; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1095 = 7'h46 == stage1_addr_line_mapping[10:4] ? way1_dirty_70 : _GEN_1094; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1096 = 7'h47 == stage1_addr_line_mapping[10:4] ? way1_dirty_71 : _GEN_1095; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1097 = 7'h48 == stage1_addr_line_mapping[10:4] ? way1_dirty_72 : _GEN_1096; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1098 = 7'h49 == stage1_addr_line_mapping[10:4] ? way1_dirty_73 : _GEN_1097; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1099 = 7'h4a == stage1_addr_line_mapping[10:4] ? way1_dirty_74 : _GEN_1098; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1100 = 7'h4b == stage1_addr_line_mapping[10:4] ? way1_dirty_75 : _GEN_1099; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1101 = 7'h4c == stage1_addr_line_mapping[10:4] ? way1_dirty_76 : _GEN_1100; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1102 = 7'h4d == stage1_addr_line_mapping[10:4] ? way1_dirty_77 : _GEN_1101; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1103 = 7'h4e == stage1_addr_line_mapping[10:4] ? way1_dirty_78 : _GEN_1102; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1104 = 7'h4f == stage1_addr_line_mapping[10:4] ? way1_dirty_79 : _GEN_1103; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1105 = 7'h50 == stage1_addr_line_mapping[10:4] ? way1_dirty_80 : _GEN_1104; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1106 = 7'h51 == stage1_addr_line_mapping[10:4] ? way1_dirty_81 : _GEN_1105; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1107 = 7'h52 == stage1_addr_line_mapping[10:4] ? way1_dirty_82 : _GEN_1106; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1108 = 7'h53 == stage1_addr_line_mapping[10:4] ? way1_dirty_83 : _GEN_1107; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1109 = 7'h54 == stage1_addr_line_mapping[10:4] ? way1_dirty_84 : _GEN_1108; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1110 = 7'h55 == stage1_addr_line_mapping[10:4] ? way1_dirty_85 : _GEN_1109; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1111 = 7'h56 == stage1_addr_line_mapping[10:4] ? way1_dirty_86 : _GEN_1110; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1112 = 7'h57 == stage1_addr_line_mapping[10:4] ? way1_dirty_87 : _GEN_1111; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1113 = 7'h58 == stage1_addr_line_mapping[10:4] ? way1_dirty_88 : _GEN_1112; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1114 = 7'h59 == stage1_addr_line_mapping[10:4] ? way1_dirty_89 : _GEN_1113; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1115 = 7'h5a == stage1_addr_line_mapping[10:4] ? way1_dirty_90 : _GEN_1114; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1116 = 7'h5b == stage1_addr_line_mapping[10:4] ? way1_dirty_91 : _GEN_1115; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1117 = 7'h5c == stage1_addr_line_mapping[10:4] ? way1_dirty_92 : _GEN_1116; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1118 = 7'h5d == stage1_addr_line_mapping[10:4] ? way1_dirty_93 : _GEN_1117; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1119 = 7'h5e == stage1_addr_line_mapping[10:4] ? way1_dirty_94 : _GEN_1118; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1120 = 7'h5f == stage1_addr_line_mapping[10:4] ? way1_dirty_95 : _GEN_1119; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1121 = 7'h60 == stage1_addr_line_mapping[10:4] ? way1_dirty_96 : _GEN_1120; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1122 = 7'h61 == stage1_addr_line_mapping[10:4] ? way1_dirty_97 : _GEN_1121; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1123 = 7'h62 == stage1_addr_line_mapping[10:4] ? way1_dirty_98 : _GEN_1122; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1124 = 7'h63 == stage1_addr_line_mapping[10:4] ? way1_dirty_99 : _GEN_1123; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1125 = 7'h64 == stage1_addr_line_mapping[10:4] ? way1_dirty_100 : _GEN_1124; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1126 = 7'h65 == stage1_addr_line_mapping[10:4] ? way1_dirty_101 : _GEN_1125; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1127 = 7'h66 == stage1_addr_line_mapping[10:4] ? way1_dirty_102 : _GEN_1126; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1128 = 7'h67 == stage1_addr_line_mapping[10:4] ? way1_dirty_103 : _GEN_1127; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1129 = 7'h68 == stage1_addr_line_mapping[10:4] ? way1_dirty_104 : _GEN_1128; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1130 = 7'h69 == stage1_addr_line_mapping[10:4] ? way1_dirty_105 : _GEN_1129; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1131 = 7'h6a == stage1_addr_line_mapping[10:4] ? way1_dirty_106 : _GEN_1130; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1132 = 7'h6b == stage1_addr_line_mapping[10:4] ? way1_dirty_107 : _GEN_1131; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1133 = 7'h6c == stage1_addr_line_mapping[10:4] ? way1_dirty_108 : _GEN_1132; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1134 = 7'h6d == stage1_addr_line_mapping[10:4] ? way1_dirty_109 : _GEN_1133; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1135 = 7'h6e == stage1_addr_line_mapping[10:4] ? way1_dirty_110 : _GEN_1134; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1136 = 7'h6f == stage1_addr_line_mapping[10:4] ? way1_dirty_111 : _GEN_1135; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1137 = 7'h70 == stage1_addr_line_mapping[10:4] ? way1_dirty_112 : _GEN_1136; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1138 = 7'h71 == stage1_addr_line_mapping[10:4] ? way1_dirty_113 : _GEN_1137; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1139 = 7'h72 == stage1_addr_line_mapping[10:4] ? way1_dirty_114 : _GEN_1138; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1140 = 7'h73 == stage1_addr_line_mapping[10:4] ? way1_dirty_115 : _GEN_1139; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1141 = 7'h74 == stage1_addr_line_mapping[10:4] ? way1_dirty_116 : _GEN_1140; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1142 = 7'h75 == stage1_addr_line_mapping[10:4] ? way1_dirty_117 : _GEN_1141; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1143 = 7'h76 == stage1_addr_line_mapping[10:4] ? way1_dirty_118 : _GEN_1142; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1144 = 7'h77 == stage1_addr_line_mapping[10:4] ? way1_dirty_119 : _GEN_1143; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1145 = 7'h78 == stage1_addr_line_mapping[10:4] ? way1_dirty_120 : _GEN_1144; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1146 = 7'h79 == stage1_addr_line_mapping[10:4] ? way1_dirty_121 : _GEN_1145; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1147 = 7'h7a == stage1_addr_line_mapping[10:4] ? way1_dirty_122 : _GEN_1146; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1148 = 7'h7b == stage1_addr_line_mapping[10:4] ? way1_dirty_123 : _GEN_1147; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1149 = 7'h7c == stage1_addr_line_mapping[10:4] ? way1_dirty_124 : _GEN_1148; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1150 = 7'h7d == stage1_addr_line_mapping[10:4] ? way1_dirty_125 : _GEN_1149; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1151 = 7'h7e == stage1_addr_line_mapping[10:4] ? way1_dirty_126 : _GEN_1150; // @[data_cache.scala 210:{12,12}]
  wire  _GEN_1152 = 7'h7f == stage1_addr_line_mapping[10:4] ? way1_dirty_127 : _GEN_1151; // @[data_cache.scala 210:{12,12}]
  wire  _way1_dirty_T_14 = _way0_dirty_T_9 & _GEN_384 | _GEN_1152; // @[data_cache.scala 210:12]
  wire  _way1_dirty_T_15 = _way0_dirty_T_5 & _GEN_384 ? 1'h0 : _way1_dirty_T_14; // @[data_cache.scala 209:12]
  wire  dirty_victim = _way0_dirty_T_7 ? _GEN_640 : _GEN_1152; // @[data_cache.scala 214:24]
  wire [10:0] _T_3 = {data_write_back_counter[6:0],4'h0}; // @[Cat.scala 31:58]
  wire  _tlb_req_T_4 = ~stage1_addr_line_mapping[31] | stage1_addr_line_mapping[31:30] == 2'h3; // @[macros.scala 492:18]
  wire  tlb_req = _tlb_req_T_4 & stage1_sram_req_reg; // @[data_cache.scala 226:51]
  wire  _lru_T_4 = _hit_T_1 ? 1'h0 : _GEN_384; // @[data_cache.scala 235:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[data_cache.scala 234:12]
  wire  _data_cache_under_write_all_back_T = work_state == 5'h18; // @[data_cache.scala 242:55]
  wire  _data_cache_under_write_all_back_T_1 = work_state == 5'h19; // @[data_cache.scala 242:90]
  wire [4:0] _state_ready_lookup_will_to_be_T_3 = stage1_sram_cache_reg ? 5'h19 : 5'h3; // @[data_cache.scala 245:16]
  wire [4:0] _state_ready_lookup_will_to_be_T_5 = stage1_sram_cache_reg ? 5'h19 : 5'h1; // @[data_cache.scala 245:88]
  wire [4:0] _state_ready_lookup_will_to_be_T_6 = stage1_sram_wr_reg ? _state_ready_lookup_will_to_be_T_3 :
    _state_ready_lookup_will_to_be_T_5; // @[data_cache.scala 244:55]
  wire [4:0] _state_ready_lookup_will_to_be_T_7 = stage1_sram_req_reg ? _state_ready_lookup_will_to_be_T_6 : 5'h19; // @[data_cache.scala 244:24]
  wire [1:0] _state_ready_lookup_will_to_be_T_12 = stage1_sram_wr_reg ? 2'h3 : 2'h1; // @[data_cache.scala 246:81]
  wire [3:0] _state_ready_lookup_will_to_be_T_15 = stage1_sram_wr_reg ? 4'h8 : 4'hc; // @[data_cache.scala 247:64]
  wire [3:0] _state_ready_lookup_will_to_be_T_16 = dirty_victim ? 4'h9 : _state_ready_lookup_will_to_be_T_15; // @[data_cache.scala 247:16]
  wire [3:0] _state_ready_lookup_will_to_be_T_17 = ~stage1_sram_cache_reg ? {{2'd0}, _state_ready_lookup_will_to_be_T_12
    } : _state_ready_lookup_will_to_be_T_16; // @[data_cache.scala 246:47]
  wire [4:0] _state_ready_lookup_will_to_be_T_18 = stage1_sram_req_reg ? {{1'd0}, _state_ready_lookup_will_to_be_T_17}
     : 5'h19; // @[data_cache.scala 246:16]
  wire [4:0] _state_ready_lookup_will_to_be_T_19 = hit ? _state_ready_lookup_will_to_be_T_7 :
    _state_ready_lookup_will_to_be_T_18; // @[data_cache.scala 244:16]
  wire [4:0] state_ready_lookup_will_to_be = io_fence_i_control ? 5'h11 : _state_ready_lookup_will_to_be_T_19; // @[data_cache.scala 243:41]
  wire [4:0] _access_work_state_T_1 = io_port_arready ? 5'h2 : work_state; // @[data_cache.scala 254:39]
  wire [4:0] _access_work_state_T_3 = io_port_rvalid ? 5'h18 : work_state; // @[data_cache.scala 255:39]
  wire [2:0] _access_work_state_T_6 = io_port_wready ? 3'h5 : 3'h4; // @[data_cache.scala 257:66]
  wire [4:0] _access_work_state_T_7 = io_port_awready ? {{2'd0}, _access_work_state_T_6} : work_state; // @[data_cache.scala 257:39]
  wire [4:0] _access_work_state_T_9 = io_port_wready ? 5'h5 : work_state; // @[data_cache.scala 258:39]
  wire [4:0] _access_work_state_T_11 = io_port_bvalid ? 5'h18 : 5'h5; // @[data_cache.scala 259:39]
  wire [4:0] _access_work_state_T_13 = io_port_arready ? 5'hd : work_state; // @[data_cache.scala 262:44]
  wire [4:0] _access_work_state_T_18 = stage1_sram_wr_reg ? 5'h10 : 5'he; // @[data_cache.scala 263:94]
  wire [4:0] _access_work_state_T_19 = io_port_rlast & io_port_rvalid ? _access_work_state_T_18 : work_state; // @[data_cache.scala 263:44]
  wire [4:0] _access_work_state_T_21 = io_port_awready ? 5'ha : work_state; // @[data_cache.scala 265:41]
  wire  _access_work_state_T_23 = write_counter == 3'h1; // @[data_cache.scala 266:81]
  wire  _access_work_state_T_24 = io_port_wready & write_counter == 3'h1; // @[data_cache.scala 266:64]
  wire [4:0] _access_work_state_T_25 = io_port_wready & write_counter == 3'h1 ? 5'hb : work_state; // @[data_cache.scala 266:41]
  wire [4:0] _access_work_state_T_27 = io_port_bvalid ? 5'hc : work_state; // @[data_cache.scala 267:41]
  wire [4:0] _access_work_state_T_29 = io_port_arready ? 5'h0 : work_state; // @[data_cache.scala 269:44]
  wire  _access_work_state_T_32 = io_port_rvalid & io_port_rlast; // @[data_cache.scala 270:68]
  wire [4:0] _access_work_state_T_33 = io_port_rvalid & io_port_rlast ? 5'h10 : work_state; // @[data_cache.scala 270:44]
  wire [4:0] _access_work_state_T_35 = io_port_awready ? 5'h6 : work_state; // @[data_cache.scala 272:41]
  wire [4:0] _access_work_state_T_39 = _access_work_state_T_24 ? 5'h7 : work_state; // @[data_cache.scala 273:41]
  wire [4:0] _access_work_state_T_41 = io_port_bvalid ? 5'h8 : work_state; // @[data_cache.scala 274:41]
  wire [4:0] _access_work_state_T_42 = data_all_write_back ? 5'h18 : work_state; // @[data_cache.scala 277:95]
  wire [4:0] _access_work_state_T_43 = data_should_write_back ? 5'h12 : _access_work_state_T_42; // @[data_cache.scala 277:42]
  wire [4:0] _access_work_state_T_45 = io_port_awready ? 5'h13 : work_state; // @[data_cache.scala 278:41]
  wire [4:0] _access_work_state_T_49 = _access_work_state_T_24 ? 5'h14 : work_state; // @[data_cache.scala 279:41]
  wire [4:0] _access_work_state_T_54 = 5'h1 == work_state ? _access_work_state_T_1 : work_state; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_56 = 5'h2 == work_state ? _access_work_state_T_3 : _access_work_state_T_54; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_58 = 5'h18 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_56; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_60 = 5'h3 == work_state ? _access_work_state_T_7 : _access_work_state_T_58; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_62 = 5'h4 == work_state ? _access_work_state_T_9 : _access_work_state_T_60; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_64 = 5'h5 == work_state ? _access_work_state_T_11 : _access_work_state_T_62; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_66 = 5'h19 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_64; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_68 = 5'hc == work_state ? _access_work_state_T_13 : _access_work_state_T_66; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_70 = 5'hd == work_state ? _access_work_state_T_19 : _access_work_state_T_68; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_72 = 5'he == work_state ? 5'h18 : _access_work_state_T_70; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_74 = 5'h9 == work_state ? _access_work_state_T_21 : _access_work_state_T_72; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_76 = 5'ha == work_state ? _access_work_state_T_25 : _access_work_state_T_74; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_78 = 5'hb == work_state ? _access_work_state_T_27 : _access_work_state_T_76; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_80 = 5'h8 == work_state ? _access_work_state_T_29 : _access_work_state_T_78; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_82 = 5'h0 == work_state ? _access_work_state_T_33 : _access_work_state_T_80; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_84 = 5'h10 == work_state ? 5'h18 : _access_work_state_T_82; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_86 = 5'hf == work_state ? _access_work_state_T_35 : _access_work_state_T_84; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_88 = 5'h6 == work_state ? _access_work_state_T_39 : _access_work_state_T_86; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_90 = 5'h7 == work_state ? _access_work_state_T_41 : _access_work_state_T_88; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_92 = 5'h11 == work_state ? _access_work_state_T_43 : _access_work_state_T_90; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_94 = 5'h12 == work_state ? _access_work_state_T_45 : _access_work_state_T_92; // @[Mux.scala 81:58]
  wire  _wait_data_T_3 = work_state == 5'hd; // @[data_cache.scala 300:24]
  wire [2:0] _GEN_3468 = {{2'd0}, stage1_addr_line_mapping[3]}; // @[data_cache.scala 300:98]
  wire  _write_counter_T = work_state == 5'ha; // @[data_cache.scala 302:37]
  wire  _write_counter_T_1 = work_state == 5'h9; // @[data_cache.scala 302:79]
  wire  _write_counter_T_2 = work_state == 5'ha | work_state == 5'h9; // @[data_cache.scala 302:65]
  wire [2:0] _write_counter_T_6 = write_counter + 3'h1; // @[data_cache.scala 302:190]
  wire [2:0] _write_counter_T_7 = _access_work_state_T_23 ? 3'h0 : _write_counter_T_6; // @[data_cache.scala 302:137]
  wire [2:0] _write_counter_T_8 = io_port_wready ? _write_counter_T_7 : write_counter; // @[data_cache.scala 302:111]
  wire  _write_counter_T_9 = work_state == 5'h6; // @[data_cache.scala 303:24]
  wire  _write_counter_T_10 = work_state == 5'hf; // @[data_cache.scala 303:67]
  wire [2:0] _read_counter_T_6 = read_counter + 3'h1; // @[data_cache.scala 305:163]
  wire [2:0] _read_counter_T_7 = io_port_rvalid ? _read_counter_T_6 : read_counter; // @[data_cache.scala 305:128]
  wire [2:0] _read_counter_T_8 = _access_work_state_T_32 ? 3'h0 : _read_counter_T_7; // @[data_cache.scala 305:72]
  wire  _read_counter_T_9 = work_state == 5'h0; // @[data_cache.scala 306:24]
  reg [31:0] stage2_sram_addr_reg; // @[Reg.scala 28:20]
  reg  stage2_hit0_reg; // @[data_cache.scala 328:34]
  wire [63:0] dcache_data_way0_0_rdata = dcache_data_io_rdata; // @[data_cache.scala 95:{36,36}]
  wire [63:0] dcache_data_way0_1_rdata = dcache_data_1_io_rdata; // @[data_cache.scala 95:{36,36}]
  wire [63:0] _GEN_2179 = stage2_sram_addr_reg[3] ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 353:{23,23}]
  wire [63:0] dcache_data_way1_0_rdata = dcache_data_2_io_rdata; // @[data_cache.scala 96:{36,36}]
  wire [63:0] dcache_data_way1_1_rdata = dcache_data_3_io_rdata; // @[data_cache.scala 96:{36,36}]
  wire [63:0] _GEN_2181 = stage2_sram_addr_reg[3] ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 353:{23,23}]
  wire [63:0] hit_word = stage2_hit0_reg ? _GEN_2179 : _GEN_2181; // @[data_cache.scala 353:23]
  wire [63:0] _GEN_2183 = write_counter[0] ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 363:{29,29}]
  wire [63:0] _GEN_2185 = write_counter[0] ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 363:{29,29}]
  wire  data_write_back_way = data_cache_under_write_back ? data_write_back_counter[7] : _GEN_384; // @[data_cache.scala 364:31]
  wire [63:0] writeback_data = data_write_back_way ? _GEN_2183 : _GEN_2185; // @[data_cache.scala 363:29]
  wire  _way0_burst_read_wen_T_2 = _wait_data_T_3 | _read_counter_T_9; // @[data_cache.scala 366:76]
  wire  _way0_burst_read_wen_T_4 = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid; // @[data_cache.scala 366:124]
  wire  way0_burst_read_wen = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid & _way0_dirty_T_7; // @[data_cache.scala 366:149]
  wire  way1_burst_read_wen = _way0_burst_read_wen_T_4 & _GEN_384; // @[data_cache.scala 367:149]
  wire  _dcache_data_way0_0_wdata_T_2 = _way0_dirty_T_9 | _way0_dirty_T; // @[data_cache.scala 370:81]
  wire [63:0] _dcache_data_way0_0_wdata_T_6 = _way0_burst_read_wen_T_2 ? io_port_rdata : 64'h0; // @[data_cache.scala 370:155]
  wire  _wen_way0_wire_0_T_1 = ~stage1_addr_line_mapping[3]; // @[data_cache.scala 380:59]
  wire  _way0_wen_0_T = 3'h0 == read_counter; // @[data_cache.scala 386:38]
  wire  way0_wen_0 = 3'h0 == read_counter & way0_burst_read_wen; // @[data_cache.scala 386:28]
  wire [7:0] _wen_way0_wire_0_T_13 = {way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,
    way0_wen_0}; // @[Cat.scala 31:58]
  wire  way1_wen_0 = _way0_wen_0_T & way1_burst_read_wen; // @[data_cache.scala 387:28]
  wire [7:0] _wen_way1_wire_0_T_13 = {way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,
    way1_wen_0}; // @[Cat.scala 31:58]
  wire  _way0_wen_1_T = 3'h1 == read_counter; // @[data_cache.scala 386:38]
  wire  way0_wen_1 = 3'h1 == read_counter & way0_burst_read_wen; // @[data_cache.scala 386:28]
  wire [7:0] _wen_way0_wire_1_T_13 = {way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,
    way0_wen_1}; // @[Cat.scala 31:58]
  wire  way1_wen_1 = _way0_wen_1_T & way1_burst_read_wen; // @[data_cache.scala 387:28]
  wire [7:0] _wen_way1_wire_1_T_13 = {way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,
    way1_wen_1}; // @[Cat.scala 31:58]
  wire [21:0] _T_27 = {1'h1,stage1_addr_line_mapping[31:11]}; // @[Cat.scala 31:58]
  wire  _io_port_araddr_T = work_state == 5'h1; // @[data_cache.scala 406:38]
  wire  _io_port_araddr_T_1 = work_state == 5'hc; // @[data_cache.scala 407:24]
  wire  _io_port_araddr_T_2 = work_state == 5'h8; // @[data_cache.scala 407:71]
  wire [31:0] _io_port_araddr_T_5 = {stage1_sram_phy_addr_reg[31:4],4'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_port_araddr_T_6 = work_state == 5'hc | work_state == 5'h8 ? _io_port_araddr_T_5 : 32'h0; // @[data_cache.scala 407:12]
  wire  stage2_addr_same_as_stage1 = stage2_sram_addr_reg == stage1_addr_line_mapping; // @[data_cache.scala 418:56]
  wire  stage2_write_stage1_read = stage2_sram_write_reg & ~stage1_sram_wr_reg; // @[data_cache.scala 419:58]
  wire  _T_35 = work_state == 5'h3; // @[data_cache.scala 420:21]
  wire  _GEN_3338 = io_port_bvalid ? 1'h0 : write_access_complete_reg; // @[data_cache.scala 422:39 423:35 425:35]
  wire  _GEN_3339 = work_state == 5'h3 | _GEN_3338; // @[data_cache.scala 420:52 421:35]
  wire [20:0] _awaddr_miss_addr_T_2 = _way0_dirty_T_7 ? dcache_tag_io_tag : dcache_tag_1_io_tag; // @[data_cache.scala 428:36]
  wire [31:0] awaddr_miss_addr = {_awaddr_miss_addr_T_2,stage1_sram_phy_addr_reg[10:4],4'h0}; // @[Cat.scala 31:58]
  wire  _io_port_arvalid_T_7 = ~(stage2_addr_same_as_stage1 & stage2_write_stage1_read & write_access_complete_reg); // @[data_cache.scala 431:53]
  wire [20:0] _io_port_awaddr_T_1 = data_write_back_way ? dcache_tag_1_io_tag : dcache_tag_io_tag; // @[data_cache.scala 439:46]
  wire [31:0] _io_port_awaddr_T_3 = {_io_port_awaddr_T_1,data_write_back_counter[6:0],4'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_port_awaddr_T_5 = 5'h3 == work_state ? stage1_sram_phy_addr_reg : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_port_awaddr_T_7 = 5'h9 == work_state ? awaddr_miss_addr : _io_port_awaddr_T_5; // @[Mux.scala 81:58]
  wire [31:0] _io_port_awaddr_T_9 = 5'hf == work_state ? awaddr_miss_addr : _io_port_awaddr_T_7; // @[Mux.scala 81:58]
  wire  _io_port_awlen_T_2 = stage1_sram_cache_reg | _data_cache_under_write_back_T_3; // @[data_cache.scala 440:57]
  wire  _io_port_awvalid_T_4 = _T_35 | _write_counter_T_10 | _write_counter_T_1; // @[data_cache.scala 449:110]
  wire [63:0] _axi_line_wdata_T_2 = {stage1_sram_wdata_reg[55:0],8'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_4 = {stage1_sram_wdata_reg[47:0],16'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_6 = {stage1_sram_wdata_reg[39:0],24'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_8 = {stage1_sram_wdata_reg[31:0],32'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_10 = {stage1_sram_wdata_reg[23:0],40'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_12 = {stage1_sram_wdata_reg[15:0],48'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_14 = {stage1_sram_wdata_reg[7:0],56'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_line_wdata_T_16 = 3'h1 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_2 : stage1_sram_wdata_reg
    ; // @[Mux.scala 81:58]
  wire [63:0] _axi_line_wdata_T_18 = 3'h2 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_4 : _axi_line_wdata_T_16; // @[Mux.scala 81:58]
  wire [63:0] _axi_line_wdata_T_20 = 3'h3 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_6 : _axi_line_wdata_T_18; // @[Mux.scala 81:58]
  wire [63:0] _axi_line_wdata_T_22 = 3'h4 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_8 : _axi_line_wdata_T_20; // @[Mux.scala 81:58]
  wire [63:0] _axi_line_wdata_T_24 = 3'h5 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_10 : _axi_line_wdata_T_22
    ; // @[Mux.scala 81:58]
  wire [63:0] _axi_line_wdata_T_26 = 3'h6 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_12 : _axi_line_wdata_T_24
    ; // @[Mux.scala 81:58]
  wire [63:0] axi_line_wdata = 3'h7 == stage1_sram_phy_addr_reg[2:0] ? _axi_line_wdata_T_14 : _axi_line_wdata_T_26; // @[Mux.scala 81:58]
  wire  _io_port_wdata_T = work_state == 5'h4; // @[data_cache.scala 464:38]
  wire  _io_port_wdata_T_2 = work_state == 5'h4 | _T_35; // @[data_cache.scala 464:67]
  wire  _io_port_wdata_T_7 = _write_counter_T_2 | _write_counter_T_10; // @[data_cache.scala 465:109]
  wire  _io_port_wdata_T_11 = _io_port_wdata_T_7 | _write_counter_T_9 | _data_cache_under_write_back_T_3; // @[data_cache.scala 466:92]
  wire  _io_port_wdata_T_13 = _io_port_wdata_T_11 | _data_cache_under_write_back_T_5; // @[data_cache.scala 467:48]
  wire [63:0] _io_port_wdata_T_14 = _io_port_wdata_T_13 ? writeback_data : 64'h0; // @[data_cache.scala 465:27]
  wire [7:0] _io_port_wstrb_T_14 = _io_port_wdata_T_13 ? 8'hff : 8'h0; // @[data_cache.scala 468:131]
  wire  _io_port_wlast_T_7 = _write_counter_T | _write_counter_T_9; // @[data_cache.scala 471:176]
  wire  _io_port_wlast_T_11 = _io_port_wlast_T_7 | _data_cache_under_write_back_T_3 | _data_cache_under_write_back_T_5; // @[data_cache.scala 472:53]
  wire  _io_port_wlast_T_13 = _io_port_wlast_T_11 & _access_work_state_T_23; // @[data_cache.scala 473:9]
  wire  _io_port_wvalid_T_8 = _io_port_wdata_T_2 | _write_counter_T | _write_counter_T_1 | _write_counter_T_10; // @[data_cache.scala 474:190]
  reg [63:0] sram_rdata_reg; // @[data_cache.scala 481:33]
  reg  stage2_stall_reg; // @[data_cache.scala 483:35]
  wire [63:0] _io_sram_rdata_T_2 = _data_cache_under_write_all_back_T_1 ? hit_word : 64'h0; // @[data_cache.scala 485:92]
  wire [63:0] _io_sram_rdata_T_3 = _data_cache_under_write_all_back_T ? wait_data : _io_sram_rdata_T_2; // @[data_cache.scala 485:46]
  ysyx_22040886_dcache_tag dcache_tag ( // @[data_cache.scala 62:30]
    .clock(dcache_tag_clock),
    .reset(dcache_tag_reset),
    .io_wen(dcache_tag_io_wen),
    .io_wdata(dcache_tag_io_wdata),
    .io_raddr(dcache_tag_io_raddr),
    .io_waddr(dcache_tag_io_waddr),
    .io_hit(dcache_tag_io_hit),
    .io_valid(dcache_tag_io_valid),
    .io_tag(dcache_tag_io_tag),
    .io_w_valid(dcache_tag_io_w_valid)
  );
  ysyx_22040886_dcache_tag dcache_tag_1 ( // @[data_cache.scala 63:30]
    .clock(dcache_tag_1_clock),
    .reset(dcache_tag_1_reset),
    .io_wen(dcache_tag_1_io_wen),
    .io_wdata(dcache_tag_1_io_wdata),
    .io_raddr(dcache_tag_1_io_raddr),
    .io_waddr(dcache_tag_1_io_waddr),
    .io_hit(dcache_tag_1_io_hit),
    .io_valid(dcache_tag_1_io_valid),
    .io_tag(dcache_tag_1_io_tag),
    .io_w_valid(dcache_tag_1_io_w_valid)
  );
  ysyx_22040886_dcache_data dcache_data ( // @[data_cache.scala 95:62]
    .clock(dcache_data_clock),
    .io_wen(dcache_data_io_wen),
    .io_addr(dcache_data_io_addr),
    .io_wdata(dcache_data_io_wdata),
    .io_rdata(dcache_data_io_rdata),
    .io_sram_addr(dcache_data_io_sram_addr),
    .io_sram_wen(dcache_data_io_sram_wen),
    .io_sram_wmask(dcache_data_io_sram_wmask),
    .io_sram_wdata(dcache_data_io_sram_wdata),
    .io_sram_rdata(dcache_data_io_sram_rdata)
  );
  ysyx_22040886_dcache_data dcache_data_1 ( // @[data_cache.scala 95:62]
    .clock(dcache_data_1_clock),
    .io_wen(dcache_data_1_io_wen),
    .io_addr(dcache_data_1_io_addr),
    .io_wdata(dcache_data_1_io_wdata),
    .io_rdata(dcache_data_1_io_rdata),
    .io_sram_addr(dcache_data_1_io_sram_addr),
    .io_sram_wen(dcache_data_1_io_sram_wen),
    .io_sram_wmask(dcache_data_1_io_sram_wmask),
    .io_sram_wdata(dcache_data_1_io_sram_wdata),
    .io_sram_rdata(dcache_data_1_io_sram_rdata)
  );
  ysyx_22040886_dcache_data dcache_data_2 ( // @[data_cache.scala 96:62]
    .clock(dcache_data_2_clock),
    .io_wen(dcache_data_2_io_wen),
    .io_addr(dcache_data_2_io_addr),
    .io_wdata(dcache_data_2_io_wdata),
    .io_rdata(dcache_data_2_io_rdata),
    .io_sram_addr(dcache_data_2_io_sram_addr),
    .io_sram_wen(dcache_data_2_io_sram_wen),
    .io_sram_wmask(dcache_data_2_io_sram_wmask),
    .io_sram_wdata(dcache_data_2_io_sram_wdata),
    .io_sram_rdata(dcache_data_2_io_sram_rdata)
  );
  ysyx_22040886_dcache_data dcache_data_3 ( // @[data_cache.scala 96:62]
    .clock(dcache_data_3_clock),
    .io_wen(dcache_data_3_io_wen),
    .io_addr(dcache_data_3_io_addr),
    .io_wdata(dcache_data_3_io_wdata),
    .io_rdata(dcache_data_3_io_rdata),
    .io_sram_addr(dcache_data_3_io_sram_addr),
    .io_sram_wen(dcache_data_3_io_sram_wen),
    .io_sram_wmask(dcache_data_3_io_sram_wmask),
    .io_sram_wdata(dcache_data_3_io_sram_wdata),
    .io_sram_rdata(dcache_data_3_io_sram_rdata)
  );
  assign io_port_araddr = work_state == 5'h1 ? stage1_sram_phy_addr_reg : _io_port_araddr_T_6; // @[data_cache.scala 406:26]
  assign io_port_arlen = {{7'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 408:20]
  assign io_port_arsize = stage1_sram_cache_reg ? 3'h3 : stage1_sram_size_reg; // @[data_cache.scala 409:27]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 413:21]
  assign io_port_arvalid = (_io_port_araddr_T | _io_port_araddr_T_1 | _io_port_araddr_T_2) & _io_port_arvalid_T_7; // @[data_cache.scala 430:27]
  assign io_port_awaddr = 5'h12 == work_state ? _io_port_awaddr_T_3 : _io_port_awaddr_T_9; // @[Mux.scala 81:58]
  assign io_port_awlen = {{7'd0}, _io_port_awlen_T_2}; // @[data_cache.scala 440:21]
  assign io_port_awsize = _io_port_awlen_T_2 ? 3'h3 : stage1_sram_size_reg; // @[data_cache.scala 441:27]
  assign io_port_awburst = {{1'd0}, _io_port_awlen_T_2}; // @[data_cache.scala 445:21]
  assign io_port_awvalid = _io_port_awvalid_T_4 | _data_cache_under_write_back_T_3; // @[data_cache.scala 450:10]
  assign io_port_wdata = work_state == 5'h4 | _T_35 ? axi_line_wdata : _io_port_wdata_T_14; // @[data_cache.scala 464:26]
  assign io_port_wstrb = _io_port_wdata_T_2 ? stage1_wstrb_reg : _io_port_wstrb_T_14; // @[data_cache.scala 468:26]
  assign io_port_wlast = _io_port_wdata_T | _T_35 & io_port_wready | _io_port_wlast_T_13; // @[data_cache.scala 471:132]
  assign io_port_wvalid = _io_port_wvalid_T_8 | _write_counter_T_9 | _data_cache_under_write_back_T_3 |
    _data_cache_under_write_back_T_5; // @[data_cache.scala 475:136]
  assign io_stage2_stall = access_work_state_for_stall == 2'h3; // @[data_cache.scala 295:48]
  assign io_v_addr_for_tlb = stage1_addr_line_mapping; // @[data_cache.scala 227:23]
  assign io_sram_rdata = stage2_stall_reg ? _io_sram_rdata_T_3 : sram_rdata_reg; // @[data_cache.scala 485:25]
  assign io_sram_0_addr = dcache_data_io_sram_addr; // @[data_cache.scala 95:{36,36}]
  assign io_sram_0_wen = dcache_data_io_sram_wen; // @[data_cache.scala 95:{36,36}]
  assign io_sram_0_wmask = dcache_data_io_sram_wmask; // @[data_cache.scala 95:{36,36}]
  assign io_sram_0_wdata = dcache_data_io_sram_wdata; // @[data_cache.scala 95:{36,36}]
  assign io_sram_1_addr = dcache_data_1_io_sram_addr; // @[data_cache.scala 95:{36,36}]
  assign io_sram_1_wen = dcache_data_1_io_sram_wen; // @[data_cache.scala 95:{36,36}]
  assign io_sram_1_wmask = dcache_data_1_io_sram_wmask; // @[data_cache.scala 95:{36,36}]
  assign io_sram_1_wdata = dcache_data_1_io_sram_wdata; // @[data_cache.scala 95:{36,36}]
  assign io_sram_2_addr = dcache_data_2_io_sram_addr; // @[data_cache.scala 96:{36,36}]
  assign io_sram_2_wen = dcache_data_2_io_sram_wen; // @[data_cache.scala 96:{36,36}]
  assign io_sram_2_wmask = dcache_data_2_io_sram_wmask; // @[data_cache.scala 96:{36,36}]
  assign io_sram_2_wdata = dcache_data_2_io_sram_wdata; // @[data_cache.scala 96:{36,36}]
  assign io_sram_3_addr = dcache_data_3_io_sram_addr; // @[data_cache.scala 96:{36,36}]
  assign io_sram_3_wen = dcache_data_3_io_sram_wen; // @[data_cache.scala 96:{36,36}]
  assign io_sram_3_wmask = dcache_data_3_io_sram_wmask; // @[data_cache.scala 96:{36,36}]
  assign io_sram_3_wdata = dcache_data_3_io_sram_wdata; // @[data_cache.scala 96:{36,36}]
  assign dcache_tag_clock = clock;
  assign dcache_tag_reset = reset;
  assign dcache_tag_io_wen = _way0_burst_read_wen_T_2 & _way0_dirty_T_7; // @[data_cache.scala 396:122]
  assign dcache_tag_io_wdata = _way0_burst_read_wen_T_2 ? _T_27 : 22'h0; // @[data_cache.scala 398:30]
  assign dcache_tag_io_raddr = io_sram_addr; // @[data_cache.scala 221:24]
  assign dcache_tag_io_waddr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 218:30]
  assign dcache_tag_1_clock = clock;
  assign dcache_tag_1_reset = reset;
  assign dcache_tag_1_io_wen = _way0_burst_read_wen_T_2 & _GEN_384; // @[data_cache.scala 397:122]
  assign dcache_tag_1_io_wdata = _way0_burst_read_wen_T_2 ? _T_27 : 22'h0; // @[data_cache.scala 399:30]
  assign dcache_tag_1_io_raddr = io_sram_addr; // @[data_cache.scala 222:24]
  assign dcache_tag_1_io_waddr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 219:30]
  assign dcache_data_clock = clock;
  assign dcache_data_io_wen = ~stage1_addr_line_mapping[3] & (_way0_dirty_T_4 | _way0_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way0_wire_0_T_13; // @[data_cache.scala 380:33]
  assign dcache_data_io_addr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 369:40]
  assign dcache_data_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 370:41]
  assign dcache_data_io_sram_rdata = io_sram_0_rdata; // @[data_cache.scala 100:16 95:36]
  assign dcache_data_1_clock = clock;
  assign dcache_data_1_io_wen = stage1_addr_line_mapping[3] & (_way0_dirty_T_4 | _way0_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way0_wire_1_T_13; // @[data_cache.scala 380:33]
  assign dcache_data_1_io_addr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 369:40]
  assign dcache_data_1_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 370:41]
  assign dcache_data_1_io_sram_rdata = io_sram_1_rdata; // @[data_cache.scala 101:16 95:36]
  assign dcache_data_2_clock = clock;
  assign dcache_data_2_io_wen = _wen_way0_wire_0_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_0_T_13; // @[data_cache.scala 382:33]
  assign dcache_data_2_io_addr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 373:40]
  assign dcache_data_2_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 374:41]
  assign dcache_data_2_io_sram_rdata = io_sram_2_rdata; // @[data_cache.scala 102:16 96:36]
  assign dcache_data_3_clock = clock;
  assign dcache_data_3_io_wen = stage1_addr_line_mapping[3] & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_1_T_13; // @[data_cache.scala 382:33]
  assign dcache_data_3_io_addr = data_cache_under_write_back ? {{21'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 373:40]
  assign dcache_data_3_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 374:41]
  assign dcache_data_3_io_sram_rdata = io_sram_3_rdata; // @[data_cache.scala 103:16 96:36]
  always @(posedge clock) begin
    if (reset) begin // @[data_cache.scala 55:29]
      work_state <= 5'h18; // @[data_cache.scala 55:29]
    end else if (5'h15 == work_state) begin // @[Mux.scala 81:58]
      if (data_all_write_back) begin // @[data_cache.scala 281:41]
        work_state <= 5'h18;
      end else begin
        work_state <= 5'h11;
      end
    end else if (5'h14 == work_state) begin // @[Mux.scala 81:58]
      if (io_port_bvalid) begin // @[data_cache.scala 280:41]
        work_state <= 5'h15;
      end
    end else if (5'h13 == work_state) begin // @[Mux.scala 81:58]
      work_state <= _access_work_state_T_49;
    end else begin
      work_state <= _access_work_state_T_94;
    end
    if (reset) begin // @[data_cache.scala 57:33]
      write_counter <= 3'h0; // @[data_cache.scala 57:33]
    end else if (work_state == 5'ha | work_state == 5'h9) begin // @[data_cache.scala 302:25]
      write_counter <= _write_counter_T_8;
    end else if (work_state == 5'h6 | work_state == 5'hf) begin // @[data_cache.scala 303:12]
      write_counter <= _write_counter_T_8;
    end else if (_data_cache_under_write_back_T_5 | _data_cache_under_write_back_T_3) begin // @[data_cache.scala 304:12]
      write_counter <= _write_counter_T_8;
    end
    if (reset) begin // @[data_cache.scala 58:32]
      read_counter <= 3'h0; // @[data_cache.scala 58:32]
    end else if (_wait_data_T_3) begin // @[data_cache.scala 305:24]
      read_counter <= _read_counter_T_8;
    end else if (work_state == 5'h0) begin // @[data_cache.scala 306:12]
      read_counter <= _read_counter_T_8;
    end
    if (reset) begin // @[data_cache.scala 59:29]
      wait_data <= 64'h0; // @[data_cache.scala 59:29]
    end else if (work_state == 5'h2 & io_port_rvalid) begin // @[data_cache.scala 299:21]
      wait_data <= io_port_rdata;
    end else if (work_state == 5'hd & io_port_rvalid & read_counter == _GEN_3468) begin // @[data_cache.scala 300:12]
      wait_data <= io_port_rdata;
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_0 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_0 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_0 <= _way0_dirty_T_7;
      end else begin
        lru_0 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_1 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_1 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_1 <= _way0_dirty_T_7;
      end else begin
        lru_1 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_2 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_2 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_2 <= _way0_dirty_T_7;
      end else begin
        lru_2 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_3 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_3 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_3 <= _way0_dirty_T_7;
      end else begin
        lru_3 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_4 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_4 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_4 <= _way0_dirty_T_7;
      end else begin
        lru_4 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_5 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_5 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_5 <= _way0_dirty_T_7;
      end else begin
        lru_5 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_6 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_6 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_6 <= _way0_dirty_T_7;
      end else begin
        lru_6 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_7 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_7 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_7 <= _way0_dirty_T_7;
      end else begin
        lru_7 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_8 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_8 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_8 <= _way0_dirty_T_7;
      end else begin
        lru_8 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_9 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_9 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_9 <= _way0_dirty_T_7;
      end else begin
        lru_9 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_10 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_10 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_10 <= _way0_dirty_T_7;
      end else begin
        lru_10 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_11 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_11 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_11 <= _way0_dirty_T_7;
      end else begin
        lru_11 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_12 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_12 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_12 <= _way0_dirty_T_7;
      end else begin
        lru_12 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_13 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_13 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_13 <= _way0_dirty_T_7;
      end else begin
        lru_13 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_14 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_14 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_14 <= _way0_dirty_T_7;
      end else begin
        lru_14 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_15 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_15 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_15 <= _way0_dirty_T_7;
      end else begin
        lru_15 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_16 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_16 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_16 <= _way0_dirty_T_7;
      end else begin
        lru_16 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_17 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_17 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_17 <= _way0_dirty_T_7;
      end else begin
        lru_17 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_18 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_18 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_18 <= _way0_dirty_T_7;
      end else begin
        lru_18 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_19 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_19 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_19 <= _way0_dirty_T_7;
      end else begin
        lru_19 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_20 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_20 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_20 <= _way0_dirty_T_7;
      end else begin
        lru_20 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_21 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_21 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_21 <= _way0_dirty_T_7;
      end else begin
        lru_21 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_22 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_22 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_22 <= _way0_dirty_T_7;
      end else begin
        lru_22 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_23 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_23 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_23 <= _way0_dirty_T_7;
      end else begin
        lru_23 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_24 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_24 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_24 <= _way0_dirty_T_7;
      end else begin
        lru_24 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_25 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_25 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_25 <= _way0_dirty_T_7;
      end else begin
        lru_25 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_26 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_26 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_26 <= _way0_dirty_T_7;
      end else begin
        lru_26 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_27 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_27 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_27 <= _way0_dirty_T_7;
      end else begin
        lru_27 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_28 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_28 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_28 <= _way0_dirty_T_7;
      end else begin
        lru_28 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_29 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_29 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_29 <= _way0_dirty_T_7;
      end else begin
        lru_29 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_30 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_30 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_30 <= _way0_dirty_T_7;
      end else begin
        lru_30 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_31 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_31 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_31 <= _way0_dirty_T_7;
      end else begin
        lru_31 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_32 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_32 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_32 <= _way0_dirty_T_7;
      end else begin
        lru_32 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_33 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_33 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_33 <= _way0_dirty_T_7;
      end else begin
        lru_33 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_34 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_34 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_34 <= _way0_dirty_T_7;
      end else begin
        lru_34 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_35 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_35 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_35 <= _way0_dirty_T_7;
      end else begin
        lru_35 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_36 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_36 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_36 <= _way0_dirty_T_7;
      end else begin
        lru_36 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_37 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_37 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_37 <= _way0_dirty_T_7;
      end else begin
        lru_37 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_38 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_38 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_38 <= _way0_dirty_T_7;
      end else begin
        lru_38 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_39 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_39 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_39 <= _way0_dirty_T_7;
      end else begin
        lru_39 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_40 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_40 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_40 <= _way0_dirty_T_7;
      end else begin
        lru_40 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_41 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_41 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_41 <= _way0_dirty_T_7;
      end else begin
        lru_41 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_42 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_42 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_42 <= _way0_dirty_T_7;
      end else begin
        lru_42 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_43 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_43 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_43 <= _way0_dirty_T_7;
      end else begin
        lru_43 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_44 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_44 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_44 <= _way0_dirty_T_7;
      end else begin
        lru_44 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_45 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_45 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_45 <= _way0_dirty_T_7;
      end else begin
        lru_45 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_46 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_46 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_46 <= _way0_dirty_T_7;
      end else begin
        lru_46 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_47 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_47 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_47 <= _way0_dirty_T_7;
      end else begin
        lru_47 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_48 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_48 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_48 <= _way0_dirty_T_7;
      end else begin
        lru_48 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_49 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_49 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_49 <= _way0_dirty_T_7;
      end else begin
        lru_49 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_50 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_50 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_50 <= _way0_dirty_T_7;
      end else begin
        lru_50 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_51 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_51 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_51 <= _way0_dirty_T_7;
      end else begin
        lru_51 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_52 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_52 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_52 <= _way0_dirty_T_7;
      end else begin
        lru_52 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_53 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_53 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_53 <= _way0_dirty_T_7;
      end else begin
        lru_53 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_54 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_54 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_54 <= _way0_dirty_T_7;
      end else begin
        lru_54 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_55 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_55 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_55 <= _way0_dirty_T_7;
      end else begin
        lru_55 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_56 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_56 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_56 <= _way0_dirty_T_7;
      end else begin
        lru_56 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_57 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_57 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_57 <= _way0_dirty_T_7;
      end else begin
        lru_57 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_58 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_58 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_58 <= _way0_dirty_T_7;
      end else begin
        lru_58 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_59 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_59 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_59 <= _way0_dirty_T_7;
      end else begin
        lru_59 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_60 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_60 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_60 <= _way0_dirty_T_7;
      end else begin
        lru_60 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_61 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_61 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_61 <= _way0_dirty_T_7;
      end else begin
        lru_61 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_62 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_62 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_62 <= _way0_dirty_T_7;
      end else begin
        lru_62 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_63 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_63 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_63 <= _way0_dirty_T_7;
      end else begin
        lru_63 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_64 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_64 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_64 <= _way0_dirty_T_7;
      end else begin
        lru_64 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_65 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_65 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_65 <= _way0_dirty_T_7;
      end else begin
        lru_65 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_66 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_66 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_66 <= _way0_dirty_T_7;
      end else begin
        lru_66 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_67 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_67 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_67 <= _way0_dirty_T_7;
      end else begin
        lru_67 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_68 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_68 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_68 <= _way0_dirty_T_7;
      end else begin
        lru_68 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_69 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_69 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_69 <= _way0_dirty_T_7;
      end else begin
        lru_69 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_70 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_70 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_70 <= _way0_dirty_T_7;
      end else begin
        lru_70 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_71 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_71 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_71 <= _way0_dirty_T_7;
      end else begin
        lru_71 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_72 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_72 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_72 <= _way0_dirty_T_7;
      end else begin
        lru_72 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_73 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_73 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_73 <= _way0_dirty_T_7;
      end else begin
        lru_73 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_74 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_74 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_74 <= _way0_dirty_T_7;
      end else begin
        lru_74 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_75 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_75 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_75 <= _way0_dirty_T_7;
      end else begin
        lru_75 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_76 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_76 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_76 <= _way0_dirty_T_7;
      end else begin
        lru_76 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_77 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_77 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_77 <= _way0_dirty_T_7;
      end else begin
        lru_77 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_78 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_78 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_78 <= _way0_dirty_T_7;
      end else begin
        lru_78 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_79 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_79 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_79 <= _way0_dirty_T_7;
      end else begin
        lru_79 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_80 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_80 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_80 <= _way0_dirty_T_7;
      end else begin
        lru_80 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_81 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_81 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_81 <= _way0_dirty_T_7;
      end else begin
        lru_81 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_82 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_82 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_82 <= _way0_dirty_T_7;
      end else begin
        lru_82 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_83 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_83 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_83 <= _way0_dirty_T_7;
      end else begin
        lru_83 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_84 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_84 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_84 <= _way0_dirty_T_7;
      end else begin
        lru_84 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_85 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_85 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_85 <= _way0_dirty_T_7;
      end else begin
        lru_85 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_86 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_86 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_86 <= _way0_dirty_T_7;
      end else begin
        lru_86 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_87 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_87 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_87 <= _way0_dirty_T_7;
      end else begin
        lru_87 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_88 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_88 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_88 <= _way0_dirty_T_7;
      end else begin
        lru_88 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_89 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_89 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_89 <= _way0_dirty_T_7;
      end else begin
        lru_89 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_90 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_90 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_90 <= _way0_dirty_T_7;
      end else begin
        lru_90 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_91 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_91 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_91 <= _way0_dirty_T_7;
      end else begin
        lru_91 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_92 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_92 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_92 <= _way0_dirty_T_7;
      end else begin
        lru_92 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_93 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_93 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_93 <= _way0_dirty_T_7;
      end else begin
        lru_93 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_94 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_94 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_94 <= _way0_dirty_T_7;
      end else begin
        lru_94 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_95 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_95 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_95 <= _way0_dirty_T_7;
      end else begin
        lru_95 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_96 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_96 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_96 <= _way0_dirty_T_7;
      end else begin
        lru_96 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_97 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_97 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_97 <= _way0_dirty_T_7;
      end else begin
        lru_97 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_98 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_98 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_98 <= _way0_dirty_T_7;
      end else begin
        lru_98 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_99 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_99 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_99 <= _way0_dirty_T_7;
      end else begin
        lru_99 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_100 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_100 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_100 <= _way0_dirty_T_7;
      end else begin
        lru_100 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_101 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_101 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_101 <= _way0_dirty_T_7;
      end else begin
        lru_101 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_102 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_102 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_102 <= _way0_dirty_T_7;
      end else begin
        lru_102 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_103 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_103 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_103 <= _way0_dirty_T_7;
      end else begin
        lru_103 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_104 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_104 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_104 <= _way0_dirty_T_7;
      end else begin
        lru_104 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_105 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_105 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_105 <= _way0_dirty_T_7;
      end else begin
        lru_105 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_106 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_106 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_106 <= _way0_dirty_T_7;
      end else begin
        lru_106 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_107 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_107 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_107 <= _way0_dirty_T_7;
      end else begin
        lru_107 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_108 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_108 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_108 <= _way0_dirty_T_7;
      end else begin
        lru_108 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_109 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_109 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_109 <= _way0_dirty_T_7;
      end else begin
        lru_109 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_110 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_110 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_110 <= _way0_dirty_T_7;
      end else begin
        lru_110 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_111 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_111 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_111 <= _way0_dirty_T_7;
      end else begin
        lru_111 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_112 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_112 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_112 <= _way0_dirty_T_7;
      end else begin
        lru_112 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_113 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_113 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_113 <= _way0_dirty_T_7;
      end else begin
        lru_113 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_114 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_114 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_114 <= _way0_dirty_T_7;
      end else begin
        lru_114 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_115 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_115 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_115 <= _way0_dirty_T_7;
      end else begin
        lru_115 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_116 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_116 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_116 <= _way0_dirty_T_7;
      end else begin
        lru_116 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_117 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_117 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_117 <= _way0_dirty_T_7;
      end else begin
        lru_117 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_118 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_118 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_118 <= _way0_dirty_T_7;
      end else begin
        lru_118 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_119 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_119 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_119 <= _way0_dirty_T_7;
      end else begin
        lru_119 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_120 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_120 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_120 <= _way0_dirty_T_7;
      end else begin
        lru_120 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_121 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_121 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_121 <= _way0_dirty_T_7;
      end else begin
        lru_121 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_122 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_122 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_122 <= _way0_dirty_T_7;
      end else begin
        lru_122 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_123 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_123 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_123 <= _way0_dirty_T_7;
      end else begin
        lru_123 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_124 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_124 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_124 <= _way0_dirty_T_7;
      end else begin
        lru_124 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_125 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_125 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_125 <= _way0_dirty_T_7;
      end else begin
        lru_125 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_126 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_126 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_126 <= _way0_dirty_T_7;
      end else begin
        lru_126 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 65:22]
      lru_127 <= 1'h0; // @[data_cache.scala 65:22]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 233:37]
      if (_way0_dirty_T) begin // @[data_cache.scala 233:43]
        lru_127 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin // @[data_cache.scala 236:12]
        lru_127 <= _way0_dirty_T_7;
      end else begin
        lru_127 <= _GEN_384;
      end
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_0 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_0 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_1 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_1 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_2 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_2 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_3 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_3 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_4 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_4 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_5 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_5 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_6 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_6 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_7 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_7 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_8 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_8 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_9 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_9 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_10 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_10 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_11 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_11 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_12 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_12 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_13 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_13 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_14 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_14 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_15 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_15 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_16 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_16 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_17 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_17 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_18 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_18 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_19 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_19 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_20 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_20 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_21 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_21 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_22 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_22 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_23 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_23 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_24 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_24 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_25 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_25 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_26 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_26 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_27 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_27 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_28 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_28 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_29 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_29 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_30 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_30 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_31 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_31 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_32 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_32 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_33 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_33 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_34 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_34 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_35 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_35 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_36 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_36 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_37 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_37 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_38 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_38 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_39 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_39 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_40 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_40 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_41 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_41 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_42 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_42 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_43 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_43 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_44 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_44 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_45 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_45 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_46 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_46 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_47 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_47 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_48 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_48 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_49 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_49 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_50 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_50 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_51 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_51 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_52 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_52 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_53 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_53 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_54 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_54 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_55 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_55 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_56 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_56 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_57 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_57 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_58 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_58 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_59 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_59 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_60 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_60 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_61 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_61 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_62 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_62 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_63 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_63 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_64 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_64 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_65 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_65 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_66 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_66 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_67 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_67 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_68 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_68 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_69 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_69 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_70 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_70 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_71 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_71 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_72 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_72 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_73 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_73 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_74 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_74 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_75 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_75 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_76 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_76 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_77 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_77 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_78 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_78 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_79 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_79 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_80 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_80 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_81 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_81 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_82 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_82 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_83 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_83 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_84 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_84 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_85 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_85 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_86 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_86 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_87 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_87 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_88 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_88 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_89 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_89 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_90 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_90 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_91 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_91 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_92 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_92 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_93 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_93 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_94 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_94 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_95 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_95 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_96 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_96 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_97 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_97 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_98 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_98 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_99 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_99 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_100 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_100 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_101 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_101 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_102 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_102 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_103 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_103 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_104 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_104 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_105 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_105 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_106 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_106 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_107 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_107 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_108 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_108 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_109 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_109 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_110 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_110 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_111 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_111 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_112 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_112 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_113 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_113 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_114 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_114 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_115 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_115 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_116 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_116 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_117 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_117 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_118 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_118 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_119 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_119 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_120 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_120 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_121 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_121 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_122 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_122 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_123 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_123 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_124 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_124 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_125 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_125 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_126 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_126 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 66:29]
      way0_dirty_127 <= 1'h0; // @[data_cache.scala 66:29]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 204:44]
      way0_dirty_127 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15; // @[data_cache.scala 204:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_0 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_0 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_1 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_1 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_2 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_2 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_3 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_3 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_4 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_4 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_5 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_5 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_6 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_6 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_7 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_7 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_8 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_8 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_9 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_9 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_10 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_10 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_11 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_11 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_12 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_12 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_13 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_13 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_14 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_14 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_15 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_15 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_16 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_16 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_17 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_17 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_18 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_18 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_19 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_19 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_20 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_20 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_21 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_21 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_22 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_22 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_23 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_23 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_24 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_24 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_25 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_25 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_26 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_26 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_27 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_27 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_28 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_28 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_29 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_29 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_30 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_30 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_31 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_31 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_32 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_32 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_33 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_33 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_34 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_34 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_35 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_35 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_36 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_36 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_37 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_37 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_38 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_38 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_39 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_39 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_40 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_40 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_41 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_41 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_42 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_42 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_43 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_43 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_44 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_44 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_45 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_45 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_46 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_46 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_47 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_47 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_48 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_48 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_49 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_49 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_50 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_50 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_51 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_51 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_52 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_52 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_53 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_53 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_54 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_54 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_55 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_55 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_56 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_56 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_57 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_57 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_58 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_58 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_59 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_59 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_60 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_60 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_61 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_61 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_62 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_62 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_63 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_63 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_64 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_64 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_65 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_65 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_66 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_66 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_67 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_67 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_68 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_68 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_69 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_69 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_70 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_70 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_71 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_71 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_72 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_72 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_73 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_73 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_74 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_74 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_75 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_75 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_76 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_76 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_77 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_77 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_78 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_78 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_79 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_79 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_80 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_80 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_81 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_81 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_82 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_82 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_83 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_83 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_84 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_84 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_85 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_85 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_86 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_86 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_87 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_87 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_88 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_88 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_89 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_89 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_90 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_90 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_91 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_91 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_92 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_92 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_93 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_93 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_94 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_94 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_95 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_95 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_96 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_96 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_97 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_97 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_98 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_98 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_99 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_99 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_100 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_100 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_101 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_101 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_102 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_102 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_103 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_103 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_104 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_104 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_105 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_105 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_106 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_106 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_107 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_107 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_108 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_108 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_109 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_109 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_110 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_110 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_111 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_111 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_112 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_112 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_113 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_113 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_114 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_114 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_115 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_115 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_116 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_116 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_117 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_117 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_118 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_118 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_119 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_119 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_120 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_120 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_121 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_121 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_122 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_122 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_123 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_123 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_124 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_124 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_125 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_125 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_126 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_126 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 67:29]
      way1_dirty_127 <= 1'h0; // @[data_cache.scala 67:29]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 208:44]
      way1_dirty_127 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15; // @[data_cache.scala 208:44]
    end
    if (reset) begin // @[data_cache.scala 71:39]
      stage1_addr_line_mapping <= 32'h0; // @[data_cache.scala 71:39]
    end else if (io_sram_req) begin // @[data_cache.scala 190:32]
      stage1_addr_line_mapping <= io_sram_addr;
    end
    if (reset) begin // @[data_cache.scala 72:40]
      stage1_sram_cache_reg <= 1'h0; // @[data_cache.scala 72:40]
    end else if (io_sram_req) begin // @[data_cache.scala 191:33]
      stage1_sram_cache_reg <= io_sram_cache;
    end
    if (reset) begin // @[data_cache.scala 73:40]
      stage1_sram_wdata_reg <= 64'h0; // @[data_cache.scala 73:40]
    end else if (io_sram_req) begin // @[data_cache.scala 192:33]
      stage1_sram_wdata_reg <= io_sram_wdata;
    end
    if (reset) begin // @[data_cache.scala 74:39]
      stage1_sram_size_reg <= 3'h0; // @[data_cache.scala 74:39]
    end else if (io_sram_req) begin // @[data_cache.scala 193:33]
      stage1_sram_size_reg <= io_sram_size;
    end
    if (reset) begin // @[data_cache.scala 75:37]
      stage1_sram_wr_reg <= 1'h0; // @[data_cache.scala 75:37]
    end else if (io_sram_req) begin // @[data_cache.scala 194:33]
      stage1_sram_wr_reg <= io_sram_wr;
    end
    if (reset) begin // @[data_cache.scala 76:38]
      stage1_sram_req_reg <= 1'h0; // @[data_cache.scala 76:38]
    end else begin
      stage1_sram_req_reg <= io_sram_req | _stage1_sram_req_reg_T_1; // @[data_cache.scala 195:27]
    end
    if (reset) begin // @[data_cache.scala 78:40]
      stage1_sram_hit0_reg <= 1'h0; // @[data_cache.scala 78:40]
    end else if (io_sram_req) begin // @[data_cache.scala 198:32]
      stage1_sram_hit0_reg <= dcache_tag_io_hit;
    end
    if (reset) begin // @[data_cache.scala 79:40]
      stage1_sram_hit1_reg <= 1'h0; // @[data_cache.scala 79:40]
    end else if (io_sram_req) begin // @[data_cache.scala 199:32]
      stage1_sram_hit1_reg <= dcache_tag_1_io_hit;
    end
    if (reset) begin // @[data_cache.scala 80:42]
      stage1_sram_valid0_reg <= 1'h0; // @[data_cache.scala 80:42]
    end else if (io_sram_req) begin // @[data_cache.scala 200:34]
      stage1_sram_valid0_reg <= dcache_tag_io_valid;
    end
    if (reset) begin // @[data_cache.scala 81:42]
      stage1_sram_valid1_reg <= 1'h0; // @[data_cache.scala 81:42]
    end else if (io_sram_req) begin // @[data_cache.scala 201:34]
      stage1_sram_valid1_reg <= dcache_tag_1_io_valid;
    end
    if (reset) begin // @[data_cache.scala 82:35]
      stage1_wstrb_reg <= 8'h0; // @[data_cache.scala 82:35]
    end else if (io_sram_req) begin // @[data_cache.scala 196:33]
      stage1_wstrb_reg <= io_data_wstrb;
    end
    if (reset) begin // @[data_cache.scala 84:43]
      stage1_sram_phy_addr_reg <= 32'h0; // @[data_cache.scala 84:43]
    end else if (stage1_stall_reg) begin // @[data_cache.scala 229:37]
      if (tlb_req) begin // @[data_cache.scala 229:73]
        stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
      end else begin
        stage1_sram_phy_addr_reg <= stage1_addr_line_mapping;
      end
    end
    if (reset) begin // @[data_cache.scala 146:42]
      data_write_back_counter <= 8'h0; // @[data_cache.scala 146:42]
    end else if (_data_write_back_counter_T_2) begin // @[Mux.scala 101:16]
      data_write_back_counter <= _data_write_back_counter_T_4;
    end else if (_data_cache_under_write_back_T_1) begin // @[Mux.scala 101:16]
      data_write_back_counter <= _data_write_back_counter_T_4;
    end
    if (reset) begin // @[data_cache.scala 176:40]
      stage2_sram_write_reg <= 1'h0; // @[data_cache.scala 176:40]
    end else if (stage2_stall) begin // @[data_cache.scala 325:54]
      stage2_sram_write_reg <= stage1_sram_wr_reg;
    end
    if (reset) begin // @[data_cache.scala 183:35]
      stage1_stall_reg <= 1'h0; // @[data_cache.scala 183:35]
    end else begin
      stage1_stall_reg <= io_sram_req; // @[data_cache.scala 184:22]
    end
    if (reset) begin // @[data_cache.scala 186:44]
      write_access_complete_reg <= 1'h0; // @[data_cache.scala 186:44]
    end else begin
      write_access_complete_reg <= _GEN_3339;
    end
    if (reset) begin // @[Reg.scala 28:20]
      stage2_sram_addr_reg <= 32'h0; // @[Reg.scala 28:20]
    end else if (stage2_stall) begin // @[Reg.scala 29:18]
      stage2_sram_addr_reg <= stage1_addr_line_mapping; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[data_cache.scala 328:34]
      stage2_hit0_reg <= 1'h0; // @[data_cache.scala 328:34]
    end else if (stage2_stall) begin // @[data_cache.scala 329:48]
      stage2_hit0_reg <= _hit_T;
    end
    if (reset) begin // @[data_cache.scala 481:33]
      sram_rdata_reg <= 64'h0; // @[data_cache.scala 481:33]
    end else if (_data_cache_under_write_all_back_T) begin // @[data_cache.scala 482:27]
      sram_rdata_reg <= wait_data;
    end else if (_data_cache_under_write_all_back_T_1) begin // @[data_cache.scala 482:73]
      if (stage2_hit0_reg) begin // @[data_cache.scala 353:23]
        sram_rdata_reg <= _GEN_2179;
      end else begin
        sram_rdata_reg <= _GEN_2181;
      end
    end
    if (reset) begin // @[data_cache.scala 483:35]
      stage2_stall_reg <= 1'h0; // @[data_cache.scala 483:35]
    end else begin
      stage2_stall_reg <= stage2_stall; // @[data_cache.scala 484:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  work_state = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  write_counter = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  read_counter = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  wait_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  lru_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_18 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_19 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_20 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_22 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_23 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_24 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_25 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_26 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_27 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_28 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_29 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_30 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_31 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_32 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_33 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_34 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_35 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_36 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_37 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_38 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_39 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_40 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_41 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_42 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_43 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_44 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_45 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_46 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_47 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_48 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_49 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_50 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_51 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_52 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_53 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_54 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_55 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_56 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_57 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_58 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_59 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_60 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_61 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_62 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_63 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_64 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_65 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_66 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_67 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_68 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_69 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_70 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_71 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_72 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_73 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_74 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_75 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_76 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_77 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_78 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_79 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_80 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_81 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_82 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_83 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_84 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_85 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_86 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_87 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_88 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_89 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_90 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_91 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_92 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_93 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_94 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_95 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_96 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_97 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_98 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_99 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_100 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_101 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_102 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_103 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_104 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_105 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_106 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_107 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_108 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_109 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_110 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_111 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_112 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_113 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_114 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_115 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_116 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_117 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_118 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_119 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_120 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_121 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_122 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_123 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  lru_124 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  lru_125 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  lru_126 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  lru_127 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way0_dirty_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way0_dirty_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way0_dirty_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way0_dirty_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way0_dirty_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way0_dirty_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way0_dirty_6 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way0_dirty_7 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way0_dirty_8 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way0_dirty_9 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way0_dirty_10 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way0_dirty_11 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way0_dirty_12 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way0_dirty_13 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way0_dirty_14 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way0_dirty_15 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way0_dirty_16 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way0_dirty_17 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  way0_dirty_18 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  way0_dirty_19 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  way0_dirty_20 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  way0_dirty_21 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  way0_dirty_22 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way0_dirty_23 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way0_dirty_24 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  way0_dirty_25 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  way0_dirty_26 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  way0_dirty_27 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  way0_dirty_28 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  way0_dirty_29 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  way0_dirty_30 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  way0_dirty_31 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  way0_dirty_32 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  way0_dirty_33 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  way0_dirty_34 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  way0_dirty_35 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  way0_dirty_36 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  way0_dirty_37 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  way0_dirty_38 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  way0_dirty_39 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  way0_dirty_40 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  way0_dirty_41 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  way0_dirty_42 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  way0_dirty_43 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  way0_dirty_44 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  way0_dirty_45 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  way0_dirty_46 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  way0_dirty_47 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  way0_dirty_48 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  way0_dirty_49 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  way0_dirty_50 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  way0_dirty_51 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  way0_dirty_52 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  way0_dirty_53 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  way0_dirty_54 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  way0_dirty_55 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  way0_dirty_56 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  way0_dirty_57 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  way0_dirty_58 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  way0_dirty_59 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  way0_dirty_60 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  way0_dirty_61 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  way0_dirty_62 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  way0_dirty_63 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  way0_dirty_64 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  way0_dirty_65 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  way0_dirty_66 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  way0_dirty_67 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  way0_dirty_68 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  way0_dirty_69 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  way0_dirty_70 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  way0_dirty_71 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  way0_dirty_72 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  way0_dirty_73 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  way0_dirty_74 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  way0_dirty_75 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  way0_dirty_76 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  way0_dirty_77 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  way0_dirty_78 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  way0_dirty_79 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  way0_dirty_80 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  way0_dirty_81 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  way0_dirty_82 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  way0_dirty_83 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  way0_dirty_84 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  way0_dirty_85 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  way0_dirty_86 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  way0_dirty_87 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  way0_dirty_88 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  way0_dirty_89 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  way0_dirty_90 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  way0_dirty_91 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  way0_dirty_92 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  way0_dirty_93 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  way0_dirty_94 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  way0_dirty_95 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  way0_dirty_96 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  way0_dirty_97 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  way0_dirty_98 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  way0_dirty_99 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  way0_dirty_100 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  way0_dirty_101 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  way0_dirty_102 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  way0_dirty_103 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  way0_dirty_104 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  way0_dirty_105 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  way0_dirty_106 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  way0_dirty_107 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  way0_dirty_108 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  way0_dirty_109 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  way0_dirty_110 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  way0_dirty_111 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  way0_dirty_112 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  way0_dirty_113 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  way0_dirty_114 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  way0_dirty_115 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  way0_dirty_116 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  way0_dirty_117 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  way0_dirty_118 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  way0_dirty_119 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  way0_dirty_120 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  way0_dirty_121 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  way0_dirty_122 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  way0_dirty_123 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  way0_dirty_124 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  way0_dirty_125 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0_dirty_126 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0_dirty_127 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way1_dirty_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way1_dirty_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way1_dirty_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way1_dirty_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way1_dirty_4 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way1_dirty_5 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way1_dirty_6 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way1_dirty_7 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way1_dirty_8 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way1_dirty_9 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way1_dirty_10 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way1_dirty_11 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way1_dirty_12 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way1_dirty_13 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way1_dirty_14 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way1_dirty_15 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way1_dirty_16 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way1_dirty_17 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way1_dirty_18 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way1_dirty_19 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way1_dirty_20 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way1_dirty_21 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way1_dirty_22 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way1_dirty_23 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way1_dirty_24 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way1_dirty_25 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way1_dirty_26 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way1_dirty_27 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way1_dirty_28 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way1_dirty_29 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way1_dirty_30 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way1_dirty_31 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way1_dirty_32 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way1_dirty_33 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way1_dirty_34 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way1_dirty_35 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way1_dirty_36 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way1_dirty_37 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way1_dirty_38 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way1_dirty_39 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way1_dirty_40 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way1_dirty_41 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way1_dirty_42 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way1_dirty_43 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way1_dirty_44 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way1_dirty_45 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way1_dirty_46 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way1_dirty_47 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way1_dirty_48 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way1_dirty_49 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way1_dirty_50 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way1_dirty_51 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way1_dirty_52 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way1_dirty_53 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way1_dirty_54 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way1_dirty_55 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way1_dirty_56 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way1_dirty_57 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way1_dirty_58 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way1_dirty_59 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way1_dirty_60 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way1_dirty_61 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way1_dirty_62 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way1_dirty_63 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way1_dirty_64 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way1_dirty_65 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way1_dirty_66 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way1_dirty_67 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way1_dirty_68 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way1_dirty_69 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way1_dirty_70 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way1_dirty_71 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way1_dirty_72 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way1_dirty_73 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way1_dirty_74 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way1_dirty_75 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way1_dirty_76 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way1_dirty_77 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way1_dirty_78 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way1_dirty_79 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way1_dirty_80 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way1_dirty_81 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way1_dirty_82 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way1_dirty_83 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way1_dirty_84 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way1_dirty_85 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way1_dirty_86 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way1_dirty_87 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way1_dirty_88 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way1_dirty_89 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way1_dirty_90 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way1_dirty_91 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way1_dirty_92 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way1_dirty_93 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way1_dirty_94 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way1_dirty_95 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way1_dirty_96 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way1_dirty_97 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way1_dirty_98 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way1_dirty_99 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way1_dirty_100 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way1_dirty_101 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way1_dirty_102 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way1_dirty_103 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way1_dirty_104 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way1_dirty_105 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way1_dirty_106 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way1_dirty_107 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way1_dirty_108 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way1_dirty_109 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way1_dirty_110 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way1_dirty_111 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way1_dirty_112 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way1_dirty_113 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way1_dirty_114 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way1_dirty_115 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way1_dirty_116 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way1_dirty_117 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way1_dirty_118 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way1_dirty_119 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way1_dirty_120 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way1_dirty_121 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way1_dirty_122 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way1_dirty_123 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way1_dirty_124 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way1_dirty_125 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way1_dirty_126 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way1_dirty_127 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  stage1_addr_line_mapping = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_389[0:0];
  _RAND_390 = {2{`RANDOM}};
  stage1_sram_wdata_reg = _RAND_390[63:0];
  _RAND_391 = {1{`RANDOM}};
  stage1_sram_size_reg = _RAND_391[2:0];
  _RAND_392 = {1{`RANDOM}};
  stage1_sram_wr_reg = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  stage1_sram_hit0_reg = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  stage1_sram_hit1_reg = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  stage1_sram_valid0_reg = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  stage1_sram_valid1_reg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  stage1_wstrb_reg = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  data_write_back_counter = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  stage2_sram_write_reg = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  write_access_complete_reg = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  stage2_sram_addr_reg = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_405[0:0];
  _RAND_406 = {2{`RANDOM}};
  sram_rdata_reg = _RAND_406[63:0];
  _RAND_407 = {1{`RANDOM}};
  stage2_stall_reg = _RAND_407[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_axi_cross_bar(
  input         clock,
  input         reset,
  input  [31:0] io_m_port_0_araddr,
  input  [7:0]  io_m_port_0_arlen,
  input  [2:0]  io_m_port_0_arsize,
  input  [1:0]  io_m_port_0_arburst,
  input         io_m_port_0_arvalid,
  output        io_m_port_0_arready,
  output [63:0] io_m_port_0_rdata,
  output        io_m_port_0_rlast,
  output        io_m_port_0_rvalid,
  input  [31:0] io_m_port_1_araddr,
  input  [7:0]  io_m_port_1_arlen,
  input  [2:0]  io_m_port_1_arsize,
  input  [1:0]  io_m_port_1_arburst,
  input         io_m_port_1_arvalid,
  output        io_m_port_1_arready,
  output [63:0] io_m_port_1_rdata,
  output        io_m_port_1_rlast,
  output        io_m_port_1_rvalid,
  input  [31:0] io_m_port_1_awaddr,
  input  [7:0]  io_m_port_1_awlen,
  input  [2:0]  io_m_port_1_awsize,
  input  [1:0]  io_m_port_1_awburst,
  input         io_m_port_1_awvalid,
  output        io_m_port_1_awready,
  input  [63:0] io_m_port_1_wdata,
  input  [7:0]  io_m_port_1_wstrb,
  input         io_m_port_1_wlast,
  input         io_m_port_1_wvalid,
  output        io_m_port_1_wready,
  output        io_m_port_1_bvalid,
  output [3:0]  io_s_port_arid,
  output [31:0] io_s_port_araddr,
  output [7:0]  io_s_port_arlen,
  output [2:0]  io_s_port_arsize,
  output [1:0]  io_s_port_arburst,
  output        io_s_port_arvalid,
  input         io_s_port_arready,
  input  [63:0] io_s_port_rdata,
  input         io_s_port_rlast,
  input         io_s_port_rvalid,
  output        io_s_port_rready,
  output [3:0]  io_s_port_awid,
  output [31:0] io_s_port_awaddr,
  output [7:0]  io_s_port_awlen,
  output [2:0]  io_s_port_awsize,
  output [1:0]  io_s_port_awburst,
  output        io_s_port_awvalid,
  input         io_s_port_awready,
  output [63:0] io_s_port_wdata,
  output [7:0]  io_s_port_wstrb,
  output        io_s_port_wlast,
  output        io_s_port_wvalid,
  input         io_s_port_wready,
  input         io_s_port_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  r_inuse_0; // @[axi_ram_port.scala 120:30]
  reg  r_inuse_1; // @[axi_ram_port.scala 120:30]
  reg  w_inuse_1; // @[axi_ram_port.scala 122:30]
  wire [1:0] _T_3 = {w_inuse_1,1'h0}; // @[axi_ram_port.scala 126:93]
  wire  _GEN_4 = io_s_port_bvalid & w_inuse_1 ? 1'h0 : w_inuse_1; // @[axi_ram_port.scala 129:67 130:41 132:41]
  wire  w_inuse_wire_1 = (io_m_port_1_awvalid | io_m_port_1_wvalid) & _T_3 == 2'h0 | _GEN_4; // @[axi_ram_port.scala 126:110 128:41]
  wire [1:0] _w_inuse_0_T = {w_inuse_wire_1,1'h0}; // @[axi_ram_port.scala 140:48]
  wire [1:0] _w_inuse_0_T_6 = 2'h2 - 2'h1; // @[axi_ram_port.scala 140:117]
  wire  _w_inuse_0_T_7 = 2'h0 == _w_inuse_0_T_6; // @[axi_ram_port.scala 140:95]
  wire [1:0] _T_11 = {r_inuse_1,r_inuse_0}; // @[axi_ram_port.scala 142:93]
  wire  _GEN_2 = io_s_port_rlast & r_inuse_0 ? 1'h0 : r_inuse_0; // @[axi_ram_port.scala 144:65 145:41 147:41]
  wire  r_inuse_wire_0 = (io_m_port_0_arvalid | io_m_port_0_rvalid) & _T_11 == 2'h0 | _GEN_2; // @[axi_ram_port.scala 142:110 143:41]
  wire  _GEN_6 = io_s_port_rlast & r_inuse_1 ? 1'h0 : r_inuse_1; // @[axi_ram_port.scala 144:65 145:41 147:41]
  wire  r_inuse_wire_1 = (io_m_port_1_arvalid | io_m_port_1_rvalid) & _T_11 == 2'h0 | _GEN_6; // @[axi_ram_port.scala 142:110 143:41]
  wire [1:0] _r_inuse_0_T = {r_inuse_wire_1,r_inuse_wire_0}; // @[axi_ram_port.scala 157:49]
  wire [1:0] _r_inuse_0_T_3 = {{1'd0}, _r_inuse_0_T[1]}; // @[axi_ram_port.scala 157:56]
  wire  _w_inuse_1_T_7 = 2'h1 == _w_inuse_0_T_6; // @[axi_ram_port.scala 140:95]
  wire [1:0] _r_select_port_T_72 = r_inuse_0 ? io_m_port_0_arburst : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _r_select_port_T_73 = r_inuse_1 ? io_m_port_1_arburst : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _r_select_port_T_75 = r_inuse_0 ? io_m_port_0_arsize : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _r_select_port_T_76 = r_inuse_1 ? io_m_port_1_arsize : 3'h0; // @[Mux.scala 27:73]
  wire [7:0] _r_select_port_T_78 = r_inuse_0 ? io_m_port_0_arlen : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _r_select_port_T_79 = r_inuse_1 ? io_m_port_1_arlen : 8'h0; // @[Mux.scala 27:73]
  wire [31:0] _r_select_port_T_81 = r_inuse_0 ? io_m_port_0_araddr : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _r_select_port_T_82 = r_inuse_1 ? io_m_port_1_araddr : 32'h0; // @[Mux.scala 27:73]
  assign io_m_port_0_arready = r_inuse_0 & io_s_port_arready; // @[axi_ram_port.scala 151:44]
  assign io_m_port_0_rdata = r_inuse_0 ? io_s_port_rdata : 64'h0; // @[axi_ram_port.scala 153:44]
  assign io_m_port_0_rlast = r_inuse_0 & io_s_port_rlast; // @[axi_ram_port.scala 155:44]
  assign io_m_port_0_rvalid = r_inuse_0 & io_s_port_rvalid; // @[axi_ram_port.scala 156:44]
  assign io_m_port_1_arready = r_inuse_1 & io_s_port_arready; // @[axi_ram_port.scala 151:44]
  assign io_m_port_1_rdata = r_inuse_1 ? io_s_port_rdata : 64'h0; // @[axi_ram_port.scala 153:44]
  assign io_m_port_1_rlast = r_inuse_1 & io_s_port_rlast; // @[axi_ram_port.scala 155:44]
  assign io_m_port_1_rvalid = r_inuse_1 & io_s_port_rvalid; // @[axi_ram_port.scala 156:44]
  assign io_m_port_1_awready = w_inuse_1 & io_s_port_awready; // @[axi_ram_port.scala 135:45]
  assign io_m_port_1_wready = w_inuse_1 & io_s_port_wready; // @[axi_ram_port.scala 136:45]
  assign io_m_port_1_bvalid = w_inuse_1 & io_s_port_bvalid; // @[axi_ram_port.scala 139:45]
  assign io_s_port_arid = r_inuse_1 ? 4'h1 : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_araddr = _r_select_port_T_81 | _r_select_port_T_82; // @[Mux.scala 27:73]
  assign io_s_port_arlen = _r_select_port_T_78 | _r_select_port_T_79; // @[Mux.scala 27:73]
  assign io_s_port_arsize = _r_select_port_T_75 | _r_select_port_T_76; // @[Mux.scala 27:73]
  assign io_s_port_arburst = _r_select_port_T_72 | _r_select_port_T_73; // @[Mux.scala 27:73]
  assign io_s_port_arvalid = r_inuse_0 & io_m_port_0_arvalid | r_inuse_1 & io_m_port_1_arvalid; // @[Mux.scala 27:73]
  assign io_s_port_rready = r_inuse_0 | r_inuse_1; // @[Mux.scala 27:73]
  assign io_s_port_awid = w_inuse_1 ? 4'h1 : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_awaddr = w_inuse_1 ? io_m_port_1_awaddr : 32'h0; // @[Mux.scala 27:73]
  assign io_s_port_awlen = w_inuse_1 ? io_m_port_1_awlen : 8'h0; // @[Mux.scala 27:73]
  assign io_s_port_awsize = w_inuse_1 ? io_m_port_1_awsize : 3'h0; // @[Mux.scala 27:73]
  assign io_s_port_awburst = w_inuse_1 ? io_m_port_1_awburst : 2'h0; // @[Mux.scala 27:73]
  assign io_s_port_awvalid = w_inuse_1 & io_m_port_1_awvalid; // @[Mux.scala 27:73]
  assign io_s_port_wdata = w_inuse_1 ? io_m_port_1_wdata : 64'h0; // @[Mux.scala 27:73]
  assign io_s_port_wstrb = w_inuse_1 ? io_m_port_1_wstrb : 8'h0; // @[Mux.scala 27:73]
  assign io_s_port_wlast = w_inuse_1 & io_m_port_1_wlast; // @[Mux.scala 27:73]
  assign io_s_port_wvalid = w_inuse_1 & io_m_port_1_wvalid; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[axi_ram_port.scala 120:30]
      r_inuse_0 <= 1'h0; // @[axi_ram_port.scala 120:30]
    end else begin
      r_inuse_0 <= (_r_inuse_0_T_3 == 2'h0 | _w_inuse_0_T_7) & r_inuse_wire_0; // @[axi_ram_port.scala 157:28]
    end
    if (reset) begin // @[axi_ram_port.scala 120:30]
      r_inuse_1 <= 1'h0; // @[axi_ram_port.scala 120:30]
    end else begin
      r_inuse_1 <= (_r_inuse_0_T == 2'h0 | _w_inuse_1_T_7) & r_inuse_wire_1; // @[axi_ram_port.scala 157:28]
    end
    if (reset) begin // @[axi_ram_port.scala 122:30]
      w_inuse_1 <= 1'h0; // @[axi_ram_port.scala 122:30]
    end else begin
      w_inuse_1 <= (_w_inuse_0_T == 2'h0 | 2'h1 == _w_inuse_0_T_6) & w_inuse_wire_1; // @[axi_ram_port.scala 140:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_inuse_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_inuse_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  w_inuse_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_axi_cross_bar_addr_switch(
  input         clock,
  input         reset,
  input  [31:0] io_m_port_0_araddr,
  input  [7:0]  io_m_port_0_arlen,
  input  [2:0]  io_m_port_0_arsize,
  input  [1:0]  io_m_port_0_arburst,
  input         io_m_port_0_arvalid,
  output        io_m_port_0_arready,
  output [63:0] io_m_port_0_rdata,
  output        io_m_port_0_rlast,
  output        io_m_port_0_rvalid,
  input  [31:0] io_m_port_1_araddr,
  input  [7:0]  io_m_port_1_arlen,
  input  [2:0]  io_m_port_1_arsize,
  input  [1:0]  io_m_port_1_arburst,
  input         io_m_port_1_arvalid,
  output        io_m_port_1_arready,
  output [63:0] io_m_port_1_rdata,
  output        io_m_port_1_rlast,
  output        io_m_port_1_rvalid,
  input  [31:0] io_m_port_1_awaddr,
  input  [7:0]  io_m_port_1_awlen,
  input  [2:0]  io_m_port_1_awsize,
  input  [1:0]  io_m_port_1_awburst,
  input         io_m_port_1_awvalid,
  output        io_m_port_1_awready,
  input  [63:0] io_m_port_1_wdata,
  input  [7:0]  io_m_port_1_wstrb,
  input         io_m_port_1_wlast,
  input         io_m_port_1_wvalid,
  output        io_m_port_1_wready,
  output        io_m_port_1_bvalid,
  output [3:0]  io_s_port_0_arid,
  output [31:0] io_s_port_0_araddr,
  output [7:0]  io_s_port_0_arlen,
  output [2:0]  io_s_port_0_arsize,
  output [1:0]  io_s_port_0_arburst,
  output        io_s_port_0_arvalid,
  input         io_s_port_0_arready,
  input  [63:0] io_s_port_0_rdata,
  input         io_s_port_0_rlast,
  input         io_s_port_0_rvalid,
  output        io_s_port_0_rready,
  output [3:0]  io_s_port_0_awid,
  output [31:0] io_s_port_0_awaddr,
  output [7:0]  io_s_port_0_awlen,
  output [2:0]  io_s_port_0_awsize,
  output [1:0]  io_s_port_0_awburst,
  output        io_s_port_0_awvalid,
  input         io_s_port_0_awready,
  output [63:0] io_s_port_0_wdata,
  output [7:0]  io_s_port_0_wstrb,
  output        io_s_port_0_wlast,
  output        io_s_port_0_wvalid,
  input         io_s_port_0_wready,
  input         io_s_port_0_bvalid,
  output        io_s_port_0_bready,
  output [31:0] io_s_port_1_araddr,
  output        io_s_port_1_arvalid,
  input  [63:0] io_s_port_1_rdata,
  input         io_s_port_1_rlast,
  input         io_s_port_1_rvalid,
  output        io_s_port_1_rready,
  output [31:0] io_s_port_1_awaddr,
  output [2:0]  io_s_port_1_awsize,
  output        io_s_port_1_awvalid,
  output [63:0] io_s_port_1_wdata,
  output        io_s_port_1_wvalid,
  input         io_s_port_1_wready,
  input         io_s_port_1_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_cross_bar_clock; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_reset; // @[axi_ram_port.scala 205:38]
  wire [31:0] axi_cross_bar_io_m_port_0_araddr; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_m_port_0_arlen; // @[axi_ram_port.scala 205:38]
  wire [2:0] axi_cross_bar_io_m_port_0_arsize; // @[axi_ram_port.scala 205:38]
  wire [1:0] axi_cross_bar_io_m_port_0_arburst; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_0_arvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_0_arready; // @[axi_ram_port.scala 205:38]
  wire [63:0] axi_cross_bar_io_m_port_0_rdata; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_0_rlast; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_0_rvalid; // @[axi_ram_port.scala 205:38]
  wire [31:0] axi_cross_bar_io_m_port_1_araddr; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_m_port_1_arlen; // @[axi_ram_port.scala 205:38]
  wire [2:0] axi_cross_bar_io_m_port_1_arsize; // @[axi_ram_port.scala 205:38]
  wire [1:0] axi_cross_bar_io_m_port_1_arburst; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_arvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_arready; // @[axi_ram_port.scala 205:38]
  wire [63:0] axi_cross_bar_io_m_port_1_rdata; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_rlast; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_rvalid; // @[axi_ram_port.scala 205:38]
  wire [31:0] axi_cross_bar_io_m_port_1_awaddr; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_m_port_1_awlen; // @[axi_ram_port.scala 205:38]
  wire [2:0] axi_cross_bar_io_m_port_1_awsize; // @[axi_ram_port.scala 205:38]
  wire [1:0] axi_cross_bar_io_m_port_1_awburst; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_awvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_awready; // @[axi_ram_port.scala 205:38]
  wire [63:0] axi_cross_bar_io_m_port_1_wdata; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_m_port_1_wstrb; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_wlast; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_wvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_wready; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_m_port_1_bvalid; // @[axi_ram_port.scala 205:38]
  wire [3:0] axi_cross_bar_io_s_port_arid; // @[axi_ram_port.scala 205:38]
  wire [31:0] axi_cross_bar_io_s_port_araddr; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_s_port_arlen; // @[axi_ram_port.scala 205:38]
  wire [2:0] axi_cross_bar_io_s_port_arsize; // @[axi_ram_port.scala 205:38]
  wire [1:0] axi_cross_bar_io_s_port_arburst; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_arready; // @[axi_ram_port.scala 205:38]
  wire [63:0] axi_cross_bar_io_s_port_rdata; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_rlast; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_rvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 205:38]
  wire [3:0] axi_cross_bar_io_s_port_awid; // @[axi_ram_port.scala 205:38]
  wire [31:0] axi_cross_bar_io_s_port_awaddr; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_s_port_awlen; // @[axi_ram_port.scala 205:38]
  wire [2:0] axi_cross_bar_io_s_port_awsize; // @[axi_ram_port.scala 205:38]
  wire [1:0] axi_cross_bar_io_s_port_awburst; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_awready; // @[axi_ram_port.scala 205:38]
  wire [63:0] axi_cross_bar_io_s_port_wdata; // @[axi_ram_port.scala 205:38]
  wire [7:0] axi_cross_bar_io_s_port_wstrb; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_wlast; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_wready; // @[axi_ram_port.scala 205:38]
  wire  axi_cross_bar_io_s_port_bvalid; // @[axi_ram_port.scala 205:38]
  reg  select_s_port_num_r_0; // @[axi_ram_port.scala 210:43]
  reg  select_s_port_num_r_1; // @[axi_ram_port.scala 210:43]
  reg  select_s_port_num_w_0; // @[axi_ram_port.scala 211:43]
  reg  select_s_port_num_w_1; // @[axi_ram_port.scala 211:43]
  wire  _access_select_s_port_num_r_1_T = axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 237:98]
  wire [63:0] _GEN_36 = {{32'd0}, axi_cross_bar_io_s_port_araddr}; // @[axi_ram_port.scala 237:137]
  wire  _access_select_s_port_num_r_1_T_2 = _GEN_36 < 64'h200bfff; // @[axi_ram_port.scala 238:64]
  wire  _access_select_s_port_num_r_1_T_3 = _GEN_36 >= 64'h2000000 & _access_select_s_port_num_r_1_T_2; // @[axi_ram_port.scala 237:182]
  wire  access_select_s_port_num_r_1 = axi_cross_bar_io_s_port_arvalid ? _GEN_36 >= 64'h2000000 &
    _access_select_s_port_num_r_1_T_2 : select_s_port_num_r_1; // @[axi_ram_port.scala 237:65]
  wire  _access_select_s_port_num_r_0_T_1 = ~access_select_s_port_num_r_1; // @[axi_ram_port.scala 219:90]
  wire  access_select_s_port_num_r_0 = _access_select_s_port_num_r_1_T ? _access_select_s_port_num_r_0_T_1 :
    select_s_port_num_r_0; // @[axi_ram_port.scala 218:69]
  wire  _access_select_s_port_num_w_1_T = axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 242:98]
  wire [63:0] _GEN_38 = {{32'd0}, axi_cross_bar_io_s_port_awaddr}; // @[axi_ram_port.scala 242:137]
  wire  _access_select_s_port_num_w_1_T_2 = _GEN_38 < 64'h200bfff; // @[axi_ram_port.scala 243:64]
  wire  _access_select_s_port_num_w_1_T_3 = _GEN_38 >= 64'h2000000 & _access_select_s_port_num_w_1_T_2; // @[axi_ram_port.scala 242:180]
  wire  access_select_s_port_num_w_1 = axi_cross_bar_io_s_port_awvalid ? _GEN_38 >= 64'h2000000 &
    _access_select_s_port_num_w_1_T_2 : select_s_port_num_w_1; // @[axi_ram_port.scala 242:65]
  wire  _access_select_s_port_num_w_0_T_1 = ~access_select_s_port_num_w_1; // @[axi_ram_port.scala 223:90]
  wire  access_select_s_port_num_w_0 = _access_select_s_port_num_w_1_T ? _access_select_s_port_num_w_0_T_1 :
    select_s_port_num_w_0; // @[axi_ram_port.scala 222:73]
  wire [63:0] _T_21 = access_select_s_port_num_r_0 ? io_s_port_0_rdata : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_22 = access_select_s_port_num_r_1 ? io_s_port_1_rdata : 64'h0; // @[Mux.scala 27:73]
  ysyx_22040886_axi_cross_bar axi_cross_bar ( // @[axi_ram_port.scala 205:38]
    .clock(axi_cross_bar_clock),
    .reset(axi_cross_bar_reset),
    .io_m_port_0_araddr(axi_cross_bar_io_m_port_0_araddr),
    .io_m_port_0_arlen(axi_cross_bar_io_m_port_0_arlen),
    .io_m_port_0_arsize(axi_cross_bar_io_m_port_0_arsize),
    .io_m_port_0_arburst(axi_cross_bar_io_m_port_0_arburst),
    .io_m_port_0_arvalid(axi_cross_bar_io_m_port_0_arvalid),
    .io_m_port_0_arready(axi_cross_bar_io_m_port_0_arready),
    .io_m_port_0_rdata(axi_cross_bar_io_m_port_0_rdata),
    .io_m_port_0_rlast(axi_cross_bar_io_m_port_0_rlast),
    .io_m_port_0_rvalid(axi_cross_bar_io_m_port_0_rvalid),
    .io_m_port_1_araddr(axi_cross_bar_io_m_port_1_araddr),
    .io_m_port_1_arlen(axi_cross_bar_io_m_port_1_arlen),
    .io_m_port_1_arsize(axi_cross_bar_io_m_port_1_arsize),
    .io_m_port_1_arburst(axi_cross_bar_io_m_port_1_arburst),
    .io_m_port_1_arvalid(axi_cross_bar_io_m_port_1_arvalid),
    .io_m_port_1_arready(axi_cross_bar_io_m_port_1_arready),
    .io_m_port_1_rdata(axi_cross_bar_io_m_port_1_rdata),
    .io_m_port_1_rlast(axi_cross_bar_io_m_port_1_rlast),
    .io_m_port_1_rvalid(axi_cross_bar_io_m_port_1_rvalid),
    .io_m_port_1_awaddr(axi_cross_bar_io_m_port_1_awaddr),
    .io_m_port_1_awlen(axi_cross_bar_io_m_port_1_awlen),
    .io_m_port_1_awsize(axi_cross_bar_io_m_port_1_awsize),
    .io_m_port_1_awburst(axi_cross_bar_io_m_port_1_awburst),
    .io_m_port_1_awvalid(axi_cross_bar_io_m_port_1_awvalid),
    .io_m_port_1_awready(axi_cross_bar_io_m_port_1_awready),
    .io_m_port_1_wdata(axi_cross_bar_io_m_port_1_wdata),
    .io_m_port_1_wstrb(axi_cross_bar_io_m_port_1_wstrb),
    .io_m_port_1_wlast(axi_cross_bar_io_m_port_1_wlast),
    .io_m_port_1_wvalid(axi_cross_bar_io_m_port_1_wvalid),
    .io_m_port_1_wready(axi_cross_bar_io_m_port_1_wready),
    .io_m_port_1_bvalid(axi_cross_bar_io_m_port_1_bvalid),
    .io_s_port_arid(axi_cross_bar_io_s_port_arid),
    .io_s_port_araddr(axi_cross_bar_io_s_port_araddr),
    .io_s_port_arlen(axi_cross_bar_io_s_port_arlen),
    .io_s_port_arsize(axi_cross_bar_io_s_port_arsize),
    .io_s_port_arburst(axi_cross_bar_io_s_port_arburst),
    .io_s_port_arvalid(axi_cross_bar_io_s_port_arvalid),
    .io_s_port_arready(axi_cross_bar_io_s_port_arready),
    .io_s_port_rdata(axi_cross_bar_io_s_port_rdata),
    .io_s_port_rlast(axi_cross_bar_io_s_port_rlast),
    .io_s_port_rvalid(axi_cross_bar_io_s_port_rvalid),
    .io_s_port_rready(axi_cross_bar_io_s_port_rready),
    .io_s_port_awid(axi_cross_bar_io_s_port_awid),
    .io_s_port_awaddr(axi_cross_bar_io_s_port_awaddr),
    .io_s_port_awlen(axi_cross_bar_io_s_port_awlen),
    .io_s_port_awsize(axi_cross_bar_io_s_port_awsize),
    .io_s_port_awburst(axi_cross_bar_io_s_port_awburst),
    .io_s_port_awvalid(axi_cross_bar_io_s_port_awvalid),
    .io_s_port_awready(axi_cross_bar_io_s_port_awready),
    .io_s_port_wdata(axi_cross_bar_io_s_port_wdata),
    .io_s_port_wstrb(axi_cross_bar_io_s_port_wstrb),
    .io_s_port_wlast(axi_cross_bar_io_s_port_wlast),
    .io_s_port_wvalid(axi_cross_bar_io_s_port_wvalid),
    .io_s_port_wready(axi_cross_bar_io_s_port_wready),
    .io_s_port_bvalid(axi_cross_bar_io_s_port_bvalid)
  );
  assign io_m_port_0_arready = axi_cross_bar_io_m_port_0_arready; // @[axi_ram_port.scala 206:34]
  assign io_m_port_0_rdata = axi_cross_bar_io_m_port_0_rdata; // @[axi_ram_port.scala 206:34]
  assign io_m_port_0_rlast = axi_cross_bar_io_m_port_0_rlast; // @[axi_ram_port.scala 206:34]
  assign io_m_port_0_rvalid = axi_cross_bar_io_m_port_0_rvalid; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_arready = axi_cross_bar_io_m_port_1_arready; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_rdata = axi_cross_bar_io_m_port_1_rdata; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_rlast = axi_cross_bar_io_m_port_1_rlast; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_rvalid = axi_cross_bar_io_m_port_1_rvalid; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_awready = axi_cross_bar_io_m_port_1_awready; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_wready = axi_cross_bar_io_m_port_1_wready; // @[axi_ram_port.scala 206:34]
  assign io_m_port_1_bvalid = axi_cross_bar_io_m_port_1_bvalid; // @[axi_ram_port.scala 206:34]
  assign io_s_port_0_arid = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arid : 4'h0; // @[axi_ram_port.scala 282:57 283:51 295:51]
  assign io_s_port_0_araddr = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_araddr : 32'h0; // @[axi_ram_port.scala 282:57 284:51 296:51]
  assign io_s_port_0_arlen = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arlen : 8'h0; // @[axi_ram_port.scala 282:57 285:51 297:51]
  assign io_s_port_0_arsize = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arsize : 3'h0; // @[axi_ram_port.scala 282:57 286:51 298:51]
  assign io_s_port_0_arburst = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arburst : 2'h0; // @[axi_ram_port.scala 282:57 287:51 299:51]
  assign io_s_port_0_arvalid = access_select_s_port_num_r_0 & axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 282:57 291:51 303:51]
  assign io_s_port_0_rready = access_select_s_port_num_r_0 & axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 282:57 292:51 304:51]
  assign io_s_port_0_awid = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awid : 4'h0; // @[axi_ram_port.scala 306:57 307:52 325:52]
  assign io_s_port_0_awaddr = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awaddr : 32'h0; // @[axi_ram_port.scala 306:57 308:52 326:52]
  assign io_s_port_0_awlen = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awlen : 8'h0; // @[axi_ram_port.scala 306:57 309:52 327:52]
  assign io_s_port_0_awsize = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awsize : 3'h0; // @[axi_ram_port.scala 306:57 310:52 328:52]
  assign io_s_port_0_awburst = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awburst : 2'h0; // @[axi_ram_port.scala 306:57 311:52 329:52]
  assign io_s_port_0_awvalid = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 306:57 315:52 333:52]
  assign io_s_port_0_wdata = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_wdata : 64'h0; // @[axi_ram_port.scala 306:57 317:52 335:52]
  assign io_s_port_0_wstrb = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_wstrb : 8'h0; // @[axi_ram_port.scala 306:57 318:52 336:52]
  assign io_s_port_0_wlast = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_wlast; // @[axi_ram_port.scala 306:57 319:52 337:52]
  assign io_s_port_0_wvalid = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 306:57 320:52 338:52]
  assign io_s_port_0_bready = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_bvalid; // @[axi_ram_port.scala 306:57 321:52 339:52]
  assign io_s_port_1_araddr = access_select_s_port_num_r_1 ? axi_cross_bar_io_s_port_araddr : 32'h0; // @[axi_ram_port.scala 282:57 284:51 296:51]
  assign io_s_port_1_arvalid = access_select_s_port_num_r_1 & axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 282:57 291:51 303:51]
  assign io_s_port_1_rready = access_select_s_port_num_r_1 & axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 282:57 292:51 304:51]
  assign io_s_port_1_awaddr = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_awaddr : 32'h0; // @[axi_ram_port.scala 306:57 308:52 326:52]
  assign io_s_port_1_awsize = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_awsize : 3'h0; // @[axi_ram_port.scala 306:57 310:52 328:52]
  assign io_s_port_1_awvalid = access_select_s_port_num_w_1 & axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 306:57 315:52 333:52]
  assign io_s_port_1_wdata = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_wdata : 64'h0; // @[axi_ram_port.scala 306:57 317:52 335:52]
  assign io_s_port_1_wvalid = access_select_s_port_num_w_1 & axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 306:57 320:52 338:52]
  assign axi_cross_bar_clock = clock;
  assign axi_cross_bar_reset = reset;
  assign axi_cross_bar_io_m_port_0_araddr = io_m_port_0_araddr; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_0_arlen = io_m_port_0_arlen; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_0_arsize = io_m_port_0_arsize; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_0_arburst = io_m_port_0_arburst; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_0_arvalid = io_m_port_0_arvalid; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_araddr = io_m_port_1_araddr; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_arlen = io_m_port_1_arlen; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_arsize = io_m_port_1_arsize; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_arburst = io_m_port_1_arburst; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_arvalid = io_m_port_1_arvalid; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_awaddr = io_m_port_1_awaddr; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_awlen = io_m_port_1_awlen; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_awsize = io_m_port_1_awsize; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_awburst = io_m_port_1_awburst; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_awvalid = io_m_port_1_awvalid; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_wdata = io_m_port_1_wdata; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_wstrb = io_m_port_1_wstrb; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_wlast = io_m_port_1_wlast; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_m_port_1_wvalid = io_m_port_1_wvalid; // @[axi_ram_port.scala 206:34]
  assign axi_cross_bar_io_s_port_arready = access_select_s_port_num_r_0 & io_s_port_0_arready |
    access_select_s_port_num_r_1; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_rdata = _T_21 | _T_22; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_rlast = access_select_s_port_num_r_0 & io_s_port_0_rlast | access_select_s_port_num_r_1
     & io_s_port_1_rlast; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_rvalid = access_select_s_port_num_r_0 & io_s_port_0_rvalid |
    access_select_s_port_num_r_1 & io_s_port_1_rvalid; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_awready = access_select_s_port_num_w_0 & io_s_port_0_awready |
    access_select_s_port_num_w_1; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_wready = access_select_s_port_num_w_0 & io_s_port_0_wready |
    access_select_s_port_num_w_1 & io_s_port_1_wready; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_bvalid = access_select_s_port_num_w_0 & io_s_port_0_bvalid |
    access_select_s_port_num_w_1 & io_s_port_1_bvalid; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (reset) begin // @[axi_ram_port.scala 210:43]
      select_s_port_num_r_0 <= 1'h0; // @[axi_ram_port.scala 210:43]
    end else if (access_select_s_port_num_r_1) begin // @[axi_ram_port.scala 217:50]
      select_s_port_num_r_0 <= 1'h0;
    end else begin
      select_s_port_num_r_0 <= 1'h1;
    end
    if (reset) begin // @[axi_ram_port.scala 210:43]
      select_s_port_num_r_1 <= 1'h0; // @[axi_ram_port.scala 210:43]
    end else if (_access_select_s_port_num_r_1_T) begin // @[axi_ram_port.scala 234:42]
      select_s_port_num_r_1 <= _access_select_s_port_num_r_1_T_3;
    end else if (io_s_port_1_rlast) begin // @[axi_ram_port.scala 235:108]
      select_s_port_num_r_1 <= 1'h0;
    end
    if (reset) begin // @[axi_ram_port.scala 211:43]
      select_s_port_num_w_0 <= 1'h0; // @[axi_ram_port.scala 211:43]
    end else if (access_select_s_port_num_w_1) begin // @[axi_ram_port.scala 221:50]
      select_s_port_num_w_0 <= 1'h0;
    end else begin
      select_s_port_num_w_0 <= 1'h1;
    end
    if (reset) begin // @[axi_ram_port.scala 211:43]
      select_s_port_num_w_1 <= 1'h0; // @[axi_ram_port.scala 211:43]
    end else if (_access_select_s_port_num_w_1_T) begin // @[axi_ram_port.scala 239:42]
      select_s_port_num_w_1 <= _access_select_s_port_num_w_1_T_3;
    end else if (io_s_port_1_bvalid) begin // @[axi_ram_port.scala 240:108]
      select_s_port_num_w_1 <= 1'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  select_s_port_num_r_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  select_s_port_num_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  select_s_port_num_w_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  select_s_port_num_w_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886_timer_periph(
  input         clock,
  input         reset,
  input  [31:0] io_axi_port_araddr,
  input         io_axi_port_arvalid,
  output [63:0] io_axi_port_rdata,
  output        io_axi_port_rlast,
  output        io_axi_port_rvalid,
  input         io_axi_port_rready,
  input  [31:0] io_axi_port_awaddr,
  input  [2:0]  io_axi_port_awsize,
  input         io_axi_port_awvalid,
  input  [63:0] io_axi_port_wdata,
  input         io_axi_port_wvalid,
  output        io_axi_port_wready,
  output        io_axi_port_bvalid,
  output        io_int_line
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[clint.scala 25:26]
  reg [63:0] mtimecmp; // @[clint.scala 26:27]
  reg [31:0] msip; // @[clint.scala 27:25]
  reg [2:0] axi_read_state; // @[clint.scala 33:33]
  reg [2:0] axi_write_state; // @[clint.scala 34:34]
  reg [63:0] axi_read_addr; // @[clint.scala 35:32]
  reg [63:0] axi_write_addr; // @[clint.scala 36:33]
  reg [3:0] axi_write_size; // @[clint.scala 37:33]
  wire [2:0] _axi_write_state_T_3 = io_axi_port_awvalid ? 3'h1 : axi_write_state; // @[clint.scala 46:26]
  wire [1:0] _axi_write_size_T_6 = 3'h1 == io_axi_port_awsize ? 2'h2 : {{1'd0}, 3'h0 == io_axi_port_awsize}; // @[Mux.scala 81:58]
  wire [2:0] _axi_write_size_T_8 = 3'h2 == io_axi_port_awsize ? 3'h4 : {{1'd0}, _axi_write_size_T_6}; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_2 = {io_axi_port_wdata[55:0],8'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_4 = {io_axi_port_wdata[47:0],16'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_6 = {io_axi_port_wdata[39:0],24'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_8 = {io_axi_port_wdata[31:0],32'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_10 = {io_axi_port_wdata[23:0],40'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_12 = {io_axi_port_wdata[15:0],48'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_14 = {io_axi_port_wdata[7:0],56'h0}; // @[Cat.scala 31:58]
  wire [63:0] _axi_write_data_T_16 = 3'h1 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_2 : io_axi_port_wdata; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_18 = 3'h2 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_4 : _axi_write_data_T_16; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_20 = 3'h3 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_6 : _axi_write_data_T_18; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_22 = 3'h4 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_8 : _axi_write_data_T_20; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_24 = 3'h5 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_10 : _axi_write_data_T_22; // @[Mux.scala 81:58]
  wire [63:0] _axi_write_data_T_26 = 3'h6 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_12 : _axi_write_data_T_24; // @[Mux.scala 81:58]
  wire [63:0] axi_write_data = 3'h7 == io_axi_port_awaddr[2:0] ? _axi_write_data_T_14 : _axi_write_data_T_26; // @[Mux.scala 81:58]
  wire [31:0] _read_data_T_7 = 64'h2000000 == axi_read_addr ? msip : 32'h0; // @[Mux.scala 81:58]
  wire [63:0] _read_data_T_9 = 64'h200bff8 == axi_read_addr ? mtime : {{32'd0}, _read_data_T_7}; // @[Mux.scala 81:58]
  wire [3:0] _mtime_to_be_0_T_3 = {1'h0,axi_write_addr[2:0]}; // @[Cat.scala 31:58]
  wire [3:0] _mtime_to_be_0_T_5 = _mtime_to_be_0_T_3 + axi_write_size; // @[clint.scala 83:109]
  wire  _mtime_to_be_0_T_7 = axi_write_addr[2:0] <= 3'h0 & _mtime_to_be_0_T_5 > 4'h0; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_0 = axi_write_addr[2:0] <= 3'h0 & _mtime_to_be_0_T_5 > 4'h0 ? axi_write_data[7:0] : mtime[7:0]; // @[clint.scala 83:38]
  wire  _mtime_to_be_1_T_7 = axi_write_addr[2:0] <= 3'h1 & _mtime_to_be_0_T_5 > 4'h1; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_1 = axi_write_addr[2:0] <= 3'h1 & _mtime_to_be_0_T_5 > 4'h1 ? axi_write_data[15:8] : mtime[15:8
    ]; // @[clint.scala 83:38]
  wire  _mtime_to_be_2_T_7 = axi_write_addr[2:0] <= 3'h2 & _mtime_to_be_0_T_5 > 4'h2; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_2 = axi_write_addr[2:0] <= 3'h2 & _mtime_to_be_0_T_5 > 4'h2 ? axi_write_data[23:16] : mtime[23:
    16]; // @[clint.scala 83:38]
  wire  _mtime_to_be_3_T_7 = axi_write_addr[2:0] <= 3'h3 & _mtime_to_be_0_T_5 > 4'h3; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_3 = axi_write_addr[2:0] <= 3'h3 & _mtime_to_be_0_T_5 > 4'h3 ? axi_write_data[31:24] : mtime[31:
    24]; // @[clint.scala 83:38]
  wire  _mtime_to_be_4_T_7 = axi_write_addr[2:0] <= 3'h4 & _mtime_to_be_0_T_5 > 4'h4; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_4 = axi_write_addr[2:0] <= 3'h4 & _mtime_to_be_0_T_5 > 4'h4 ? axi_write_data[39:32] : mtime[39:
    32]; // @[clint.scala 83:38]
  wire  _mtime_to_be_5_T_7 = axi_write_addr[2:0] <= 3'h5 & _mtime_to_be_0_T_5 > 4'h5; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_5 = axi_write_addr[2:0] <= 3'h5 & _mtime_to_be_0_T_5 > 4'h5 ? axi_write_data[47:40] : mtime[47:
    40]; // @[clint.scala 83:38]
  wire  _mtime_to_be_6_T_7 = axi_write_addr[2:0] <= 3'h6 & _mtime_to_be_0_T_5 > 4'h6; // @[clint.scala 83:70]
  wire [7:0] mtime_to_be_6 = axi_write_addr[2:0] <= 3'h6 & _mtime_to_be_0_T_5 > 4'h6 ? axi_write_data[55:48] : mtime[55:
    48]; // @[clint.scala 83:38]
  wire  _mtime_to_be_7_T_6 = _mtime_to_be_0_T_5 > 4'h7; // @[clint.scala 83:126]
  wire [7:0] mtime_to_be_7 = _mtime_to_be_0_T_5 > 4'h7 ? axi_write_data[63:56] : mtime[63:56]; // @[clint.scala 83:38]
  wire  _mtime_T_2 = axi_write_state == 3'h1 & io_axi_port_wvalid; // @[clint.scala 86:48]
  wire [63:0] _mtime_T_9 = {mtime_to_be_7,mtime_to_be_6,mtime_to_be_5,mtime_to_be_4,mtime_to_be_3,mtime_to_be_2,
    mtime_to_be_1,mtime_to_be_0}; // @[clint.scala 87:21]
  wire [63:0] _mtime_T_11 = mtime + 64'h1; // @[clint.scala 87:34]
  wire [7:0] mtimecmp_to_be_0 = _mtime_to_be_0_T_7 ? axi_write_data[7:0] : mtimecmp[7:0]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_1 = _mtime_to_be_1_T_7 ? axi_write_data[15:8] : mtimecmp[15:8]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_2 = _mtime_to_be_2_T_7 ? axi_write_data[23:16] : mtimecmp[23:16]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_3 = _mtime_to_be_3_T_7 ? axi_write_data[31:24] : mtimecmp[31:24]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_4 = _mtime_to_be_4_T_7 ? axi_write_data[39:32] : mtimecmp[39:32]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_5 = _mtime_to_be_5_T_7 ? axi_write_data[47:40] : mtimecmp[47:40]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_6 = _mtime_to_be_6_T_7 ? axi_write_data[55:48] : mtimecmp[55:48]; // @[clint.scala 90:41]
  wire [7:0] mtimecmp_to_be_7 = _mtime_to_be_7_T_6 ? axi_write_data[63:56] : mtimecmp[63:56]; // @[clint.scala 90:41]
  wire [63:0] _mtimecmp_T_9 = {mtimecmp_to_be_7,mtimecmp_to_be_6,mtimecmp_to_be_5,mtimecmp_to_be_4,mtimecmp_to_be_3,
    mtimecmp_to_be_2,mtimecmp_to_be_1,mtimecmp_to_be_0}; // @[clint.scala 94:24]
  wire [31:0] _msip_T_8 = {31'h0,axi_write_data[0]}; // @[Cat.scala 31:58]
  assign io_axi_port_rdata = 64'h2004000 == axi_read_addr ? mtimecmp : _read_data_T_9; // @[Mux.scala 81:58]
  assign io_axi_port_rlast = axi_read_state == 3'h1 & io_axi_port_rready; // @[clint.scala 74:55]
  assign io_axi_port_rvalid = axi_read_state == 3'h1; // @[clint.scala 75:42]
  assign io_axi_port_wready = axi_write_state == 3'h1; // @[clint.scala 99:45]
  assign io_axi_port_bvalid = axi_write_state == 3'h2; // @[clint.scala 102:45]
  assign io_int_line = mtime >= mtimecmp; // @[clint.scala 104:26]
  always @(posedge clock) begin
    if (reset) begin // @[clint.scala 25:26]
      mtime <= 64'h0; // @[clint.scala 25:26]
    end else if (axi_write_state == 3'h1 & io_axi_port_wvalid & axi_write_addr[63:3] == 61'h4017ff) begin // @[clint.scala 86:17]
      mtime <= _mtime_T_9;
    end else begin
      mtime <= _mtime_T_11;
    end
    if (reset) begin // @[clint.scala 26:27]
      mtimecmp <= 64'h0; // @[clint.scala 26:27]
    end else if (_mtime_T_2 & axi_write_addr[63:3] == 61'h400800) begin // @[clint.scala 93:20]
      mtimecmp <= _mtimecmp_T_9;
    end
    if (reset) begin // @[clint.scala 27:25]
      msip <= 32'h0; // @[clint.scala 27:25]
    end else if (axi_read_addr == 64'h1 & io_axi_port_wvalid & axi_write_addr == 64'h2000000) begin // @[clint.scala 95:16]
      msip <= _msip_T_8;
    end
    if (reset) begin // @[clint.scala 33:33]
      axi_read_state <= 3'h0; // @[clint.scala 33:33]
    end else if (3'h1 == axi_read_state) begin // @[Mux.scala 81:58]
      if (!(io_axi_port_rready)) begin // @[clint.scala 42:26]
        axi_read_state <= 3'h0;
      end
    end else if (3'h0 == axi_read_state) begin // @[Mux.scala 81:58]
      if (io_axi_port_arvalid) begin // @[clint.scala 41:26]
        axi_read_state <= 3'h1;
      end
    end
    if (reset) begin // @[clint.scala 34:34]
      axi_write_state <= 3'h0; // @[clint.scala 34:34]
    end else if (3'h2 == axi_write_state) begin // @[Mux.scala 81:58]
      axi_write_state <= 3'h0;
    end else if (3'h1 == axi_write_state) begin // @[Mux.scala 81:58]
      if (io_axi_port_wready) begin // @[clint.scala 47:26]
        axi_write_state <= 3'h2;
      end
    end else if (3'h0 == axi_write_state) begin // @[Mux.scala 81:58]
      axi_write_state <= _axi_write_state_T_3;
    end
    if (reset) begin // @[clint.scala 35:32]
      axi_read_addr <= 64'h0; // @[clint.scala 35:32]
    end else if (io_axi_port_arvalid) begin // @[clint.scala 51:25]
      axi_read_addr <= {{32'd0}, io_axi_port_araddr};
    end
    if (reset) begin // @[clint.scala 36:33]
      axi_write_addr <= 64'h0; // @[clint.scala 36:33]
    end else if (io_axi_port_awvalid) begin // @[clint.scala 52:26]
      axi_write_addr <= {{32'd0}, io_axi_port_awaddr};
    end
    if (reset) begin // @[clint.scala 37:33]
      axi_write_size <= 4'h0; // @[clint.scala 37:33]
    end else if (io_axi_port_awvalid) begin // @[clint.scala 53:26]
      if (3'h3 == io_axi_port_awsize) begin // @[Mux.scala 81:58]
        axi_write_size <= 4'h8;
      end else begin
        axi_write_size <= {{1'd0}, _axi_write_size_T_8};
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  msip = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  axi_read_state = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  axi_write_state = _RAND_4[2:0];
  _RAND_5 = {2{`RANDOM}};
  axi_read_addr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  axi_write_addr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  axi_write_size = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_22040886(
  input          clock,
  input          reset,
  output [3:0]   io_master_arid,
  output [31:0]  io_master_araddr,
  output [7:0]   io_master_arlen,
  output [2:0]   io_master_arsize,
  output [1:0]   io_master_arburst,
  output         io_master_arvalid,
  input          io_master_arready,
  input  [3:0]   io_master_rid,
  input  [63:0]  io_master_rdata,
  input  [1:0]   io_master_rresp,
  input          io_master_rlast,
  input          io_master_rvalid,
  output         io_master_rready,
  output [3:0]   io_master_awid,
  output [31:0]  io_master_awaddr,
  output [7:0]   io_master_awlen,
  output [2:0]   io_master_awsize,
  output [1:0]   io_master_awburst,
  output         io_master_awvalid,
  input          io_master_awready,
  output [63:0]  io_master_wdata,
  output [7:0]   io_master_wstrb,
  output         io_master_wlast,
  output         io_master_wvalid,
  input          io_master_wready,
  input  [3:0]   io_master_bid,
  input  [1:0]   io_master_bresp,
  input          io_master_bvalid,
  output         io_master_bready,
  input  [3:0]   io_slave_arid,
  input  [31:0]  io_slave_araddr,
  input  [7:0]   io_slave_arlen,
  input  [2:0]   io_slave_arsize,
  input  [1:0]   io_slave_arburst,
  input          io_slave_arvalid,
  output         io_slave_arready,
  output [3:0]   io_slave_rid,
  output [63:0]  io_slave_rdata,
  output [1:0]   io_slave_rresp,
  output         io_slave_rlast,
  output         io_slave_rvalid,
  input          io_slave_rready,
  input  [3:0]   io_slave_awid,
  input  [31:0]  io_slave_awaddr,
  input  [7:0]   io_slave_awlen,
  input  [2:0]   io_slave_awsize,
  input  [1:0]   io_slave_awburst,
  input          io_slave_awvalid,
  output         io_slave_awready,
  input  [63:0]  io_slave_wdata,
  input  [7:0]   io_slave_wstrb,
  input          io_slave_wlast,
  input          io_slave_wvalid,
  output         io_slave_wready,
  output [3:0]   io_slave_bid,
  output [1:0]   io_slave_bresp,
  output         io_slave_bvalid,
  input          io_slave_bready,
  input          io_interrupt,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wmask,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wmask,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wmask,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wmask,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wmask,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wmask,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wmask,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wmask,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata
);
  wire  u_riscv_cpu_clock; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_reset; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_ext_int_timer; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_ext_int_out_int; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_inst_cache; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_inst_sram_en; // @[my_cpu_top.scala 139:29]
  wire [63:0] u_riscv_cpu_inst_sram_addr; // @[my_cpu_top.scala 139:29]
  wire [39:0] u_riscv_cpu_inst_sram_rdata_L; // @[my_cpu_top.scala 139:29]
  wire [1:0] u_riscv_cpu_inst_write_en; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_stage2_flush; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_stage2_stall; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_stage1_valid_flush; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_inst_ready_to_use; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_inst_buffer_full; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_data_sram_en; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_data_sram_wen; // @[my_cpu_top.scala 139:29]
  wire [1:0] u_riscv_cpu_data_size; // @[my_cpu_top.scala 139:29]
  wire [31:0] u_riscv_cpu_data_sram_addr; // @[my_cpu_top.scala 139:29]
  wire [63:0] u_riscv_cpu_data_sram_wdata; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_data_cache; // @[my_cpu_top.scala 139:29]
  wire [63:0] u_riscv_cpu_data_sram_rdata; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_data_stage2_stall; // @[my_cpu_top.scala 139:29]
  wire [7:0] u_riscv_cpu_data_wstrb; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_data_fence_i_control; // @[my_cpu_top.scala 139:29]
  wire  u_riscv_cpu_icache_tag_flush; // @[my_cpu_top.scala 139:29]
  wire  inst_cache_clock; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_reset; // @[my_cpu_top.scala 140:30]
  wire [31:0] inst_cache_io_port_araddr; // @[my_cpu_top.scala 140:30]
  wire [7:0] inst_cache_io_port_arlen; // @[my_cpu_top.scala 140:30]
  wire [2:0] inst_cache_io_port_arsize; // @[my_cpu_top.scala 140:30]
  wire [1:0] inst_cache_io_port_arburst; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_port_arvalid; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_port_arready; // @[my_cpu_top.scala 140:30]
  wire [63:0] inst_cache_io_port_rdata; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_port_rlast; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_port_rvalid; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_stage2_flush; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_stage2_stall; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_stage1_valid_flush; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_inst_ready_to_use; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_inst_buffer_full; // @[my_cpu_top.scala 140:30]
  wire [63:0] inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 140:30]
  wire [63:0] inst_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_req; // @[my_cpu_top.scala 140:30]
  wire [63:0] inst_cache_io_sram_addr; // @[my_cpu_top.scala 140:30]
  wire [1:0] inst_cache_io_sram_write_en; // @[my_cpu_top.scala 140:30]
  wire [39:0] inst_cache_io_sram_rdata_L; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_cache; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_tag_valid_flush; // @[my_cpu_top.scala 140:30]
  wire [5:0] inst_cache_io_sram_0_addr; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_0_wen; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_0_wmask; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_0_wdata; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_0_rdata; // @[my_cpu_top.scala 140:30]
  wire [5:0] inst_cache_io_sram_1_addr; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_1_wen; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_1_wmask; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_1_wdata; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_1_rdata; // @[my_cpu_top.scala 140:30]
  wire [5:0] inst_cache_io_sram_2_addr; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_2_wen; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_2_wmask; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_2_wdata; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_2_rdata; // @[my_cpu_top.scala 140:30]
  wire [5:0] inst_cache_io_sram_3_addr; // @[my_cpu_top.scala 140:30]
  wire  inst_cache_io_sram_3_wen; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_3_wmask; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_3_wdata; // @[my_cpu_top.scala 140:30]
  wire [127:0] inst_cache_io_sram_3_rdata; // @[my_cpu_top.scala 140:30]
  wire  data_cache_clock; // @[my_cpu_top.scala 142:30]
  wire  data_cache_reset; // @[my_cpu_top.scala 142:30]
  wire [31:0] data_cache_io_port_araddr; // @[my_cpu_top.scala 142:30]
  wire [7:0] data_cache_io_port_arlen; // @[my_cpu_top.scala 142:30]
  wire [2:0] data_cache_io_port_arsize; // @[my_cpu_top.scala 142:30]
  wire [1:0] data_cache_io_port_arburst; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_arvalid; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_arready; // @[my_cpu_top.scala 142:30]
  wire [63:0] data_cache_io_port_rdata; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_rlast; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_rvalid; // @[my_cpu_top.scala 142:30]
  wire [31:0] data_cache_io_port_awaddr; // @[my_cpu_top.scala 142:30]
  wire [7:0] data_cache_io_port_awlen; // @[my_cpu_top.scala 142:30]
  wire [2:0] data_cache_io_port_awsize; // @[my_cpu_top.scala 142:30]
  wire [1:0] data_cache_io_port_awburst; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_awvalid; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_awready; // @[my_cpu_top.scala 142:30]
  wire [63:0] data_cache_io_port_wdata; // @[my_cpu_top.scala 142:30]
  wire [7:0] data_cache_io_port_wstrb; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_wlast; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_wvalid; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_wready; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_port_bvalid; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_stage2_stall; // @[my_cpu_top.scala 142:30]
  wire [31:0] data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 142:30]
  wire [31:0] data_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 142:30]
  wire [7:0] data_cache_io_data_wstrb; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_req; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_wr; // @[my_cpu_top.scala 142:30]
  wire [2:0] data_cache_io_sram_size; // @[my_cpu_top.scala 142:30]
  wire [31:0] data_cache_io_sram_addr; // @[my_cpu_top.scala 142:30]
  wire [63:0] data_cache_io_sram_wdata; // @[my_cpu_top.scala 142:30]
  wire [63:0] data_cache_io_sram_rdata; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_cache; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_fence_i_control; // @[my_cpu_top.scala 142:30]
  wire [5:0] data_cache_io_sram_0_addr; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_0_wen; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_0_wmask; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_0_wdata; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_0_rdata; // @[my_cpu_top.scala 142:30]
  wire [5:0] data_cache_io_sram_1_addr; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_1_wen; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_1_wmask; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_1_wdata; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_1_rdata; // @[my_cpu_top.scala 142:30]
  wire [5:0] data_cache_io_sram_2_addr; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_2_wen; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_2_wmask; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_2_wdata; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_2_rdata; // @[my_cpu_top.scala 142:30]
  wire [5:0] data_cache_io_sram_3_addr; // @[my_cpu_top.scala 142:30]
  wire  data_cache_io_sram_3_wen; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_3_wmask; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_3_wdata; // @[my_cpu_top.scala 142:30]
  wire [127:0] data_cache_io_sram_3_rdata; // @[my_cpu_top.scala 142:30]
  wire  _axi_cross_bar_clock; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_reset; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_m_port_0_araddr; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_m_port_0_arlen; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_m_port_0_arsize; // @[my_cpu_top.scala 144:32]
  wire [1:0] _axi_cross_bar_io_m_port_0_arburst; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_0_arvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_0_arready; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_m_port_0_rdata; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_0_rlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_0_rvalid; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_m_port_1_araddr; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_m_port_1_arlen; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_m_port_1_arsize; // @[my_cpu_top.scala 144:32]
  wire [1:0] _axi_cross_bar_io_m_port_1_arburst; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_arvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_arready; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_rdata; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_rlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_rvalid; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_m_port_1_awaddr; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_m_port_1_awlen; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_m_port_1_awsize; // @[my_cpu_top.scala 144:32]
  wire [1:0] _axi_cross_bar_io_m_port_1_awburst; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_awvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_awready; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_wdata; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_m_port_1_wstrb; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_wlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_wvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_wready; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_m_port_1_bvalid; // @[my_cpu_top.scala 144:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_arid; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_s_port_0_araddr; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_s_port_0_arlen; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_s_port_0_arsize; // @[my_cpu_top.scala 144:32]
  wire [1:0] _axi_cross_bar_io_s_port_0_arburst; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_arvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_arready; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_rdata; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_rlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_rvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_rready; // @[my_cpu_top.scala 144:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_awid; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_s_port_0_awaddr; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_s_port_0_awlen; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_s_port_0_awsize; // @[my_cpu_top.scala 144:32]
  wire [1:0] _axi_cross_bar_io_s_port_0_awburst; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_awvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_awready; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_wdata; // @[my_cpu_top.scala 144:32]
  wire [7:0] _axi_cross_bar_io_s_port_0_wstrb; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_wlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_wvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_wready; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_bvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_0_bready; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_s_port_1_araddr; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_arvalid; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_rdata; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_rlast; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_rvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_rready; // @[my_cpu_top.scala 144:32]
  wire [31:0] _axi_cross_bar_io_s_port_1_awaddr; // @[my_cpu_top.scala 144:32]
  wire [2:0] _axi_cross_bar_io_s_port_1_awsize; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_awvalid; // @[my_cpu_top.scala 144:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_wdata; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_wvalid; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_wready; // @[my_cpu_top.scala 144:32]
  wire  _axi_cross_bar_io_s_port_1_bvalid; // @[my_cpu_top.scala 144:32]
  wire  timer_periph_clock; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_reset; // @[my_cpu_top.scala 252:27]
  wire [31:0] timer_periph_io_axi_port_araddr; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_arvalid; // @[my_cpu_top.scala 252:27]
  wire [63:0] timer_periph_io_axi_port_rdata; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_rlast; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_rvalid; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_rready; // @[my_cpu_top.scala 252:27]
  wire [31:0] timer_periph_io_axi_port_awaddr; // @[my_cpu_top.scala 252:27]
  wire [2:0] timer_periph_io_axi_port_awsize; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_awvalid; // @[my_cpu_top.scala 252:27]
  wire [63:0] timer_periph_io_axi_port_wdata; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_wvalid; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_wready; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_axi_port_bvalid; // @[my_cpu_top.scala 252:27]
  wire  timer_periph_io_int_line; // @[my_cpu_top.scala 252:27]
  ysyx_22040886_lys_cpu u_riscv_cpu ( // @[my_cpu_top.scala 139:29]
    .clock(u_riscv_cpu_clock),
    .reset(u_riscv_cpu_reset),
    .ext_int_timer(u_riscv_cpu_ext_int_timer),
    .ext_int_out_int(u_riscv_cpu_ext_int_out_int),
    .inst_cache(u_riscv_cpu_inst_cache),
    .inst_sram_en(u_riscv_cpu_inst_sram_en),
    .inst_sram_addr(u_riscv_cpu_inst_sram_addr),
    .inst_sram_rdata_L(u_riscv_cpu_inst_sram_rdata_L),
    .inst_write_en(u_riscv_cpu_inst_write_en),
    .stage2_flush(u_riscv_cpu_stage2_flush),
    .stage2_stall(u_riscv_cpu_stage2_stall),
    .stage1_valid_flush(u_riscv_cpu_stage1_valid_flush),
    .inst_ready_to_use(u_riscv_cpu_inst_ready_to_use),
    .inst_buffer_full(u_riscv_cpu_inst_buffer_full),
    .data_sram_en(u_riscv_cpu_data_sram_en),
    .data_sram_wen(u_riscv_cpu_data_sram_wen),
    .data_size(u_riscv_cpu_data_size),
    .data_sram_addr(u_riscv_cpu_data_sram_addr),
    .data_sram_wdata(u_riscv_cpu_data_sram_wdata),
    .data_cache(u_riscv_cpu_data_cache),
    .data_sram_rdata(u_riscv_cpu_data_sram_rdata),
    .data_stage2_stall(u_riscv_cpu_data_stage2_stall),
    .data_wstrb(u_riscv_cpu_data_wstrb),
    .data_fence_i_control(u_riscv_cpu_data_fence_i_control),
    .icache_tag_flush(u_riscv_cpu_icache_tag_flush)
  );
  ysyx_22040886_inst_cache inst_cache ( // @[my_cpu_top.scala 140:30]
    .clock(inst_cache_clock),
    .reset(inst_cache_reset),
    .io_port_araddr(inst_cache_io_port_araddr),
    .io_port_arlen(inst_cache_io_port_arlen),
    .io_port_arsize(inst_cache_io_port_arsize),
    .io_port_arburst(inst_cache_io_port_arburst),
    .io_port_arvalid(inst_cache_io_port_arvalid),
    .io_port_arready(inst_cache_io_port_arready),
    .io_port_rdata(inst_cache_io_port_rdata),
    .io_port_rlast(inst_cache_io_port_rlast),
    .io_port_rvalid(inst_cache_io_port_rvalid),
    .io_stage2_flush(inst_cache_io_stage2_flush),
    .io_stage2_stall(inst_cache_io_stage2_stall),
    .io_stage1_valid_flush(inst_cache_io_stage1_valid_flush),
    .io_inst_ready_to_use(inst_cache_io_inst_ready_to_use),
    .io_inst_buffer_full(inst_cache_io_inst_buffer_full),
    .io_v_addr_for_tlb(inst_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(inst_cache_io_p_addr_for_tlb),
    .io_sram_req(inst_cache_io_sram_req),
    .io_sram_addr(inst_cache_io_sram_addr),
    .io_sram_write_en(inst_cache_io_sram_write_en),
    .io_sram_rdata_L(inst_cache_io_sram_rdata_L),
    .io_sram_cache(inst_cache_io_sram_cache),
    .io_tag_valid_flush(inst_cache_io_tag_valid_flush),
    .io_sram_0_addr(inst_cache_io_sram_0_addr),
    .io_sram_0_wen(inst_cache_io_sram_0_wen),
    .io_sram_0_wmask(inst_cache_io_sram_0_wmask),
    .io_sram_0_wdata(inst_cache_io_sram_0_wdata),
    .io_sram_0_rdata(inst_cache_io_sram_0_rdata),
    .io_sram_1_addr(inst_cache_io_sram_1_addr),
    .io_sram_1_wen(inst_cache_io_sram_1_wen),
    .io_sram_1_wmask(inst_cache_io_sram_1_wmask),
    .io_sram_1_wdata(inst_cache_io_sram_1_wdata),
    .io_sram_1_rdata(inst_cache_io_sram_1_rdata),
    .io_sram_2_addr(inst_cache_io_sram_2_addr),
    .io_sram_2_wen(inst_cache_io_sram_2_wen),
    .io_sram_2_wmask(inst_cache_io_sram_2_wmask),
    .io_sram_2_wdata(inst_cache_io_sram_2_wdata),
    .io_sram_2_rdata(inst_cache_io_sram_2_rdata),
    .io_sram_3_addr(inst_cache_io_sram_3_addr),
    .io_sram_3_wen(inst_cache_io_sram_3_wen),
    .io_sram_3_wmask(inst_cache_io_sram_3_wmask),
    .io_sram_3_wdata(inst_cache_io_sram_3_wdata),
    .io_sram_3_rdata(inst_cache_io_sram_3_rdata)
  );
  ysyx_22040886_data_cache data_cache ( // @[my_cpu_top.scala 142:30]
    .clock(data_cache_clock),
    .reset(data_cache_reset),
    .io_port_araddr(data_cache_io_port_araddr),
    .io_port_arlen(data_cache_io_port_arlen),
    .io_port_arsize(data_cache_io_port_arsize),
    .io_port_arburst(data_cache_io_port_arburst),
    .io_port_arvalid(data_cache_io_port_arvalid),
    .io_port_arready(data_cache_io_port_arready),
    .io_port_rdata(data_cache_io_port_rdata),
    .io_port_rlast(data_cache_io_port_rlast),
    .io_port_rvalid(data_cache_io_port_rvalid),
    .io_port_awaddr(data_cache_io_port_awaddr),
    .io_port_awlen(data_cache_io_port_awlen),
    .io_port_awsize(data_cache_io_port_awsize),
    .io_port_awburst(data_cache_io_port_awburst),
    .io_port_awvalid(data_cache_io_port_awvalid),
    .io_port_awready(data_cache_io_port_awready),
    .io_port_wdata(data_cache_io_port_wdata),
    .io_port_wstrb(data_cache_io_port_wstrb),
    .io_port_wlast(data_cache_io_port_wlast),
    .io_port_wvalid(data_cache_io_port_wvalid),
    .io_port_wready(data_cache_io_port_wready),
    .io_port_bvalid(data_cache_io_port_bvalid),
    .io_stage2_stall(data_cache_io_stage2_stall),
    .io_v_addr_for_tlb(data_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(data_cache_io_p_addr_for_tlb),
    .io_data_wstrb(data_cache_io_data_wstrb),
    .io_sram_req(data_cache_io_sram_req),
    .io_sram_wr(data_cache_io_sram_wr),
    .io_sram_size(data_cache_io_sram_size),
    .io_sram_addr(data_cache_io_sram_addr),
    .io_sram_wdata(data_cache_io_sram_wdata),
    .io_sram_rdata(data_cache_io_sram_rdata),
    .io_sram_cache(data_cache_io_sram_cache),
    .io_fence_i_control(data_cache_io_fence_i_control),
    .io_sram_0_addr(data_cache_io_sram_0_addr),
    .io_sram_0_wen(data_cache_io_sram_0_wen),
    .io_sram_0_wmask(data_cache_io_sram_0_wmask),
    .io_sram_0_wdata(data_cache_io_sram_0_wdata),
    .io_sram_0_rdata(data_cache_io_sram_0_rdata),
    .io_sram_1_addr(data_cache_io_sram_1_addr),
    .io_sram_1_wen(data_cache_io_sram_1_wen),
    .io_sram_1_wmask(data_cache_io_sram_1_wmask),
    .io_sram_1_wdata(data_cache_io_sram_1_wdata),
    .io_sram_1_rdata(data_cache_io_sram_1_rdata),
    .io_sram_2_addr(data_cache_io_sram_2_addr),
    .io_sram_2_wen(data_cache_io_sram_2_wen),
    .io_sram_2_wmask(data_cache_io_sram_2_wmask),
    .io_sram_2_wdata(data_cache_io_sram_2_wdata),
    .io_sram_2_rdata(data_cache_io_sram_2_rdata),
    .io_sram_3_addr(data_cache_io_sram_3_addr),
    .io_sram_3_wen(data_cache_io_sram_3_wen),
    .io_sram_3_wmask(data_cache_io_sram_3_wmask),
    .io_sram_3_wdata(data_cache_io_sram_3_wdata),
    .io_sram_3_rdata(data_cache_io_sram_3_rdata)
  );
  ysyx_22040886_axi_cross_bar_addr_switch _axi_cross_bar ( // @[my_cpu_top.scala 144:32]
    .clock(_axi_cross_bar_clock),
    .reset(_axi_cross_bar_reset),
    .io_m_port_0_araddr(_axi_cross_bar_io_m_port_0_araddr),
    .io_m_port_0_arlen(_axi_cross_bar_io_m_port_0_arlen),
    .io_m_port_0_arsize(_axi_cross_bar_io_m_port_0_arsize),
    .io_m_port_0_arburst(_axi_cross_bar_io_m_port_0_arburst),
    .io_m_port_0_arvalid(_axi_cross_bar_io_m_port_0_arvalid),
    .io_m_port_0_arready(_axi_cross_bar_io_m_port_0_arready),
    .io_m_port_0_rdata(_axi_cross_bar_io_m_port_0_rdata),
    .io_m_port_0_rlast(_axi_cross_bar_io_m_port_0_rlast),
    .io_m_port_0_rvalid(_axi_cross_bar_io_m_port_0_rvalid),
    .io_m_port_1_araddr(_axi_cross_bar_io_m_port_1_araddr),
    .io_m_port_1_arlen(_axi_cross_bar_io_m_port_1_arlen),
    .io_m_port_1_arsize(_axi_cross_bar_io_m_port_1_arsize),
    .io_m_port_1_arburst(_axi_cross_bar_io_m_port_1_arburst),
    .io_m_port_1_arvalid(_axi_cross_bar_io_m_port_1_arvalid),
    .io_m_port_1_arready(_axi_cross_bar_io_m_port_1_arready),
    .io_m_port_1_rdata(_axi_cross_bar_io_m_port_1_rdata),
    .io_m_port_1_rlast(_axi_cross_bar_io_m_port_1_rlast),
    .io_m_port_1_rvalid(_axi_cross_bar_io_m_port_1_rvalid),
    .io_m_port_1_awaddr(_axi_cross_bar_io_m_port_1_awaddr),
    .io_m_port_1_awlen(_axi_cross_bar_io_m_port_1_awlen),
    .io_m_port_1_awsize(_axi_cross_bar_io_m_port_1_awsize),
    .io_m_port_1_awburst(_axi_cross_bar_io_m_port_1_awburst),
    .io_m_port_1_awvalid(_axi_cross_bar_io_m_port_1_awvalid),
    .io_m_port_1_awready(_axi_cross_bar_io_m_port_1_awready),
    .io_m_port_1_wdata(_axi_cross_bar_io_m_port_1_wdata),
    .io_m_port_1_wstrb(_axi_cross_bar_io_m_port_1_wstrb),
    .io_m_port_1_wlast(_axi_cross_bar_io_m_port_1_wlast),
    .io_m_port_1_wvalid(_axi_cross_bar_io_m_port_1_wvalid),
    .io_m_port_1_wready(_axi_cross_bar_io_m_port_1_wready),
    .io_m_port_1_bvalid(_axi_cross_bar_io_m_port_1_bvalid),
    .io_s_port_0_arid(_axi_cross_bar_io_s_port_0_arid),
    .io_s_port_0_araddr(_axi_cross_bar_io_s_port_0_araddr),
    .io_s_port_0_arlen(_axi_cross_bar_io_s_port_0_arlen),
    .io_s_port_0_arsize(_axi_cross_bar_io_s_port_0_arsize),
    .io_s_port_0_arburst(_axi_cross_bar_io_s_port_0_arburst),
    .io_s_port_0_arvalid(_axi_cross_bar_io_s_port_0_arvalid),
    .io_s_port_0_arready(_axi_cross_bar_io_s_port_0_arready),
    .io_s_port_0_rdata(_axi_cross_bar_io_s_port_0_rdata),
    .io_s_port_0_rlast(_axi_cross_bar_io_s_port_0_rlast),
    .io_s_port_0_rvalid(_axi_cross_bar_io_s_port_0_rvalid),
    .io_s_port_0_rready(_axi_cross_bar_io_s_port_0_rready),
    .io_s_port_0_awid(_axi_cross_bar_io_s_port_0_awid),
    .io_s_port_0_awaddr(_axi_cross_bar_io_s_port_0_awaddr),
    .io_s_port_0_awlen(_axi_cross_bar_io_s_port_0_awlen),
    .io_s_port_0_awsize(_axi_cross_bar_io_s_port_0_awsize),
    .io_s_port_0_awburst(_axi_cross_bar_io_s_port_0_awburst),
    .io_s_port_0_awvalid(_axi_cross_bar_io_s_port_0_awvalid),
    .io_s_port_0_awready(_axi_cross_bar_io_s_port_0_awready),
    .io_s_port_0_wdata(_axi_cross_bar_io_s_port_0_wdata),
    .io_s_port_0_wstrb(_axi_cross_bar_io_s_port_0_wstrb),
    .io_s_port_0_wlast(_axi_cross_bar_io_s_port_0_wlast),
    .io_s_port_0_wvalid(_axi_cross_bar_io_s_port_0_wvalid),
    .io_s_port_0_wready(_axi_cross_bar_io_s_port_0_wready),
    .io_s_port_0_bvalid(_axi_cross_bar_io_s_port_0_bvalid),
    .io_s_port_0_bready(_axi_cross_bar_io_s_port_0_bready),
    .io_s_port_1_araddr(_axi_cross_bar_io_s_port_1_araddr),
    .io_s_port_1_arvalid(_axi_cross_bar_io_s_port_1_arvalid),
    .io_s_port_1_rdata(_axi_cross_bar_io_s_port_1_rdata),
    .io_s_port_1_rlast(_axi_cross_bar_io_s_port_1_rlast),
    .io_s_port_1_rvalid(_axi_cross_bar_io_s_port_1_rvalid),
    .io_s_port_1_rready(_axi_cross_bar_io_s_port_1_rready),
    .io_s_port_1_awaddr(_axi_cross_bar_io_s_port_1_awaddr),
    .io_s_port_1_awsize(_axi_cross_bar_io_s_port_1_awsize),
    .io_s_port_1_awvalid(_axi_cross_bar_io_s_port_1_awvalid),
    .io_s_port_1_wdata(_axi_cross_bar_io_s_port_1_wdata),
    .io_s_port_1_wvalid(_axi_cross_bar_io_s_port_1_wvalid),
    .io_s_port_1_wready(_axi_cross_bar_io_s_port_1_wready),
    .io_s_port_1_bvalid(_axi_cross_bar_io_s_port_1_bvalid)
  );
  ysyx_22040886_timer_periph timer_periph ( // @[my_cpu_top.scala 252:27]
    .clock(timer_periph_clock),
    .reset(timer_periph_reset),
    .io_axi_port_araddr(timer_periph_io_axi_port_araddr),
    .io_axi_port_arvalid(timer_periph_io_axi_port_arvalid),
    .io_axi_port_rdata(timer_periph_io_axi_port_rdata),
    .io_axi_port_rlast(timer_periph_io_axi_port_rlast),
    .io_axi_port_rvalid(timer_periph_io_axi_port_rvalid),
    .io_axi_port_rready(timer_periph_io_axi_port_rready),
    .io_axi_port_awaddr(timer_periph_io_axi_port_awaddr),
    .io_axi_port_awsize(timer_periph_io_axi_port_awsize),
    .io_axi_port_awvalid(timer_periph_io_axi_port_awvalid),
    .io_axi_port_wdata(timer_periph_io_axi_port_wdata),
    .io_axi_port_wvalid(timer_periph_io_axi_port_wvalid),
    .io_axi_port_wready(timer_periph_io_axi_port_wready),
    .io_axi_port_bvalid(timer_periph_io_axi_port_bvalid),
    .io_int_line(timer_periph_io_int_line)
  );
  assign io_master_arid = _axi_cross_bar_io_s_port_0_arid; // @[my_cpu_top.scala 246:15]
  assign io_master_araddr = _axi_cross_bar_io_s_port_0_araddr; // @[my_cpu_top.scala 246:15]
  assign io_master_arlen = _axi_cross_bar_io_s_port_0_arlen; // @[my_cpu_top.scala 246:15]
  assign io_master_arsize = _axi_cross_bar_io_s_port_0_arsize; // @[my_cpu_top.scala 246:15]
  assign io_master_arburst = _axi_cross_bar_io_s_port_0_arburst; // @[my_cpu_top.scala 246:15]
  assign io_master_arvalid = _axi_cross_bar_io_s_port_0_arvalid; // @[my_cpu_top.scala 246:15]
  assign io_master_rready = _axi_cross_bar_io_s_port_0_rready; // @[my_cpu_top.scala 246:15]
  assign io_master_awid = _axi_cross_bar_io_s_port_0_awid; // @[my_cpu_top.scala 246:15]
  assign io_master_awaddr = _axi_cross_bar_io_s_port_0_awaddr; // @[my_cpu_top.scala 246:15]
  assign io_master_awlen = _axi_cross_bar_io_s_port_0_awlen; // @[my_cpu_top.scala 246:15]
  assign io_master_awsize = _axi_cross_bar_io_s_port_0_awsize; // @[my_cpu_top.scala 246:15]
  assign io_master_awburst = _axi_cross_bar_io_s_port_0_awburst; // @[my_cpu_top.scala 246:15]
  assign io_master_awvalid = _axi_cross_bar_io_s_port_0_awvalid; // @[my_cpu_top.scala 246:15]
  assign io_master_wdata = _axi_cross_bar_io_s_port_0_wdata; // @[my_cpu_top.scala 246:15]
  assign io_master_wstrb = _axi_cross_bar_io_s_port_0_wstrb; // @[my_cpu_top.scala 246:15]
  assign io_master_wlast = _axi_cross_bar_io_s_port_0_wlast; // @[my_cpu_top.scala 246:15]
  assign io_master_wvalid = _axi_cross_bar_io_s_port_0_wvalid; // @[my_cpu_top.scala 246:15]
  assign io_master_bready = _axi_cross_bar_io_s_port_0_bready; // @[my_cpu_top.scala 246:15]
  assign io_slave_arready = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_rid = 4'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_rdata = 64'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_rresp = 2'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_rlast = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_rvalid = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_awready = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_wready = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_bid = 4'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_bresp = 2'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_slave_bvalid = 1'h0; // @[my_cpu_top.scala 137:{29,29}]
  assign io_sram0_addr = inst_cache_io_sram_0_addr; // @[my_cpu_top.scala 364:14]
  assign io_sram0_cen = 1'h0; // @[my_cpu_top.scala 364:14]
  assign io_sram0_wen = inst_cache_io_sram_0_wen; // @[my_cpu_top.scala 364:14]
  assign io_sram0_wmask = inst_cache_io_sram_0_wmask; // @[my_cpu_top.scala 364:14]
  assign io_sram0_wdata = inst_cache_io_sram_0_wdata; // @[my_cpu_top.scala 364:14]
  assign io_sram1_addr = inst_cache_io_sram_1_addr; // @[my_cpu_top.scala 365:14]
  assign io_sram1_cen = 1'h0; // @[my_cpu_top.scala 365:14]
  assign io_sram1_wen = inst_cache_io_sram_1_wen; // @[my_cpu_top.scala 365:14]
  assign io_sram1_wmask = inst_cache_io_sram_1_wmask; // @[my_cpu_top.scala 365:14]
  assign io_sram1_wdata = inst_cache_io_sram_1_wdata; // @[my_cpu_top.scala 365:14]
  assign io_sram2_addr = inst_cache_io_sram_2_addr; // @[my_cpu_top.scala 366:14]
  assign io_sram2_cen = 1'h0; // @[my_cpu_top.scala 366:14]
  assign io_sram2_wen = inst_cache_io_sram_2_wen; // @[my_cpu_top.scala 366:14]
  assign io_sram2_wmask = inst_cache_io_sram_2_wmask; // @[my_cpu_top.scala 366:14]
  assign io_sram2_wdata = inst_cache_io_sram_2_wdata; // @[my_cpu_top.scala 366:14]
  assign io_sram3_addr = inst_cache_io_sram_3_addr; // @[my_cpu_top.scala 367:14]
  assign io_sram3_cen = 1'h0; // @[my_cpu_top.scala 367:14]
  assign io_sram3_wen = inst_cache_io_sram_3_wen; // @[my_cpu_top.scala 367:14]
  assign io_sram3_wmask = inst_cache_io_sram_3_wmask; // @[my_cpu_top.scala 367:14]
  assign io_sram3_wdata = inst_cache_io_sram_3_wdata; // @[my_cpu_top.scala 367:14]
  assign io_sram4_addr = data_cache_io_sram_0_addr; // @[my_cpu_top.scala 368:14]
  assign io_sram4_cen = 1'h0; // @[my_cpu_top.scala 368:14]
  assign io_sram4_wen = data_cache_io_sram_0_wen; // @[my_cpu_top.scala 368:14]
  assign io_sram4_wmask = data_cache_io_sram_0_wmask; // @[my_cpu_top.scala 368:14]
  assign io_sram4_wdata = data_cache_io_sram_0_wdata; // @[my_cpu_top.scala 368:14]
  assign io_sram5_addr = data_cache_io_sram_1_addr; // @[my_cpu_top.scala 369:14]
  assign io_sram5_cen = 1'h0; // @[my_cpu_top.scala 369:14]
  assign io_sram5_wen = data_cache_io_sram_1_wen; // @[my_cpu_top.scala 369:14]
  assign io_sram5_wmask = data_cache_io_sram_1_wmask; // @[my_cpu_top.scala 369:14]
  assign io_sram5_wdata = data_cache_io_sram_1_wdata; // @[my_cpu_top.scala 369:14]
  assign io_sram6_addr = data_cache_io_sram_2_addr; // @[my_cpu_top.scala 370:14]
  assign io_sram6_cen = 1'h0; // @[my_cpu_top.scala 370:14]
  assign io_sram6_wen = data_cache_io_sram_2_wen; // @[my_cpu_top.scala 370:14]
  assign io_sram6_wmask = data_cache_io_sram_2_wmask; // @[my_cpu_top.scala 370:14]
  assign io_sram6_wdata = data_cache_io_sram_2_wdata; // @[my_cpu_top.scala 370:14]
  assign io_sram7_addr = data_cache_io_sram_3_addr; // @[my_cpu_top.scala 371:14]
  assign io_sram7_cen = 1'h0; // @[my_cpu_top.scala 371:14]
  assign io_sram7_wen = data_cache_io_sram_3_wen; // @[my_cpu_top.scala 371:14]
  assign io_sram7_wmask = data_cache_io_sram_3_wmask; // @[my_cpu_top.scala 371:14]
  assign io_sram7_wdata = data_cache_io_sram_3_wdata; // @[my_cpu_top.scala 371:14]
  assign u_riscv_cpu_clock = clock;
  assign u_riscv_cpu_reset = reset;
  assign u_riscv_cpu_ext_int_timer = timer_periph_io_int_line; // @[my_cpu_top.scala 255:31]
  assign u_riscv_cpu_ext_int_out_int = io_interrupt; // @[my_cpu_top.scala 256:33]
  assign u_riscv_cpu_inst_sram_rdata_L = inst_cache_io_sram_rdata_L; // @[my_cpu_top.scala 222:32]
  assign u_riscv_cpu_inst_write_en = inst_cache_io_sram_write_en; // @[my_cpu_top.scala 230:31]
  assign u_riscv_cpu_stage2_stall = inst_cache_io_stage2_stall; // @[my_cpu_top.scala 240:35]
  assign u_riscv_cpu_data_sram_rdata = data_cache_io_sram_rdata; // @[my_cpu_top.scala 209:28]
  assign u_riscv_cpu_data_stage2_stall = data_cache_io_stage2_stall; // @[my_cpu_top.scala 231:35]
  assign inst_cache_clock = clock;
  assign inst_cache_reset = reset;
  assign inst_cache_io_port_arready = _axi_cross_bar_io_m_port_0_arready; // @[my_cpu_top.scala 248:33]
  assign inst_cache_io_port_rdata = _axi_cross_bar_io_m_port_0_rdata; // @[my_cpu_top.scala 248:33]
  assign inst_cache_io_port_rlast = _axi_cross_bar_io_m_port_0_rlast; // @[my_cpu_top.scala 248:33]
  assign inst_cache_io_port_rvalid = _axi_cross_bar_io_m_port_0_rvalid; // @[my_cpu_top.scala 248:33]
  assign inst_cache_io_stage2_flush = u_riscv_cpu_stage2_flush; // @[my_cpu_top.scala 243:31]
  assign inst_cache_io_stage1_valid_flush = u_riscv_cpu_stage1_valid_flush; // @[my_cpu_top.scala 361:37]
  assign inst_cache_io_inst_ready_to_use = u_riscv_cpu_inst_ready_to_use; // @[my_cpu_top.scala 362:36]
  assign inst_cache_io_inst_buffer_full = u_riscv_cpu_inst_buffer_full; // @[my_cpu_top.scala 363:37]
  assign inst_cache_io_p_addr_for_tlb = inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 180:38]
  assign inst_cache_io_sram_req = u_riscv_cpu_inst_sram_en; // @[my_cpu_top.scala 216:29]
  assign inst_cache_io_sram_addr = u_riscv_cpu_inst_sram_addr; // @[my_cpu_top.scala 213:29]
  assign inst_cache_io_sram_cache = u_riscv_cpu_inst_cache; // @[my_cpu_top.scala 215:29]
  assign inst_cache_io_tag_valid_flush = u_riscv_cpu_icache_tag_flush; // @[my_cpu_top.scala 244:34]
  assign inst_cache_io_sram_0_rdata = io_sram0_rdata; // @[my_cpu_top.scala 364:14]
  assign inst_cache_io_sram_1_rdata = io_sram1_rdata; // @[my_cpu_top.scala 365:14]
  assign inst_cache_io_sram_2_rdata = io_sram2_rdata; // @[my_cpu_top.scala 366:14]
  assign inst_cache_io_sram_3_rdata = io_sram3_rdata; // @[my_cpu_top.scala 367:14]
  assign data_cache_clock = clock;
  assign data_cache_reset = reset;
  assign data_cache_io_port_arready = _axi_cross_bar_io_m_port_1_arready; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_rdata = _axi_cross_bar_io_m_port_1_rdata; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_rlast = _axi_cross_bar_io_m_port_1_rlast; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_rvalid = _axi_cross_bar_io_m_port_1_rvalid; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_awready = _axi_cross_bar_io_m_port_1_awready; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_wready = _axi_cross_bar_io_m_port_1_wready; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_port_bvalid = _axi_cross_bar_io_m_port_1_bvalid; // @[my_cpu_top.scala 249:33]
  assign data_cache_io_p_addr_for_tlb = data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 181:38]
  assign data_cache_io_data_wstrb = u_riscv_cpu_data_wstrb; // @[my_cpu_top.scala 208:29]
  assign data_cache_io_sram_req = u_riscv_cpu_data_sram_en; // @[my_cpu_top.scala 204:23]
  assign data_cache_io_sram_wr = u_riscv_cpu_data_sram_wen; // @[my_cpu_top.scala 205:23]
  assign data_cache_io_sram_size = {{1'd0}, u_riscv_cpu_data_size}; // @[my_cpu_top.scala 202:22]
  assign data_cache_io_sram_addr = u_riscv_cpu_data_sram_addr; // @[my_cpu_top.scala 201:22]
  assign data_cache_io_sram_wdata = u_riscv_cpu_data_sram_wdata; // @[my_cpu_top.scala 206:23]
  assign data_cache_io_sram_cache = u_riscv_cpu_data_cache; // @[my_cpu_top.scala 203:23]
  assign data_cache_io_fence_i_control = u_riscv_cpu_data_fence_i_control; // @[my_cpu_top.scala 207:28]
  assign data_cache_io_sram_0_rdata = io_sram4_rdata; // @[my_cpu_top.scala 368:14]
  assign data_cache_io_sram_1_rdata = io_sram5_rdata; // @[my_cpu_top.scala 369:14]
  assign data_cache_io_sram_2_rdata = io_sram6_rdata; // @[my_cpu_top.scala 370:14]
  assign data_cache_io_sram_3_rdata = io_sram7_rdata; // @[my_cpu_top.scala 371:14]
  assign _axi_cross_bar_clock = clock;
  assign _axi_cross_bar_reset = reset;
  assign _axi_cross_bar_io_m_port_0_araddr = inst_cache_io_port_araddr; // @[my_cpu_top.scala 248:33]
  assign _axi_cross_bar_io_m_port_0_arlen = inst_cache_io_port_arlen; // @[my_cpu_top.scala 248:33]
  assign _axi_cross_bar_io_m_port_0_arsize = inst_cache_io_port_arsize; // @[my_cpu_top.scala 248:33]
  assign _axi_cross_bar_io_m_port_0_arburst = inst_cache_io_port_arburst; // @[my_cpu_top.scala 248:33]
  assign _axi_cross_bar_io_m_port_0_arvalid = inst_cache_io_port_arvalid; // @[my_cpu_top.scala 248:33]
  assign _axi_cross_bar_io_m_port_1_araddr = data_cache_io_port_araddr; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_arlen = data_cache_io_port_arlen; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_arsize = data_cache_io_port_arsize; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_arburst = data_cache_io_port_arburst; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_arvalid = data_cache_io_port_arvalid; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_awaddr = data_cache_io_port_awaddr; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_awlen = data_cache_io_port_awlen; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_awsize = data_cache_io_port_awsize; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_awburst = data_cache_io_port_awburst; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_awvalid = data_cache_io_port_awvalid; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_wdata = data_cache_io_port_wdata; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_wstrb = data_cache_io_port_wstrb; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_wlast = data_cache_io_port_wlast; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_m_port_1_wvalid = data_cache_io_port_wvalid; // @[my_cpu_top.scala 249:33]
  assign _axi_cross_bar_io_s_port_0_arready = io_master_arready; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_rdata = io_master_rdata; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_rlast = io_master_rlast; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_rvalid = io_master_rvalid; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_awready = io_master_awready; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_wready = io_master_wready; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_0_bvalid = io_master_bvalid; // @[my_cpu_top.scala 246:15]
  assign _axi_cross_bar_io_s_port_1_rdata = timer_periph_io_axi_port_rdata; // @[my_cpu_top.scala 253:33]
  assign _axi_cross_bar_io_s_port_1_rlast = timer_periph_io_axi_port_rlast; // @[my_cpu_top.scala 253:33]
  assign _axi_cross_bar_io_s_port_1_rvalid = timer_periph_io_axi_port_rvalid; // @[my_cpu_top.scala 253:33]
  assign _axi_cross_bar_io_s_port_1_wready = timer_periph_io_axi_port_wready; // @[my_cpu_top.scala 253:33]
  assign _axi_cross_bar_io_s_port_1_bvalid = timer_periph_io_axi_port_bvalid; // @[my_cpu_top.scala 253:33]
  assign timer_periph_clock = clock;
  assign timer_periph_reset = reset;
  assign timer_periph_io_axi_port_araddr = _axi_cross_bar_io_s_port_1_araddr; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_arvalid = _axi_cross_bar_io_s_port_1_arvalid; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_rready = _axi_cross_bar_io_s_port_1_rready; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_awaddr = _axi_cross_bar_io_s_port_1_awaddr; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_awsize = _axi_cross_bar_io_s_port_1_awsize; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_awvalid = _axi_cross_bar_io_s_port_1_awvalid; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_wdata = _axi_cross_bar_io_s_port_1_wdata; // @[my_cpu_top.scala 253:33]
  assign timer_periph_io_axi_port_wvalid = _axi_cross_bar_io_s_port_1_wvalid; // @[my_cpu_top.scala 253:33]
endmodule
